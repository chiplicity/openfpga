magic
tech EFS8A
magscale 1 2
timestamp 1603800963
<< locali >>
rect 9861 17051 9895 17289
<< viali >>
rect 13148 25313 13182 25347
rect 20784 25313 20818 25347
rect 13219 25109 13253 25143
rect 20855 25109 20889 25143
rect 13173 24905 13207 24939
rect 20809 24905 20843 24939
rect 11333 24769 11367 24803
rect 24305 24769 24339 24803
rect 25409 24769 25443 24803
rect 10940 24701 10974 24735
rect 12656 24701 12690 24735
rect 13449 24701 13483 24735
rect 14277 24701 14311 24735
rect 14829 24701 14863 24735
rect 15448 24701 15482 24735
rect 15841 24701 15875 24735
rect 19705 24701 19739 24735
rect 20165 24701 20199 24735
rect 21488 24701 21522 24735
rect 21913 24701 21947 24735
rect 23912 24701 23946 24735
rect 24924 24701 24958 24735
rect 12759 24633 12793 24667
rect 20533 24633 20567 24667
rect 11011 24565 11045 24599
rect 14461 24565 14495 24599
rect 15519 24565 15553 24599
rect 17681 24565 17715 24599
rect 21591 24565 21625 24599
rect 23983 24565 24017 24599
rect 24995 24565 25029 24599
rect 15013 24361 15047 24395
rect 18509 24361 18543 24395
rect 22281 24361 22315 24395
rect 23569 24361 23603 24395
rect 20625 24293 20659 24327
rect 5972 24225 6006 24259
rect 8088 24225 8122 24259
rect 9284 24225 9318 24259
rect 12805 24225 12839 24259
rect 13792 24225 13826 24259
rect 14829 24225 14863 24259
rect 16853 24225 16887 24259
rect 18325 24225 18359 24259
rect 22097 24225 22131 24259
rect 23385 24225 23419 24259
rect 24556 24225 24590 24259
rect 11149 24157 11183 24191
rect 12161 24157 12195 24191
rect 20533 24157 20567 24191
rect 20809 24157 20843 24191
rect 24627 24089 24661 24123
rect 6043 24021 6077 24055
rect 8159 24021 8193 24055
rect 9355 24021 9389 24055
rect 13863 24021 13897 24055
rect 17221 24021 17255 24055
rect 17773 24021 17807 24055
rect 1903 23817 1937 23851
rect 2225 23817 2259 23851
rect 3237 23817 3271 23851
rect 5353 23817 5387 23851
rect 5997 23817 6031 23851
rect 7377 23817 7411 23851
rect 8389 23817 8423 23851
rect 9309 23817 9343 23851
rect 10321 23817 10355 23851
rect 10965 23817 10999 23851
rect 11701 23817 11735 23851
rect 12161 23817 12195 23851
rect 13817 23817 13851 23851
rect 14047 23817 14081 23851
rect 14369 23817 14403 23851
rect 19705 23817 19739 23851
rect 20533 23817 20567 23851
rect 22097 23817 22131 23851
rect 22649 23817 22683 23851
rect 24581 23817 24615 23851
rect 25317 23817 25351 23851
rect 8113 23749 8147 23783
rect 16623 23749 16657 23783
rect 18693 23749 18727 23783
rect 12437 23681 12471 23715
rect 20717 23681 20751 23715
rect 21637 23681 21671 23715
rect 1832 23613 1866 23647
rect 2844 23613 2878 23647
rect 4960 23613 4994 23647
rect 6984 23613 7018 23647
rect 8608 23613 8642 23647
rect 9836 23613 9870 23647
rect 10781 23613 10815 23647
rect 11333 23613 11367 23647
rect 13944 23613 13978 23647
rect 15289 23613 15323 23647
rect 16520 23613 16554 23647
rect 19521 23613 19555 23647
rect 23017 23613 23051 23647
rect 23293 23613 23327 23647
rect 24832 23613 24866 23647
rect 12529 23545 12563 23579
rect 13081 23545 13115 23579
rect 14829 23545 14863 23579
rect 17773 23545 17807 23579
rect 17865 23545 17899 23579
rect 18417 23545 18451 23579
rect 20809 23545 20843 23579
rect 21361 23545 21395 23579
rect 23201 23545 23235 23579
rect 2915 23477 2949 23511
rect 5031 23477 5065 23511
rect 7055 23477 7089 23511
rect 8711 23477 8745 23511
rect 9907 23477 9941 23511
rect 15197 23477 15231 23511
rect 16301 23477 16335 23511
rect 16945 23477 16979 23511
rect 17405 23477 17439 23511
rect 19429 23477 19463 23511
rect 20165 23477 20199 23511
rect 24903 23477 24937 23511
rect 20993 23273 21027 23307
rect 24627 23273 24661 23307
rect 10873 23205 10907 23239
rect 10965 23205 10999 23239
rect 12253 23205 12287 23239
rect 12529 23205 12563 23239
rect 13081 23205 13115 23239
rect 13909 23205 13943 23239
rect 15197 23205 15231 23239
rect 16761 23205 16795 23239
rect 18325 23205 18359 23239
rect 21453 23205 21487 23239
rect 21545 23205 21579 23239
rect 23017 23205 23051 23239
rect 23109 23205 23143 23239
rect 9861 23137 9895 23171
rect 24556 23137 24590 23171
rect 9217 23069 9251 23103
rect 11517 23069 11551 23103
rect 12437 23069 12471 23103
rect 15105 23069 15139 23103
rect 15749 23069 15783 23103
rect 16669 23069 16703 23103
rect 17313 23069 17347 23103
rect 18233 23069 18267 23103
rect 18509 23069 18543 23103
rect 22097 23069 22131 23103
rect 23293 23069 23327 23103
rect 17681 23001 17715 23035
rect 16025 22933 16059 22967
rect 20717 22933 20751 22967
rect 9217 22729 9251 22763
rect 10321 22729 10355 22763
rect 11011 22729 11045 22763
rect 11333 22729 11367 22763
rect 15381 22729 15415 22763
rect 16945 22729 16979 22763
rect 17313 22729 17347 22763
rect 18969 22729 19003 22763
rect 19291 22729 19325 22763
rect 21637 22729 21671 22763
rect 23017 22729 23051 22763
rect 24213 22729 24247 22763
rect 22005 22661 22039 22695
rect 12437 22593 12471 22627
rect 13357 22593 13391 22627
rect 14093 22593 14127 22627
rect 15105 22593 15139 22627
rect 15657 22593 15691 22627
rect 15933 22593 15967 22627
rect 17957 22593 17991 22627
rect 21361 22593 21395 22627
rect 23293 22593 23327 22627
rect 23569 22593 23603 22627
rect 24581 22593 24615 22627
rect 10908 22525 10942 22559
rect 14737 22525 14771 22559
rect 19188 22525 19222 22559
rect 19613 22525 19647 22559
rect 8297 22457 8331 22491
rect 8849 22457 8883 22491
rect 9401 22457 9435 22491
rect 9493 22457 9527 22491
rect 10045 22457 10079 22491
rect 10689 22457 10723 22491
rect 12069 22457 12103 22491
rect 12161 22457 12195 22491
rect 14185 22457 14219 22491
rect 15749 22457 15783 22491
rect 17681 22457 17715 22491
rect 17773 22457 17807 22491
rect 20717 22457 20751 22491
rect 20809 22457 20843 22491
rect 23385 22457 23419 22491
rect 11793 22389 11827 22423
rect 12989 22389 13023 22423
rect 13817 22389 13851 22423
rect 16669 22389 16703 22423
rect 18601 22389 18635 22423
rect 20533 22389 20567 22423
rect 22649 22389 22683 22423
rect 10873 22185 10907 22219
rect 11885 22185 11919 22219
rect 14185 22185 14219 22219
rect 19337 22185 19371 22219
rect 23845 22185 23879 22219
rect 9585 22117 9619 22151
rect 10137 22117 10171 22151
rect 15013 22117 15047 22151
rect 15565 22117 15599 22151
rect 18141 22117 18175 22151
rect 20625 22117 20659 22151
rect 23017 22117 23051 22151
rect 23569 22117 23603 22151
rect 1004 22049 1038 22083
rect 11701 22049 11735 22083
rect 13817 22049 13851 22083
rect 13909 22049 13943 22083
rect 17773 22049 17807 22083
rect 24464 22049 24498 22083
rect 9493 21981 9527 22015
rect 14921 21981 14955 22015
rect 20533 21981 20567 22015
rect 20809 21981 20843 22015
rect 22925 21981 22959 22015
rect 1075 21845 1109 21879
rect 12713 21845 12747 21879
rect 15841 21845 15875 21879
rect 18509 21845 18543 21879
rect 24535 21845 24569 21879
rect 1121 21641 1155 21675
rect 4249 21641 4283 21675
rect 9953 21641 9987 21675
rect 11609 21641 11643 21675
rect 12529 21641 12563 21675
rect 13081 21641 13115 21675
rect 14461 21641 14495 21675
rect 14921 21641 14955 21675
rect 17773 21641 17807 21675
rect 20625 21641 20659 21675
rect 22097 21641 22131 21675
rect 22557 21641 22591 21675
rect 24489 21641 24523 21675
rect 25317 21641 25351 21675
rect 15841 21573 15875 21607
rect 21361 21573 21395 21607
rect 7469 21505 7503 21539
rect 8113 21505 8147 21539
rect 9309 21505 9343 21539
rect 10321 21505 10355 21539
rect 15289 21505 15323 21539
rect 18969 21505 19003 21539
rect 22925 21505 22959 21539
rect 23201 21505 23235 21539
rect 3856 21437 3890 21471
rect 12136 21437 12170 21471
rect 13541 21437 13575 21471
rect 19889 21437 19923 21471
rect 20717 21437 20751 21471
rect 21913 21437 21947 21471
rect 23293 21437 23327 21471
rect 24832 21437 24866 21471
rect 7285 21369 7319 21403
rect 7561 21369 7595 21403
rect 9033 21369 9067 21403
rect 9125 21369 9159 21403
rect 13357 21369 13391 21403
rect 13862 21369 13896 21403
rect 18509 21369 18543 21403
rect 18601 21369 18635 21403
rect 3927 21301 3961 21335
rect 8757 21301 8791 21335
rect 12207 21301 12241 21335
rect 18325 21301 18359 21335
rect 20257 21301 20291 21335
rect 21729 21301 21763 21335
rect 24903 21301 24937 21335
rect 7469 21097 7503 21131
rect 10229 21097 10263 21131
rect 12253 21097 12287 21131
rect 17313 21097 17347 21131
rect 22925 21097 22959 21131
rect 24305 21097 24339 21131
rect 8297 21029 8331 21063
rect 9671 21029 9705 21063
rect 11695 21029 11729 21063
rect 16755 21029 16789 21063
rect 18693 21029 18727 21063
rect 18969 21029 19003 21063
rect 20441 21029 20475 21063
rect 8205 20961 8239 20995
rect 15105 20961 15139 20995
rect 15381 20961 15415 20995
rect 20533 20961 20567 20995
rect 24121 20961 24155 20995
rect 9309 20893 9343 20927
rect 11333 20893 11367 20927
rect 15565 20893 15599 20927
rect 15841 20893 15875 20927
rect 16393 20893 16427 20927
rect 18877 20893 18911 20927
rect 19521 20893 19555 20927
rect 9033 20757 9067 20791
rect 13633 20757 13667 20791
rect 14001 20757 14035 20791
rect 17681 20757 17715 20791
rect 23385 20757 23419 20791
rect 7653 20553 7687 20587
rect 9953 20553 9987 20587
rect 12897 20553 12931 20587
rect 14921 20553 14955 20587
rect 16669 20553 16703 20587
rect 20533 20553 20567 20587
rect 22189 20553 22223 20587
rect 24949 20553 24983 20587
rect 25271 20553 25305 20587
rect 24581 20485 24615 20519
rect 10229 20417 10263 20451
rect 15749 20417 15783 20451
rect 18325 20417 18359 20451
rect 19521 20417 19555 20451
rect 8205 20349 8239 20383
rect 9033 20349 9067 20383
rect 11977 20349 12011 20383
rect 14001 20349 14035 20383
rect 16945 20349 16979 20383
rect 21269 20349 21303 20383
rect 24188 20349 24222 20383
rect 25200 20349 25234 20383
rect 25593 20349 25627 20383
rect 8573 20281 8607 20315
rect 8941 20281 8975 20315
rect 9395 20281 9429 20315
rect 11057 20281 11091 20315
rect 12339 20281 12373 20315
rect 13817 20281 13851 20315
rect 14322 20281 14356 20315
rect 15565 20281 15599 20315
rect 16070 20281 16104 20315
rect 17313 20281 17347 20315
rect 17681 20281 17715 20315
rect 17773 20281 17807 20315
rect 19245 20281 19279 20315
rect 19337 20281 19371 20315
rect 21590 20281 21624 20315
rect 11333 20213 11367 20247
rect 11701 20213 11735 20247
rect 15289 20213 15323 20247
rect 18601 20213 18635 20247
rect 18969 20213 19003 20247
rect 21085 20213 21119 20247
rect 24259 20213 24293 20247
rect 9585 20009 9619 20043
rect 17405 20009 17439 20043
rect 18601 20009 18635 20043
rect 18969 20009 19003 20043
rect 20579 20009 20613 20043
rect 22465 20009 22499 20043
rect 13909 19941 13943 19975
rect 15657 19941 15691 19975
rect 16806 19941 16840 19975
rect 21866 19941 21900 19975
rect 9493 19873 9527 19907
rect 9953 19873 9987 19907
rect 11517 19873 11551 19907
rect 11977 19873 12011 19907
rect 13357 19873 13391 19907
rect 13725 19873 13759 19907
rect 14921 19873 14955 19907
rect 15381 19873 15415 19907
rect 17681 19873 17715 19907
rect 18877 19873 18911 19907
rect 20476 19873 20510 19907
rect 23661 19873 23695 19907
rect 24924 19873 24958 19907
rect 12069 19805 12103 19839
rect 12529 19805 12563 19839
rect 16485 19805 16519 19839
rect 21545 19805 21579 19839
rect 24995 19737 25029 19771
rect 14645 19669 14679 19703
rect 21269 19669 21303 19703
rect 23569 19669 23603 19703
rect 16485 19465 16519 19499
rect 18877 19465 18911 19499
rect 20993 19465 21027 19499
rect 25409 19465 25443 19499
rect 14921 19397 14955 19431
rect 17313 19329 17347 19363
rect 24029 19329 24063 19363
rect 9217 19261 9251 19295
rect 9493 19261 9527 19295
rect 9769 19261 9803 19295
rect 11517 19261 11551 19295
rect 12069 19261 12103 19295
rect 12529 19261 12563 19295
rect 13725 19261 13759 19295
rect 14001 19261 14035 19295
rect 14553 19261 14587 19295
rect 15289 19261 15323 19295
rect 15749 19261 15783 19295
rect 16025 19261 16059 19295
rect 16853 19261 16887 19295
rect 17589 19261 17623 19295
rect 18509 19261 18543 19295
rect 19797 19261 19831 19295
rect 20717 19261 20751 19295
rect 22649 19261 22683 19295
rect 24924 19261 24958 19295
rect 25777 19261 25811 19295
rect 8849 19193 8883 19227
rect 13173 19193 13207 19227
rect 17910 19193 17944 19227
rect 19613 19193 19647 19227
rect 20118 19193 20152 19227
rect 21545 19193 21579 19227
rect 22097 19193 22131 19227
rect 23385 19193 23419 19227
rect 23477 19193 23511 19227
rect 9401 19125 9435 19159
rect 10321 19125 10355 19159
rect 10873 19125 10907 19159
rect 11149 19125 11183 19159
rect 12069 19125 12103 19159
rect 13633 19125 13667 19159
rect 21913 19125 21947 19159
rect 23017 19125 23051 19159
rect 24995 19125 25029 19159
rect 13265 18921 13299 18955
rect 17773 18921 17807 18955
rect 23385 18921 23419 18955
rect 9861 18853 9895 18887
rect 9953 18853 9987 18887
rect 16577 18853 16611 18887
rect 17589 18853 17623 18887
rect 19521 18853 19555 18887
rect 19797 18853 19831 18887
rect 21177 18853 21211 18887
rect 23661 18853 23695 18887
rect 24213 18853 24247 18887
rect 15289 18785 15323 18819
rect 15841 18785 15875 18819
rect 16301 18785 16335 18819
rect 18877 18785 18911 18819
rect 19245 18785 19279 18819
rect 20717 18785 20751 18819
rect 20993 18785 21027 18819
rect 10505 18717 10539 18751
rect 11333 18717 11367 18751
rect 11977 18717 12011 18751
rect 13909 18717 13943 18751
rect 14645 18717 14679 18751
rect 23569 18717 23603 18751
rect 9585 18581 9619 18615
rect 10781 18581 10815 18615
rect 12345 18581 12379 18615
rect 13633 18581 13667 18615
rect 15657 18581 15691 18615
rect 21453 18581 21487 18615
rect 11333 18377 11367 18411
rect 13679 18377 13713 18411
rect 14001 18377 14035 18411
rect 15841 18377 15875 18411
rect 16577 18377 16611 18411
rect 19061 18377 19095 18411
rect 20165 18377 20199 18411
rect 21177 18377 21211 18411
rect 22281 18377 22315 18411
rect 22649 18377 22683 18411
rect 12621 18309 12655 18343
rect 13817 18309 13851 18343
rect 10413 18241 10447 18275
rect 10689 18241 10723 18275
rect 12069 18241 12103 18275
rect 13909 18241 13943 18275
rect 19245 18241 19279 18275
rect 24213 18241 24247 18275
rect 8665 18173 8699 18207
rect 9401 18173 9435 18207
rect 9861 18173 9895 18207
rect 18233 18173 18267 18207
rect 18693 18173 18727 18207
rect 21361 18173 21395 18207
rect 9493 18105 9527 18139
rect 10137 18105 10171 18139
rect 10505 18105 10539 18139
rect 11793 18105 11827 18139
rect 12161 18105 12195 18139
rect 13081 18105 13115 18139
rect 13541 18105 13575 18139
rect 19566 18105 19600 18139
rect 21682 18105 21716 18139
rect 23017 18105 23051 18139
rect 23937 18105 23971 18139
rect 24029 18105 24063 18139
rect 13449 18037 13483 18071
rect 14553 18037 14587 18071
rect 15013 18037 15047 18071
rect 15289 18037 15323 18071
rect 16209 18037 16243 18071
rect 18141 18037 18175 18071
rect 18417 18037 18451 18071
rect 20441 18037 20475 18071
rect 20809 18037 20843 18071
rect 23661 18037 23695 18071
rect 10413 17833 10447 17867
rect 13817 17833 13851 17867
rect 14553 17833 14587 17867
rect 16577 17833 16611 17867
rect 23569 17833 23603 17867
rect 9814 17765 9848 17799
rect 11701 17765 11735 17799
rect 12253 17765 12287 17799
rect 13081 17765 13115 17799
rect 15565 17765 15599 17799
rect 19429 17765 19463 17799
rect 19705 17765 19739 17799
rect 21177 17765 21211 17799
rect 22326 17765 22360 17799
rect 23937 17765 23971 17799
rect 13173 17697 13207 17731
rect 14829 17697 14863 17731
rect 14976 17697 15010 17731
rect 16393 17697 16427 17731
rect 18693 17697 18727 17731
rect 19153 17697 19187 17731
rect 20717 17697 20751 17731
rect 20993 17697 21027 17731
rect 22925 17697 22959 17731
rect 9493 17629 9527 17663
rect 11609 17629 11643 17663
rect 13541 17629 13575 17663
rect 15197 17629 15231 17663
rect 22005 17629 22039 17663
rect 23845 17629 23879 17663
rect 15933 17561 15967 17595
rect 24397 17561 24431 17595
rect 10689 17493 10723 17527
rect 12713 17493 12747 17527
rect 13311 17493 13345 17527
rect 13449 17493 13483 17527
rect 14277 17493 14311 17527
rect 15105 17493 15139 17527
rect 16853 17493 16887 17527
rect 17681 17493 17715 17527
rect 20165 17493 20199 17527
rect 21453 17493 21487 17527
rect 9677 17289 9711 17323
rect 9861 17289 9895 17323
rect 9953 17289 9987 17323
rect 11609 17289 11643 17323
rect 12970 17289 13004 17323
rect 13449 17289 13483 17323
rect 15013 17289 15047 17323
rect 16577 17289 16611 17323
rect 18693 17289 18727 17323
rect 21637 17289 21671 17323
rect 23661 17289 23695 17323
rect 25087 17289 25121 17323
rect 25501 17289 25535 17323
rect 9309 17153 9343 17187
rect 8849 17085 8883 17119
rect 9125 17085 9159 17119
rect 13081 17221 13115 17255
rect 14645 17221 14679 17255
rect 15381 17221 15415 17255
rect 16209 17221 16243 17255
rect 17037 17221 17071 17255
rect 12713 17153 12747 17187
rect 13173 17153 13207 17187
rect 14737 17153 14771 17187
rect 16301 17153 16335 17187
rect 17681 17153 17715 17187
rect 17957 17153 17991 17187
rect 21361 17153 21395 17187
rect 10137 17085 10171 17119
rect 11057 17085 11091 17119
rect 12345 17085 12379 17119
rect 14516 17085 14550 17119
rect 15749 17085 15783 17119
rect 16080 17085 16114 17119
rect 19153 17085 19187 17119
rect 20165 17085 20199 17119
rect 20533 17085 20567 17119
rect 20809 17085 20843 17119
rect 21085 17085 21119 17119
rect 22005 17085 22039 17119
rect 23017 17085 23051 17119
rect 24029 17085 24063 17119
rect 24397 17085 24431 17119
rect 25016 17085 25050 17119
rect 8481 17017 8515 17051
rect 9861 17017 9895 17051
rect 10458 17017 10492 17051
rect 12805 17017 12839 17051
rect 14369 17017 14403 17051
rect 15933 17017 15967 17051
rect 17773 17017 17807 17051
rect 19613 17017 19647 17051
rect 13817 16949 13851 16983
rect 14185 16949 14219 16983
rect 17313 16949 17347 16983
rect 19337 16949 19371 16983
rect 22373 16949 22407 16983
rect 8665 16745 8699 16779
rect 9493 16745 9527 16779
rect 11333 16745 11367 16779
rect 11793 16745 11827 16779
rect 12897 16745 12931 16779
rect 13817 16745 13851 16779
rect 15013 16745 15047 16779
rect 15289 16745 15323 16779
rect 18693 16745 18727 16779
rect 24121 16745 24155 16779
rect 10689 16677 10723 16711
rect 15657 16677 15691 16711
rect 16025 16677 16059 16711
rect 16117 16677 16151 16711
rect 21361 16677 21395 16711
rect 23339 16677 23373 16711
rect 10229 16609 10263 16643
rect 10413 16609 10447 16643
rect 11793 16609 11827 16643
rect 13173 16609 13207 16643
rect 14829 16609 14863 16643
rect 17589 16609 17623 16643
rect 18233 16609 18267 16643
rect 19061 16609 19095 16643
rect 20717 16609 20751 16643
rect 21085 16609 21119 16643
rect 23236 16609 23270 16643
rect 23661 16609 23695 16643
rect 24280 16609 24314 16643
rect 13541 16541 13575 16575
rect 16669 16541 16703 16575
rect 13449 16473 13483 16507
rect 13311 16405 13345 16439
rect 14369 16405 14403 16439
rect 24351 16405 24385 16439
rect 9677 16201 9711 16235
rect 10321 16201 10355 16235
rect 10781 16201 10815 16235
rect 11609 16201 11643 16235
rect 12897 16201 12931 16235
rect 14231 16201 14265 16235
rect 14737 16201 14771 16235
rect 15105 16201 15139 16235
rect 18877 16201 18911 16235
rect 24305 16201 24339 16235
rect 24949 16201 24983 16235
rect 14369 16133 14403 16167
rect 13633 16065 13667 16099
rect 14001 16065 14035 16099
rect 14461 16065 14495 16099
rect 16669 16065 16703 16099
rect 19521 16065 19555 16099
rect 20165 16065 20199 16099
rect 22649 16065 22683 16099
rect 23293 16065 23327 16099
rect 9493 15997 9527 16031
rect 16577 15997 16611 16031
rect 16945 15997 16979 16031
rect 18509 15997 18543 16031
rect 24765 15997 24799 16031
rect 25317 15997 25351 16031
rect 14093 15929 14127 15963
rect 18601 15929 18635 15963
rect 19613 15929 19647 15963
rect 20717 15929 20751 15963
rect 23385 15929 23419 15963
rect 23937 15929 23971 15963
rect 10045 15861 10079 15895
rect 12529 15861 12563 15895
rect 13265 15861 13299 15895
rect 15473 15861 15507 15895
rect 17313 15861 17347 15895
rect 19337 15861 19371 15895
rect 20993 15861 21027 15895
rect 23017 15861 23051 15895
rect 14093 15657 14127 15691
rect 15841 15657 15875 15691
rect 16209 15657 16243 15691
rect 17589 15657 17623 15691
rect 17957 15657 17991 15691
rect 18233 15657 18267 15691
rect 23569 15657 23603 15691
rect 15283 15589 15317 15623
rect 16485 15589 16519 15623
rect 16990 15589 17024 15623
rect 18601 15589 18635 15623
rect 19153 15589 19187 15623
rect 21913 15589 21947 15623
rect 22465 15589 22499 15623
rect 23385 15521 23419 15555
rect 24892 15521 24926 15555
rect 14921 15453 14955 15487
rect 16669 15453 16703 15487
rect 18509 15453 18543 15487
rect 20441 15453 20475 15487
rect 21821 15453 21855 15487
rect 13265 15317 13299 15351
rect 14461 15317 14495 15351
rect 19429 15317 19463 15351
rect 20993 15317 21027 15351
rect 24995 15317 25029 15351
rect 15749 15113 15783 15147
rect 16761 15113 16795 15147
rect 17221 15113 17255 15147
rect 18601 15113 18635 15147
rect 19061 15113 19095 15147
rect 21913 15113 21947 15147
rect 22281 15113 22315 15147
rect 23385 15113 23419 15147
rect 24029 15113 24063 15147
rect 22557 15045 22591 15079
rect 17681 14977 17715 15011
rect 14277 14909 14311 14943
rect 14645 14909 14679 14943
rect 14829 14909 14863 14943
rect 15197 14909 15231 14943
rect 16301 14909 16335 14943
rect 20993 14909 21027 14943
rect 24121 14909 24155 14943
rect 16117 14841 16151 14875
rect 17773 14841 17807 14875
rect 18325 14841 18359 14875
rect 19245 14841 19279 14875
rect 19337 14841 19371 14875
rect 19889 14841 19923 14875
rect 20901 14841 20935 14875
rect 21355 14841 21389 14875
rect 13909 14773 13943 14807
rect 15473 14773 15507 14807
rect 16485 14773 16519 14807
rect 24305 14773 24339 14807
rect 24857 14773 24891 14807
rect 14001 14569 14035 14603
rect 14921 14569 14955 14603
rect 16669 14569 16703 14603
rect 17681 14569 17715 14603
rect 22097 14569 22131 14603
rect 23201 14569 23235 14603
rect 14461 14501 14495 14535
rect 18094 14501 18128 14535
rect 20625 14501 20659 14535
rect 14921 14433 14955 14467
rect 15289 14433 15323 14467
rect 15657 14433 15691 14467
rect 22005 14433 22039 14467
rect 22465 14433 22499 14467
rect 24213 14433 24247 14467
rect 17773 14365 17807 14399
rect 20533 14365 20567 14399
rect 20809 14365 20843 14399
rect 23569 14365 23603 14399
rect 18693 14229 18727 14263
rect 19153 14229 19187 14263
rect 21453 14229 21487 14263
rect 13173 14025 13207 14059
rect 15749 14025 15783 14059
rect 17865 14025 17899 14059
rect 20809 14025 20843 14059
rect 22281 14025 22315 14059
rect 23017 14025 23051 14059
rect 24213 14025 24247 14059
rect 14185 13957 14219 13991
rect 22557 13957 22591 13991
rect 19797 13889 19831 13923
rect 20441 13889 20475 13923
rect 21269 13889 21303 13923
rect 23293 13889 23327 13923
rect 12989 13821 13023 13855
rect 13449 13821 13483 13855
rect 13909 13821 13943 13855
rect 14369 13821 14403 13855
rect 15013 13821 15047 13855
rect 15197 13821 15231 13855
rect 16117 13821 16151 13855
rect 16485 13821 16519 13855
rect 18141 13821 18175 13855
rect 18969 13821 19003 13855
rect 19153 13821 19187 13855
rect 21361 13821 21395 13855
rect 21682 13753 21716 13787
rect 23385 13753 23419 13787
rect 23937 13753 23971 13787
rect 15473 13685 15507 13719
rect 24765 13685 24799 13719
rect 12345 13481 12379 13515
rect 16209 13481 16243 13515
rect 22327 13481 22361 13515
rect 24949 13481 24983 13515
rect 13909 13413 13943 13447
rect 15933 13413 15967 13447
rect 17865 13413 17899 13447
rect 18877 13413 18911 13447
rect 21361 13413 21395 13447
rect 23385 13413 23419 13447
rect 23937 13413 23971 13447
rect 12161 13345 12195 13379
rect 13173 13345 13207 13379
rect 14829 13345 14863 13379
rect 15657 13345 15691 13379
rect 17773 13345 17807 13379
rect 20809 13345 20843 13379
rect 21085 13345 21119 13379
rect 22005 13345 22039 13379
rect 22224 13345 22258 13379
rect 24765 13345 24799 13379
rect 13541 13277 13575 13311
rect 15565 13277 15599 13311
rect 18785 13277 18819 13311
rect 19061 13277 19095 13311
rect 23293 13277 23327 13311
rect 13081 13209 13115 13243
rect 13338 13209 13372 13243
rect 13449 13141 13483 13175
rect 14185 13141 14219 13175
rect 14553 13141 14587 13175
rect 12897 12937 12931 12971
rect 13890 12937 13924 12971
rect 14369 12937 14403 12971
rect 14829 12937 14863 12971
rect 15565 12937 15599 12971
rect 16577 12937 16611 12971
rect 17037 12937 17071 12971
rect 18785 12937 18819 12971
rect 21821 12937 21855 12971
rect 23477 12937 23511 12971
rect 24213 12937 24247 12971
rect 24765 12937 24799 12971
rect 14001 12869 14035 12903
rect 14093 12801 14127 12835
rect 15657 12801 15691 12835
rect 19337 12801 19371 12835
rect 21361 12801 21395 12835
rect 23017 12801 23051 12835
rect 12253 12733 12287 12767
rect 13725 12733 13759 12767
rect 17405 12733 17439 12767
rect 17681 12733 17715 12767
rect 20809 12733 20843 12767
rect 21269 12733 21303 12767
rect 23728 12733 23762 12767
rect 15978 12665 16012 12699
rect 18325 12665 18359 12699
rect 19429 12665 19463 12699
rect 19981 12665 20015 12699
rect 22189 12665 22223 12699
rect 13265 12597 13299 12631
rect 13541 12597 13575 12631
rect 19061 12597 19095 12631
rect 20349 12597 20383 12631
rect 20717 12597 20751 12631
rect 23799 12597 23833 12631
rect 12897 12393 12931 12427
rect 14185 12393 14219 12427
rect 15013 12393 15047 12427
rect 16209 12393 16243 12427
rect 15841 12325 15875 12359
rect 17497 12325 17531 12359
rect 19153 12325 19187 12359
rect 19613 12325 19647 12359
rect 12713 12257 12747 12291
rect 13725 12257 13759 12291
rect 14829 12257 14863 12291
rect 20809 12257 20843 12291
rect 20993 12257 21027 12291
rect 21545 12257 21579 12291
rect 22925 12257 22959 12291
rect 13633 12189 13667 12223
rect 17405 12189 17439 12223
rect 18049 12189 18083 12223
rect 21269 12189 21303 12223
rect 23477 12189 23511 12223
rect 13265 12121 13299 12155
rect 13909 12053 13943 12087
rect 14553 12053 14587 12087
rect 15473 12053 15507 12087
rect 18785 12053 18819 12087
rect 13081 11849 13115 11883
rect 16485 11849 16519 11883
rect 17037 11849 17071 11883
rect 20625 11849 20659 11883
rect 21269 11849 21303 11883
rect 22281 11849 22315 11883
rect 22649 11849 22683 11883
rect 22925 11849 22959 11883
rect 14185 11781 14219 11815
rect 14921 11781 14955 11815
rect 15749 11781 15783 11815
rect 17313 11781 17347 11815
rect 19981 11781 20015 11815
rect 12805 11713 12839 11747
rect 14277 11713 14311 11747
rect 15841 11713 15875 11747
rect 19429 11713 19463 11747
rect 21361 11713 21395 11747
rect 12897 11645 12931 11679
rect 14056 11645 14090 11679
rect 15620 11645 15654 11679
rect 17589 11645 17623 11679
rect 13449 11577 13483 11611
rect 13909 11577 13943 11611
rect 15473 11577 15507 11611
rect 16209 11577 16243 11611
rect 17910 11577 17944 11611
rect 19521 11577 19555 11611
rect 21682 11577 21716 11611
rect 23293 11577 23327 11611
rect 23385 11577 23419 11611
rect 23937 11577 23971 11611
rect 13725 11509 13759 11543
rect 14553 11509 14587 11543
rect 15289 11509 15323 11543
rect 18509 11509 18543 11543
rect 19153 11509 19187 11543
rect 12713 11305 12747 11339
rect 13725 11305 13759 11339
rect 17313 11305 17347 11339
rect 21361 11305 21395 11339
rect 23293 11305 23327 11339
rect 15841 11237 15875 11271
rect 16755 11237 16789 11271
rect 17957 11237 17991 11271
rect 18325 11237 18359 11271
rect 20625 11237 20659 11271
rect 22142 11237 22176 11271
rect 23753 11237 23787 11271
rect 12529 11169 12563 11203
rect 13541 11169 13575 11203
rect 14829 11169 14863 11203
rect 15289 11169 15323 11203
rect 14369 11101 14403 11135
rect 15565 11101 15599 11135
rect 16393 11101 16427 11135
rect 18233 11101 18267 11135
rect 18509 11101 18543 11135
rect 19337 11101 19371 11135
rect 21821 11101 21855 11135
rect 23661 11101 23695 11135
rect 14001 11033 14035 11067
rect 17589 11033 17623 11067
rect 22741 11033 22775 11067
rect 24213 11033 24247 11067
rect 12529 10761 12563 10795
rect 13357 10761 13391 10795
rect 14093 10761 14127 10795
rect 14829 10761 14863 10795
rect 15749 10761 15783 10795
rect 17221 10761 17255 10795
rect 18233 10761 18267 10795
rect 18601 10761 18635 10795
rect 18969 10761 19003 10795
rect 22557 10761 22591 10795
rect 24397 10761 24431 10795
rect 24765 10761 24799 10795
rect 25133 10761 25167 10795
rect 16853 10693 16887 10727
rect 16577 10625 16611 10659
rect 19705 10625 19739 10659
rect 20165 10625 20199 10659
rect 23477 10625 23511 10659
rect 13541 10557 13575 10591
rect 14645 10557 14679 10591
rect 15105 10557 15139 10591
rect 15841 10557 15875 10591
rect 16301 10557 16335 10591
rect 18785 10557 18819 10591
rect 20533 10557 20567 10591
rect 20717 10557 20751 10591
rect 24949 10557 24983 10591
rect 25501 10557 25535 10591
rect 20993 10489 21027 10523
rect 23569 10489 23603 10523
rect 24121 10489 24155 10523
rect 12989 10421 13023 10455
rect 14553 10421 14587 10455
rect 17865 10421 17899 10455
rect 21821 10421 21855 10455
rect 22097 10421 22131 10455
rect 23017 10421 23051 10455
rect 14553 10217 14587 10251
rect 16301 10217 16335 10251
rect 20717 10217 20751 10251
rect 22695 10217 22729 10251
rect 24581 10217 24615 10251
rect 13909 10149 13943 10183
rect 23753 10149 23787 10183
rect 13541 10081 13575 10115
rect 14829 10081 14863 10115
rect 18877 10081 18911 10115
rect 20533 10081 20567 10115
rect 20901 10081 20935 10115
rect 22624 10081 22658 10115
rect 14976 10013 15010 10047
rect 15197 10013 15231 10047
rect 23661 10013 23695 10047
rect 23937 10013 23971 10047
rect 14277 9945 14311 9979
rect 15289 9945 15323 9979
rect 15105 9877 15139 9911
rect 15841 9877 15875 9911
rect 18969 9877 19003 9911
rect 23293 9877 23327 9911
rect 12621 9673 12655 9707
rect 21269 9673 21303 9707
rect 22925 9673 22959 9707
rect 15565 9605 15599 9639
rect 16301 9605 16335 9639
rect 18417 9605 18451 9639
rect 18785 9605 18819 9639
rect 24949 9605 24983 9639
rect 14093 9537 14127 9571
rect 15436 9537 15470 9571
rect 15657 9537 15691 9571
rect 20901 9537 20935 9571
rect 23937 9537 23971 9571
rect 24213 9537 24247 9571
rect 12253 9469 12287 9503
rect 12529 9469 12563 9503
rect 13725 9469 13759 9503
rect 14277 9469 14311 9503
rect 14829 9469 14863 9503
rect 16669 9469 16703 9503
rect 22132 9469 22166 9503
rect 22557 9469 22591 9503
rect 23293 9469 23327 9503
rect 24765 9469 24799 9503
rect 12345 9401 12379 9435
rect 13633 9401 13667 9435
rect 15289 9401 15323 9435
rect 18049 9401 18083 9435
rect 18969 9401 19003 9435
rect 19061 9401 19095 9435
rect 19613 9401 19647 9435
rect 22235 9401 22269 9435
rect 25317 9401 25351 9435
rect 13265 9333 13299 9367
rect 15105 9333 15139 9367
rect 15933 9333 15967 9367
rect 20441 9333 20475 9367
rect 13817 9129 13851 9163
rect 14645 9129 14679 9163
rect 16025 9129 16059 9163
rect 19429 9129 19463 9163
rect 21913 9129 21947 9163
rect 22649 9129 22683 9163
rect 24673 9129 24707 9163
rect 12437 9061 12471 9095
rect 16898 9061 16932 9095
rect 18509 9061 18543 9095
rect 21079 9061 21113 9095
rect 23109 9061 23143 9095
rect 13173 8993 13207 9027
rect 14185 8993 14219 9027
rect 15013 8993 15047 9027
rect 15565 8993 15599 9027
rect 20717 8993 20751 9027
rect 24489 8993 24523 9027
rect 13541 8925 13575 8959
rect 15749 8925 15783 8959
rect 16577 8925 16611 8959
rect 18417 8925 18451 8959
rect 18785 8925 18819 8959
rect 23017 8925 23051 8959
rect 13338 8857 13372 8891
rect 23569 8857 23603 8891
rect 13449 8789 13483 8823
rect 16393 8789 16427 8823
rect 17497 8789 17531 8823
rect 21637 8789 21671 8823
rect 23937 8789 23971 8823
rect 12897 8585 12931 8619
rect 13633 8585 13667 8619
rect 15473 8585 15507 8619
rect 15749 8585 15783 8619
rect 16945 8585 16979 8619
rect 17313 8585 17347 8619
rect 18509 8585 18543 8619
rect 19153 8585 19187 8619
rect 20441 8585 20475 8619
rect 20809 8585 20843 8619
rect 21269 8585 21303 8619
rect 22649 8585 22683 8619
rect 24949 8585 24983 8619
rect 13265 8449 13299 8483
rect 19429 8449 19463 8483
rect 19705 8449 19739 8483
rect 21361 8449 21395 8483
rect 23293 8449 23327 8483
rect 23569 8449 23603 8483
rect 14369 8381 14403 8415
rect 15013 8381 15047 8415
rect 15933 8381 15967 8415
rect 16393 8381 16427 8415
rect 16669 8381 16703 8415
rect 17589 8381 17623 8415
rect 22281 8381 22315 8415
rect 24765 8381 24799 8415
rect 25317 8381 25351 8415
rect 13725 8313 13759 8347
rect 17910 8313 17944 8347
rect 19521 8313 19555 8347
rect 21682 8313 21716 8347
rect 23385 8313 23419 8347
rect 24213 8313 24247 8347
rect 24581 8313 24615 8347
rect 18785 8245 18819 8279
rect 23017 8245 23051 8279
rect 13265 8041 13299 8075
rect 13817 8041 13851 8075
rect 16945 8041 16979 8075
rect 17589 8041 17623 8075
rect 18325 8041 18359 8075
rect 24765 8041 24799 8075
rect 14185 7973 14219 8007
rect 18601 7973 18635 8007
rect 21637 7973 21671 8007
rect 23201 7973 23235 8007
rect 16117 7905 16151 7939
rect 16485 7905 16519 7939
rect 24581 7905 24615 7939
rect 16669 7837 16703 7871
rect 18509 7837 18543 7871
rect 18877 7837 18911 7871
rect 21545 7837 21579 7871
rect 23109 7837 23143 7871
rect 23385 7837 23419 7871
rect 22097 7769 22131 7803
rect 15381 7701 15415 7735
rect 15749 7701 15783 7735
rect 15197 7497 15231 7531
rect 15657 7497 15691 7531
rect 16393 7497 16427 7531
rect 20993 7497 21027 7531
rect 21453 7497 21487 7531
rect 22005 7497 22039 7531
rect 23017 7497 23051 7531
rect 24949 7497 24983 7531
rect 14093 7429 14127 7463
rect 14921 7429 14955 7463
rect 15546 7429 15580 7463
rect 12621 7361 12655 7395
rect 13265 7361 13299 7395
rect 14185 7361 14219 7395
rect 15749 7361 15783 7395
rect 18509 7361 18543 7395
rect 18785 7361 18819 7395
rect 23201 7361 23235 7395
rect 12253 7293 12287 7327
rect 12897 7293 12931 7327
rect 13964 7293 13998 7327
rect 17405 7293 17439 7327
rect 17865 7293 17899 7327
rect 21637 7293 21671 7327
rect 23385 7293 23419 7327
rect 24765 7293 24799 7327
rect 25317 7293 25351 7327
rect 11793 7225 11827 7259
rect 12069 7225 12103 7259
rect 13817 7225 13851 7259
rect 15381 7225 15415 7259
rect 16117 7225 16151 7259
rect 22649 7225 22683 7259
rect 13633 7157 13667 7191
rect 14461 7157 14495 7191
rect 16853 7157 16887 7191
rect 19245 7157 19279 7191
rect 20165 7157 20199 7191
rect 24581 7157 24615 7191
rect 21637 6953 21671 6987
rect 23385 6953 23419 6987
rect 14185 6885 14219 6919
rect 17129 6885 17163 6919
rect 18877 6885 18911 6919
rect 11885 6817 11919 6851
rect 11977 6817 12011 6851
rect 12161 6817 12195 6851
rect 13449 6817 13483 6851
rect 13725 6817 13759 6851
rect 15105 6817 15139 6851
rect 15289 6817 15323 6851
rect 16577 6817 16611 6851
rect 16945 6817 16979 6851
rect 18509 6817 18543 6851
rect 21085 6817 21119 6851
rect 22833 6817 22867 6851
rect 23880 6817 23914 6851
rect 23983 6817 24017 6851
rect 24924 6817 24958 6851
rect 13909 6749 13943 6783
rect 15565 6749 15599 6783
rect 15841 6749 15875 6783
rect 18785 6749 18819 6783
rect 19429 6749 19463 6783
rect 24995 6681 25029 6715
rect 20901 6613 20935 6647
rect 12253 6409 12287 6443
rect 13541 6409 13575 6443
rect 14921 6409 14955 6443
rect 16577 6409 16611 6443
rect 16945 6409 16979 6443
rect 18509 6409 18543 6443
rect 18877 6409 18911 6443
rect 20533 6409 20567 6443
rect 20901 6409 20935 6443
rect 22097 6409 22131 6443
rect 23845 6409 23879 6443
rect 24765 6409 24799 6443
rect 13265 6341 13299 6375
rect 14553 6341 14587 6375
rect 23339 6341 23373 6375
rect 15381 6273 15415 6307
rect 17589 6273 17623 6307
rect 19337 6273 19371 6307
rect 21177 6273 21211 6307
rect 21453 6273 21487 6307
rect 22925 6273 22959 6307
rect 24351 6273 24385 6307
rect 11333 6205 11367 6239
rect 12069 6205 12103 6239
rect 23236 6205 23270 6239
rect 24264 6205 24298 6239
rect 15702 6137 15736 6171
rect 17405 6137 17439 6171
rect 17951 6137 17985 6171
rect 19245 6137 19279 6171
rect 19699 6137 19733 6171
rect 21269 6137 21303 6171
rect 11609 6069 11643 6103
rect 15197 6069 15231 6103
rect 16301 6069 16335 6103
rect 20257 6069 20291 6103
rect 25133 6069 25167 6103
rect 17589 5865 17623 5899
rect 19337 5865 19371 5899
rect 23247 5865 23281 5899
rect 15150 5797 15184 5831
rect 16761 5797 16795 5831
rect 20625 5797 20659 5831
rect 21177 5797 21211 5831
rect 14829 5729 14863 5763
rect 18233 5729 18267 5763
rect 23144 5729 23178 5763
rect 24188 5729 24222 5763
rect 16669 5661 16703 5695
rect 17313 5661 17347 5695
rect 18141 5661 18175 5695
rect 20533 5661 20567 5695
rect 11977 5593 12011 5627
rect 24259 5593 24293 5627
rect 15749 5525 15783 5559
rect 14001 5321 14035 5355
rect 14829 5321 14863 5355
rect 16393 5321 16427 5355
rect 16945 5321 16979 5355
rect 18601 5321 18635 5355
rect 20533 5321 20567 5355
rect 23385 5321 23419 5355
rect 24259 5321 24293 5355
rect 24673 5321 24707 5355
rect 25041 5321 25075 5355
rect 15013 5185 15047 5219
rect 15473 5185 15507 5219
rect 17957 5185 17991 5219
rect 19889 5185 19923 5219
rect 20901 5185 20935 5219
rect 24188 5117 24222 5151
rect 14461 5049 14495 5083
rect 15105 5049 15139 5083
rect 16485 5049 16519 5083
rect 17681 5049 17715 5083
rect 17773 5049 17807 5083
rect 19061 5049 19095 5083
rect 19613 5049 19647 5083
rect 19705 5049 19739 5083
rect 17405 4981 17439 5015
rect 19429 4981 19463 5015
rect 15013 4777 15047 4811
rect 17681 4777 17715 4811
rect 24259 4777 24293 4811
rect 15933 4709 15967 4743
rect 16485 4709 16519 4743
rect 19521 4709 19555 4743
rect 18877 4641 18911 4675
rect 24188 4641 24222 4675
rect 15841 4573 15875 4607
rect 14921 4233 14955 4267
rect 18877 4233 18911 4267
rect 15841 4097 15875 4131
rect 16117 4097 16151 4131
rect 16485 4097 16519 4131
rect 25041 4097 25075 4131
rect 15197 4029 15231 4063
rect 24172 4029 24206 4063
rect 24259 3961 24293 3995
rect 24673 3893 24707 3927
rect 16347 3689 16381 3723
rect 16276 3553 16310 3587
rect 16301 2941 16335 2975
rect 24259 2601 24293 2635
rect 24188 2465 24222 2499
rect 24673 2261 24707 2295
<< metal1 >>
rect 632 25594 26392 25616
rect 632 25542 9843 25594
rect 9895 25542 9907 25594
rect 9959 25542 9971 25594
rect 10023 25542 10035 25594
rect 10087 25542 19176 25594
rect 19228 25542 19240 25594
rect 19292 25542 19304 25594
rect 19356 25542 19368 25594
rect 19420 25542 26392 25594
rect 632 25520 26392 25542
rect 13136 25347 13194 25353
rect 13136 25313 13148 25347
rect 13182 25344 13194 25347
rect 13250 25344 13256 25356
rect 13182 25316 13256 25344
rect 13182 25313 13194 25316
rect 13136 25307 13194 25313
rect 13250 25304 13256 25316
rect 13308 25304 13314 25356
rect 20794 25353 20800 25356
rect 20772 25347 20800 25353
rect 20772 25313 20784 25347
rect 20772 25307 20800 25313
rect 20794 25304 20800 25307
rect 20852 25304 20858 25356
rect 13207 25143 13265 25149
rect 13207 25109 13219 25143
rect 13253 25140 13265 25143
rect 17114 25140 17120 25152
rect 13253 25112 17120 25140
rect 13253 25109 13265 25112
rect 13207 25103 13265 25109
rect 17114 25100 17120 25112
rect 17172 25100 17178 25152
rect 20843 25143 20901 25149
rect 20843 25109 20855 25143
rect 20889 25140 20901 25143
rect 21990 25140 21996 25152
rect 20889 25112 21996 25140
rect 20889 25109 20901 25112
rect 20843 25103 20901 25109
rect 21990 25100 21996 25112
rect 22048 25100 22054 25152
rect 632 25050 26392 25072
rect 632 24998 5176 25050
rect 5228 24998 5240 25050
rect 5292 24998 5304 25050
rect 5356 24998 5368 25050
rect 5420 24998 14510 25050
rect 14562 24998 14574 25050
rect 14626 24998 14638 25050
rect 14690 24998 14702 25050
rect 14754 24998 23843 25050
rect 23895 24998 23907 25050
rect 23959 24998 23971 25050
rect 24023 24998 24035 25050
rect 24087 24998 26392 25050
rect 632 24976 26392 24998
rect 13161 24939 13219 24945
rect 13161 24905 13173 24939
rect 13207 24936 13219 24939
rect 13250 24936 13256 24948
rect 13207 24908 13256 24936
rect 13207 24905 13219 24908
rect 13161 24899 13219 24905
rect 13250 24896 13256 24908
rect 13308 24896 13314 24948
rect 20794 24936 20800 24948
rect 20755 24908 20800 24936
rect 20794 24896 20800 24908
rect 20852 24896 20858 24948
rect 11318 24800 11324 24812
rect 11279 24772 11324 24800
rect 11318 24760 11324 24772
rect 11376 24760 11382 24812
rect 24290 24800 24296 24812
rect 24251 24772 24296 24800
rect 24290 24760 24296 24772
rect 24348 24760 24354 24812
rect 25394 24800 25400 24812
rect 25355 24772 25400 24800
rect 25394 24760 25400 24772
rect 25452 24760 25458 24812
rect 10928 24735 10986 24741
rect 10928 24701 10940 24735
rect 10974 24732 10986 24735
rect 11336 24732 11364 24760
rect 10974 24704 11364 24732
rect 10974 24701 10986 24704
rect 10928 24695 10986 24701
rect 12606 24692 12612 24744
rect 12664 24741 12670 24744
rect 12664 24735 12702 24741
rect 12690 24732 12702 24735
rect 13437 24735 13495 24741
rect 13437 24732 13449 24735
rect 12690 24704 13449 24732
rect 12690 24701 12702 24704
rect 12664 24695 12702 24701
rect 13437 24701 13449 24704
rect 13483 24701 13495 24735
rect 13437 24695 13495 24701
rect 12664 24692 12670 24695
rect 14078 24692 14084 24744
rect 14136 24732 14142 24744
rect 15458 24741 15464 24744
rect 14265 24735 14323 24741
rect 14265 24732 14277 24735
rect 14136 24704 14277 24732
rect 14136 24692 14142 24704
rect 14265 24701 14277 24704
rect 14311 24732 14323 24735
rect 14817 24735 14875 24741
rect 14817 24732 14829 24735
rect 14311 24704 14829 24732
rect 14311 24701 14323 24704
rect 14265 24695 14323 24701
rect 14817 24701 14829 24704
rect 14863 24701 14875 24735
rect 14817 24695 14875 24701
rect 15436 24735 15464 24741
rect 15436 24701 15448 24735
rect 15516 24732 15522 24744
rect 15829 24735 15887 24741
rect 15829 24732 15841 24735
rect 15516 24704 15841 24732
rect 15436 24695 15464 24701
rect 15458 24692 15464 24695
rect 15516 24692 15522 24704
rect 15829 24701 15841 24704
rect 15875 24701 15887 24735
rect 15829 24695 15887 24701
rect 19693 24735 19751 24741
rect 19693 24701 19705 24735
rect 19739 24732 19751 24735
rect 20150 24732 20156 24744
rect 19739 24704 20156 24732
rect 19739 24701 19751 24704
rect 19693 24695 19751 24701
rect 20150 24692 20156 24704
rect 20208 24692 20214 24744
rect 21346 24692 21352 24744
rect 21404 24732 21410 24744
rect 21476 24735 21534 24741
rect 21476 24732 21488 24735
rect 21404 24704 21488 24732
rect 21404 24692 21410 24704
rect 21476 24701 21488 24704
rect 21522 24732 21534 24735
rect 21901 24735 21959 24741
rect 21901 24732 21913 24735
rect 21522 24704 21913 24732
rect 21522 24701 21534 24704
rect 21476 24695 21534 24701
rect 21901 24701 21913 24704
rect 21947 24701 21959 24735
rect 21901 24695 21959 24701
rect 23900 24735 23958 24741
rect 23900 24701 23912 24735
rect 23946 24732 23958 24735
rect 24308 24732 24336 24760
rect 23946 24704 24336 24732
rect 24912 24735 24970 24741
rect 23946 24701 23958 24704
rect 23900 24695 23958 24701
rect 24912 24701 24924 24735
rect 24958 24732 24970 24735
rect 25412 24732 25440 24760
rect 24958 24704 25440 24732
rect 24958 24701 24970 24704
rect 24912 24695 24970 24701
rect 12747 24667 12805 24673
rect 12747 24633 12759 24667
rect 12793 24664 12805 24667
rect 14170 24664 14176 24676
rect 12793 24636 14176 24664
rect 12793 24633 12805 24636
rect 12747 24627 12805 24633
rect 14170 24624 14176 24636
rect 14228 24624 14234 24676
rect 20518 24664 20524 24676
rect 20479 24636 20524 24664
rect 20518 24624 20524 24636
rect 20576 24624 20582 24676
rect 11042 24605 11048 24608
rect 10999 24599 11048 24605
rect 10999 24565 11011 24599
rect 11045 24565 11048 24599
rect 10999 24559 11048 24565
rect 11042 24556 11048 24559
rect 11100 24556 11106 24608
rect 14446 24596 14452 24608
rect 14407 24568 14452 24596
rect 14446 24556 14452 24568
rect 14504 24556 14510 24608
rect 15507 24599 15565 24605
rect 15507 24565 15519 24599
rect 15553 24596 15565 24599
rect 16010 24596 16016 24608
rect 15553 24568 16016 24596
rect 15553 24565 15565 24568
rect 15507 24559 15565 24565
rect 16010 24556 16016 24568
rect 16068 24556 16074 24608
rect 17669 24599 17727 24605
rect 17669 24565 17681 24599
rect 17715 24596 17727 24599
rect 18034 24596 18040 24608
rect 17715 24568 18040 24596
rect 17715 24565 17727 24568
rect 17669 24559 17727 24565
rect 18034 24556 18040 24568
rect 18092 24556 18098 24608
rect 21579 24599 21637 24605
rect 21579 24565 21591 24599
rect 21625 24596 21637 24599
rect 21806 24596 21812 24608
rect 21625 24568 21812 24596
rect 21625 24565 21637 24568
rect 21579 24559 21637 24565
rect 21806 24556 21812 24568
rect 21864 24556 21870 24608
rect 23971 24599 24029 24605
rect 23971 24565 23983 24599
rect 24017 24596 24029 24599
rect 24198 24596 24204 24608
rect 24017 24568 24204 24596
rect 24017 24565 24029 24568
rect 23971 24559 24029 24565
rect 24198 24556 24204 24568
rect 24256 24556 24262 24608
rect 25026 24605 25032 24608
rect 24983 24599 25032 24605
rect 24983 24565 24995 24599
rect 25029 24565 25032 24599
rect 24983 24559 25032 24565
rect 25026 24556 25032 24559
rect 25084 24556 25090 24608
rect 632 24506 26392 24528
rect 632 24454 9843 24506
rect 9895 24454 9907 24506
rect 9959 24454 9971 24506
rect 10023 24454 10035 24506
rect 10087 24454 19176 24506
rect 19228 24454 19240 24506
rect 19292 24454 19304 24506
rect 19356 24454 19368 24506
rect 19420 24454 26392 24506
rect 632 24432 26392 24454
rect 14998 24392 15004 24404
rect 14959 24364 15004 24392
rect 14998 24352 15004 24364
rect 15056 24352 15062 24404
rect 18494 24392 18500 24404
rect 18455 24364 18500 24392
rect 18494 24352 18500 24364
rect 18552 24352 18558 24404
rect 22266 24392 22272 24404
rect 22227 24364 22272 24392
rect 22266 24352 22272 24364
rect 22324 24352 22330 24404
rect 23557 24395 23615 24401
rect 23557 24361 23569 24395
rect 23603 24392 23615 24395
rect 24842 24392 24848 24404
rect 23603 24364 24848 24392
rect 23603 24361 23615 24364
rect 23557 24355 23615 24361
rect 24842 24352 24848 24364
rect 24900 24352 24906 24404
rect 20518 24284 20524 24336
rect 20576 24324 20582 24336
rect 20613 24327 20671 24333
rect 20613 24324 20625 24327
rect 20576 24296 20625 24324
rect 20576 24284 20582 24296
rect 20613 24293 20625 24296
rect 20659 24293 20671 24327
rect 20613 24287 20671 24293
rect 5960 24259 6018 24265
rect 5960 24225 5972 24259
rect 6006 24256 6018 24259
rect 6166 24256 6172 24268
rect 6006 24228 6172 24256
rect 6006 24225 6018 24228
rect 5960 24219 6018 24225
rect 6166 24216 6172 24228
rect 6224 24216 6230 24268
rect 8076 24259 8134 24265
rect 8076 24225 8088 24259
rect 8122 24256 8134 24259
rect 8282 24256 8288 24268
rect 8122 24228 8288 24256
rect 8122 24225 8134 24228
rect 8076 24219 8134 24225
rect 8282 24216 8288 24228
rect 8340 24216 8346 24268
rect 9294 24265 9300 24268
rect 9272 24259 9300 24265
rect 9272 24225 9284 24259
rect 9272 24219 9300 24225
rect 9294 24216 9300 24219
rect 9352 24216 9358 24268
rect 12793 24259 12851 24265
rect 12793 24225 12805 24259
rect 12839 24256 12851 24259
rect 12882 24256 12888 24268
rect 12839 24228 12888 24256
rect 12839 24225 12851 24228
rect 12793 24219 12851 24225
rect 12882 24216 12888 24228
rect 12940 24216 12946 24268
rect 13802 24265 13808 24268
rect 13780 24259 13808 24265
rect 13780 24256 13792 24259
rect 13715 24228 13792 24256
rect 13780 24225 13792 24228
rect 13860 24256 13866 24268
rect 14354 24256 14360 24268
rect 13860 24228 14360 24256
rect 13780 24219 13808 24225
rect 13802 24216 13808 24219
rect 13860 24216 13866 24228
rect 14354 24216 14360 24228
rect 14412 24216 14418 24268
rect 14817 24259 14875 24265
rect 14817 24225 14829 24259
rect 14863 24225 14875 24259
rect 14817 24219 14875 24225
rect 11137 24191 11195 24197
rect 11137 24157 11149 24191
rect 11183 24188 11195 24191
rect 11686 24188 11692 24200
rect 11183 24160 11692 24188
rect 11183 24157 11195 24160
rect 11137 24151 11195 24157
rect 11686 24148 11692 24160
rect 11744 24148 11750 24200
rect 12146 24188 12152 24200
rect 12107 24160 12152 24188
rect 12146 24148 12152 24160
rect 12204 24148 12210 24200
rect 14170 24148 14176 24200
rect 14228 24188 14234 24200
rect 14832 24188 14860 24219
rect 16746 24216 16752 24268
rect 16804 24256 16810 24268
rect 16841 24259 16899 24265
rect 16841 24256 16853 24259
rect 16804 24228 16853 24256
rect 16804 24216 16810 24228
rect 16841 24225 16853 24228
rect 16887 24225 16899 24259
rect 18310 24256 18316 24268
rect 18271 24228 18316 24256
rect 16841 24219 16899 24225
rect 18310 24216 18316 24228
rect 18368 24216 18374 24268
rect 21806 24216 21812 24268
rect 21864 24256 21870 24268
rect 22085 24259 22143 24265
rect 22085 24256 22097 24259
rect 21864 24228 22097 24256
rect 21864 24216 21870 24228
rect 22085 24225 22097 24228
rect 22131 24225 22143 24259
rect 22085 24219 22143 24225
rect 22634 24216 22640 24268
rect 22692 24256 22698 24268
rect 23373 24259 23431 24265
rect 23373 24256 23385 24259
rect 22692 24228 23385 24256
rect 22692 24216 22698 24228
rect 23373 24225 23385 24228
rect 23419 24256 23431 24259
rect 24290 24256 24296 24268
rect 23419 24228 24296 24256
rect 23419 24225 23431 24228
rect 23373 24219 23431 24225
rect 24290 24216 24296 24228
rect 24348 24216 24354 24268
rect 24566 24265 24572 24268
rect 24544 24259 24572 24265
rect 24544 24225 24556 24259
rect 24544 24219 24572 24225
rect 24566 24216 24572 24219
rect 24624 24216 24630 24268
rect 14228 24160 14860 24188
rect 20521 24191 20579 24197
rect 14228 24148 14234 24160
rect 20521 24157 20533 24191
rect 20567 24188 20579 24191
rect 20610 24188 20616 24200
rect 20567 24160 20616 24188
rect 20567 24157 20579 24160
rect 20521 24151 20579 24157
rect 20610 24148 20616 24160
rect 20668 24148 20674 24200
rect 20797 24191 20855 24197
rect 20797 24157 20809 24191
rect 20843 24157 20855 24191
rect 20797 24151 20855 24157
rect 20812 24064 20840 24151
rect 24474 24080 24480 24132
rect 24532 24120 24538 24132
rect 24615 24123 24673 24129
rect 24615 24120 24627 24123
rect 24532 24092 24627 24120
rect 24532 24080 24538 24092
rect 24615 24089 24627 24092
rect 24661 24089 24673 24123
rect 24615 24083 24673 24089
rect 6031 24055 6089 24061
rect 6031 24021 6043 24055
rect 6077 24052 6089 24055
rect 6258 24052 6264 24064
rect 6077 24024 6264 24052
rect 6077 24021 6089 24024
rect 6031 24015 6089 24021
rect 6258 24012 6264 24024
rect 6316 24012 6322 24064
rect 8190 24061 8196 24064
rect 8147 24055 8196 24061
rect 8147 24021 8159 24055
rect 8193 24021 8196 24055
rect 8147 24015 8196 24021
rect 8190 24012 8196 24015
rect 8248 24012 8254 24064
rect 9386 24061 9392 24064
rect 9343 24055 9392 24061
rect 9343 24021 9355 24055
rect 9389 24021 9392 24055
rect 9343 24015 9392 24021
rect 9386 24012 9392 24015
rect 9444 24012 9450 24064
rect 13851 24055 13909 24061
rect 13851 24021 13863 24055
rect 13897 24052 13909 24055
rect 14262 24052 14268 24064
rect 13897 24024 14268 24052
rect 13897 24021 13909 24024
rect 13851 24015 13909 24021
rect 14262 24012 14268 24024
rect 14320 24012 14326 24064
rect 17206 24052 17212 24064
rect 17167 24024 17212 24052
rect 17206 24012 17212 24024
rect 17264 24012 17270 24064
rect 17758 24052 17764 24064
rect 17719 24024 17764 24052
rect 17758 24012 17764 24024
rect 17816 24012 17822 24064
rect 20794 24012 20800 24064
rect 20852 24012 20858 24064
rect 632 23962 26392 23984
rect 632 23910 5176 23962
rect 5228 23910 5240 23962
rect 5292 23910 5304 23962
rect 5356 23910 5368 23962
rect 5420 23910 14510 23962
rect 14562 23910 14574 23962
rect 14626 23910 14638 23962
rect 14690 23910 14702 23962
rect 14754 23910 23843 23962
rect 23895 23910 23907 23962
rect 23959 23910 23971 23962
rect 24023 23910 24035 23962
rect 24087 23910 26392 23962
rect 632 23888 26392 23910
rect 1934 23857 1940 23860
rect 1891 23851 1940 23857
rect 1891 23817 1903 23851
rect 1937 23817 1940 23851
rect 1891 23811 1940 23817
rect 1934 23808 1940 23811
rect 1992 23808 1998 23860
rect 2026 23808 2032 23860
rect 2084 23848 2090 23860
rect 2213 23851 2271 23857
rect 2213 23848 2225 23851
rect 2084 23820 2225 23848
rect 2084 23808 2090 23820
rect 2213 23817 2225 23820
rect 2259 23817 2271 23851
rect 2213 23811 2271 23817
rect 3038 23808 3044 23860
rect 3096 23848 3102 23860
rect 3225 23851 3283 23857
rect 3225 23848 3237 23851
rect 3096 23820 3237 23848
rect 3096 23808 3102 23820
rect 3225 23817 3237 23820
rect 3271 23817 3283 23851
rect 3225 23811 3283 23817
rect 5062 23808 5068 23860
rect 5120 23848 5126 23860
rect 5341 23851 5399 23857
rect 5341 23848 5353 23851
rect 5120 23820 5353 23848
rect 5120 23808 5126 23820
rect 5341 23817 5353 23820
rect 5387 23817 5399 23851
rect 5341 23811 5399 23817
rect 5985 23851 6043 23857
rect 5985 23817 5997 23851
rect 6031 23848 6043 23851
rect 6166 23848 6172 23860
rect 6031 23820 6172 23848
rect 6031 23817 6043 23820
rect 5985 23811 6043 23817
rect 6166 23808 6172 23820
rect 6224 23808 6230 23860
rect 7178 23808 7184 23860
rect 7236 23848 7242 23860
rect 7365 23851 7423 23857
rect 7365 23848 7377 23851
rect 7236 23820 7377 23848
rect 7236 23808 7242 23820
rect 7365 23817 7377 23820
rect 7411 23817 7423 23851
rect 8374 23848 8380 23860
rect 8335 23820 8380 23848
rect 7365 23811 7423 23817
rect 8374 23808 8380 23820
rect 8432 23808 8438 23860
rect 9294 23848 9300 23860
rect 9255 23820 9300 23848
rect 9294 23808 9300 23820
rect 9352 23808 9358 23860
rect 10306 23848 10312 23860
rect 10267 23820 10312 23848
rect 10306 23808 10312 23820
rect 10364 23808 10370 23860
rect 10950 23848 10956 23860
rect 10911 23820 10956 23848
rect 10950 23808 10956 23820
rect 11008 23808 11014 23860
rect 11686 23848 11692 23860
rect 11647 23820 11692 23848
rect 11686 23808 11692 23820
rect 11744 23808 11750 23860
rect 12146 23848 12152 23860
rect 12107 23820 12152 23848
rect 12146 23808 12152 23820
rect 12204 23808 12210 23860
rect 13802 23848 13808 23860
rect 13763 23820 13808 23848
rect 13802 23808 13808 23820
rect 13860 23808 13866 23860
rect 14078 23857 14084 23860
rect 14035 23851 14084 23857
rect 14035 23817 14047 23851
rect 14081 23817 14084 23851
rect 14035 23811 14084 23817
rect 14078 23808 14084 23811
rect 14136 23808 14142 23860
rect 14170 23808 14176 23860
rect 14228 23848 14234 23860
rect 14357 23851 14415 23857
rect 14357 23848 14369 23851
rect 14228 23820 14369 23848
rect 14228 23808 14234 23820
rect 14357 23817 14369 23820
rect 14403 23817 14415 23851
rect 19690 23848 19696 23860
rect 19651 23820 19696 23848
rect 14357 23811 14415 23817
rect 19690 23808 19696 23820
rect 19748 23808 19754 23860
rect 20518 23848 20524 23860
rect 20479 23820 20524 23848
rect 20518 23808 20524 23820
rect 20576 23808 20582 23860
rect 21806 23808 21812 23860
rect 21864 23848 21870 23860
rect 22085 23851 22143 23857
rect 22085 23848 22097 23851
rect 21864 23820 22097 23848
rect 21864 23808 21870 23820
rect 22085 23817 22097 23820
rect 22131 23817 22143 23851
rect 22634 23848 22640 23860
rect 22595 23820 22640 23848
rect 22085 23811 22143 23817
rect 22634 23808 22640 23820
rect 22692 23808 22698 23860
rect 24566 23848 24572 23860
rect 24527 23820 24572 23848
rect 24566 23808 24572 23820
rect 24624 23808 24630 23860
rect 25302 23848 25308 23860
rect 25263 23820 25308 23848
rect 25302 23808 25308 23820
rect 25360 23808 25366 23860
rect 8101 23783 8159 23789
rect 8101 23749 8113 23783
rect 8147 23780 8159 23783
rect 8282 23780 8288 23792
rect 8147 23752 8288 23780
rect 8147 23749 8159 23752
rect 8101 23743 8159 23749
rect 8282 23740 8288 23752
rect 8340 23740 8346 23792
rect 11704 23712 11732 23808
rect 16611 23783 16669 23789
rect 16611 23749 16623 23783
rect 16657 23780 16669 23783
rect 18310 23780 18316 23792
rect 16657 23752 18316 23780
rect 16657 23749 16669 23752
rect 16611 23743 16669 23749
rect 18310 23740 18316 23752
rect 18368 23780 18374 23792
rect 18681 23783 18739 23789
rect 18681 23780 18693 23783
rect 18368 23752 18693 23780
rect 18368 23740 18374 23752
rect 18681 23749 18693 23752
rect 18727 23749 18739 23783
rect 18681 23743 18739 23749
rect 12425 23715 12483 23721
rect 12425 23712 12437 23715
rect 11704 23684 12437 23712
rect 12425 23681 12437 23684
rect 12471 23681 12483 23715
rect 12425 23675 12483 23681
rect 20705 23715 20763 23721
rect 20705 23681 20717 23715
rect 20751 23712 20763 23715
rect 20794 23712 20800 23724
rect 20751 23684 20800 23712
rect 20751 23681 20763 23684
rect 20705 23675 20763 23681
rect 20794 23672 20800 23684
rect 20852 23712 20858 23724
rect 21625 23715 21683 23721
rect 21625 23712 21637 23715
rect 20852 23684 21637 23712
rect 20852 23672 20858 23684
rect 21625 23681 21637 23684
rect 21671 23681 21683 23715
rect 21625 23675 21683 23681
rect 1820 23647 1878 23653
rect 1820 23613 1832 23647
rect 1866 23644 1878 23647
rect 2026 23644 2032 23656
rect 1866 23616 2032 23644
rect 1866 23613 1878 23616
rect 1820 23607 1878 23613
rect 2026 23604 2032 23616
rect 2084 23604 2090 23656
rect 2832 23647 2890 23653
rect 2832 23613 2844 23647
rect 2878 23644 2890 23647
rect 3038 23644 3044 23656
rect 2878 23616 3044 23644
rect 2878 23613 2890 23616
rect 2832 23607 2890 23613
rect 3038 23604 3044 23616
rect 3096 23604 3102 23656
rect 4948 23647 5006 23653
rect 4948 23613 4960 23647
rect 4994 23644 5006 23647
rect 5062 23644 5068 23656
rect 4994 23616 5068 23644
rect 4994 23613 5006 23616
rect 4948 23607 5006 23613
rect 5062 23604 5068 23616
rect 5120 23604 5126 23656
rect 6972 23647 7030 23653
rect 6972 23613 6984 23647
rect 7018 23644 7030 23647
rect 7178 23644 7184 23656
rect 7018 23616 7184 23644
rect 7018 23613 7030 23616
rect 6972 23607 7030 23613
rect 7178 23604 7184 23616
rect 7236 23604 7242 23656
rect 8374 23604 8380 23656
rect 8432 23644 8438 23656
rect 8596 23647 8654 23653
rect 8596 23644 8608 23647
rect 8432 23616 8608 23644
rect 8432 23604 8438 23616
rect 8596 23613 8608 23616
rect 8642 23613 8654 23647
rect 8596 23607 8654 23613
rect 9824 23647 9882 23653
rect 9824 23613 9836 23647
rect 9870 23644 9882 23647
rect 10306 23644 10312 23656
rect 9870 23616 10312 23644
rect 9870 23613 9882 23616
rect 9824 23607 9882 23613
rect 10306 23604 10312 23616
rect 10364 23604 10370 23656
rect 10769 23647 10827 23653
rect 10769 23613 10781 23647
rect 10815 23644 10827 23647
rect 10950 23644 10956 23656
rect 10815 23616 10956 23644
rect 10815 23613 10827 23616
rect 10769 23607 10827 23613
rect 10950 23604 10956 23616
rect 11008 23644 11014 23656
rect 11321 23647 11379 23653
rect 11321 23644 11333 23647
rect 11008 23616 11333 23644
rect 11008 23604 11014 23616
rect 11321 23613 11333 23616
rect 11367 23613 11379 23647
rect 13932 23647 13990 23653
rect 13932 23644 13944 23647
rect 11321 23607 11379 23613
rect 13084 23616 13944 23644
rect 13084 23588 13112 23616
rect 13932 23613 13944 23616
rect 13978 23613 13990 23647
rect 13932 23607 13990 23613
rect 15277 23647 15335 23653
rect 15277 23613 15289 23647
rect 15323 23644 15335 23647
rect 16508 23647 16566 23653
rect 16508 23644 16520 23647
rect 15323 23616 15357 23644
rect 16304 23616 16520 23644
rect 15323 23613 15335 23616
rect 15277 23607 15335 23613
rect 12146 23536 12152 23588
rect 12204 23576 12210 23588
rect 12517 23579 12575 23585
rect 12517 23576 12529 23579
rect 12204 23548 12529 23576
rect 12204 23536 12210 23548
rect 12517 23545 12529 23548
rect 12563 23545 12575 23579
rect 13066 23576 13072 23588
rect 13027 23548 13072 23576
rect 12517 23539 12575 23545
rect 13066 23536 13072 23548
rect 13124 23536 13130 23588
rect 14817 23579 14875 23585
rect 14817 23545 14829 23579
rect 14863 23576 14875 23579
rect 15292 23576 15320 23607
rect 15826 23576 15832 23588
rect 14863 23548 15832 23576
rect 14863 23545 14875 23548
rect 14817 23539 14875 23545
rect 15826 23536 15832 23548
rect 15884 23536 15890 23588
rect 16304 23520 16332 23616
rect 16508 23613 16520 23616
rect 16554 23613 16566 23647
rect 16508 23607 16566 23613
rect 19509 23647 19567 23653
rect 19509 23613 19521 23647
rect 19555 23613 19567 23647
rect 23002 23644 23008 23656
rect 22915 23616 23008 23644
rect 19509 23607 19567 23613
rect 17758 23576 17764 23588
rect 17719 23548 17764 23576
rect 17758 23536 17764 23548
rect 17816 23536 17822 23588
rect 17853 23579 17911 23585
rect 17853 23545 17865 23579
rect 17899 23545 17911 23579
rect 17853 23539 17911 23545
rect 18405 23579 18463 23585
rect 18405 23545 18417 23579
rect 18451 23576 18463 23579
rect 18494 23576 18500 23588
rect 18451 23548 18500 23576
rect 18451 23545 18463 23548
rect 18405 23539 18463 23545
rect 2903 23511 2961 23517
rect 2903 23477 2915 23511
rect 2949 23508 2961 23511
rect 3590 23508 3596 23520
rect 2949 23480 3596 23508
rect 2949 23477 2961 23480
rect 2903 23471 2961 23477
rect 3590 23468 3596 23480
rect 3648 23468 3654 23520
rect 4970 23468 4976 23520
rect 5028 23517 5034 23520
rect 5028 23511 5077 23517
rect 5028 23477 5031 23511
rect 5065 23477 5077 23511
rect 5028 23471 5077 23477
rect 7043 23511 7101 23517
rect 7043 23477 7055 23511
rect 7089 23508 7101 23511
rect 7730 23508 7736 23520
rect 7089 23480 7736 23508
rect 7089 23477 7101 23480
rect 7043 23471 7101 23477
rect 5028 23468 5034 23471
rect 7730 23468 7736 23480
rect 7788 23468 7794 23520
rect 8699 23511 8757 23517
rect 8699 23477 8711 23511
rect 8745 23508 8757 23511
rect 8926 23508 8932 23520
rect 8745 23480 8932 23508
rect 8745 23477 8757 23480
rect 8699 23471 8757 23477
rect 8926 23468 8932 23480
rect 8984 23468 8990 23520
rect 9895 23511 9953 23517
rect 9895 23477 9907 23511
rect 9941 23508 9953 23511
rect 10306 23508 10312 23520
rect 9941 23480 10312 23508
rect 9941 23477 9953 23480
rect 9895 23471 9953 23477
rect 10306 23468 10312 23480
rect 10364 23468 10370 23520
rect 15182 23508 15188 23520
rect 15143 23480 15188 23508
rect 15182 23468 15188 23480
rect 15240 23468 15246 23520
rect 16286 23508 16292 23520
rect 16247 23480 16292 23508
rect 16286 23468 16292 23480
rect 16344 23468 16350 23520
rect 16746 23468 16752 23520
rect 16804 23508 16810 23520
rect 16933 23511 16991 23517
rect 16933 23508 16945 23511
rect 16804 23480 16945 23508
rect 16804 23468 16810 23480
rect 16933 23477 16945 23480
rect 16979 23477 16991 23511
rect 17390 23508 17396 23520
rect 17303 23480 17396 23508
rect 16933 23471 16991 23477
rect 17390 23468 17396 23480
rect 17448 23508 17454 23520
rect 17868 23508 17896 23539
rect 18494 23536 18500 23548
rect 18552 23536 18558 23588
rect 19524 23520 19552 23607
rect 23002 23604 23008 23616
rect 23060 23644 23066 23656
rect 23281 23647 23339 23653
rect 23281 23644 23293 23647
rect 23060 23616 23293 23644
rect 23060 23604 23066 23616
rect 23281 23613 23293 23616
rect 23327 23613 23339 23647
rect 23281 23607 23339 23613
rect 24820 23647 24878 23653
rect 24820 23613 24832 23647
rect 24866 23644 24878 23647
rect 25302 23644 25308 23656
rect 24866 23616 25308 23644
rect 24866 23613 24878 23616
rect 24820 23607 24878 23613
rect 25302 23604 25308 23616
rect 25360 23604 25366 23656
rect 20797 23579 20855 23585
rect 20797 23545 20809 23579
rect 20843 23545 20855 23579
rect 21346 23576 21352 23588
rect 21307 23548 21352 23576
rect 20797 23539 20855 23545
rect 17448 23480 17896 23508
rect 19417 23511 19475 23517
rect 17448 23468 17454 23480
rect 19417 23477 19429 23511
rect 19463 23508 19475 23511
rect 19506 23508 19512 23520
rect 19463 23480 19512 23508
rect 19463 23477 19475 23480
rect 19417 23471 19475 23477
rect 19506 23468 19512 23480
rect 19564 23468 19570 23520
rect 20150 23508 20156 23520
rect 20111 23480 20156 23508
rect 20150 23468 20156 23480
rect 20208 23508 20214 23520
rect 20812 23508 20840 23539
rect 21346 23536 21352 23548
rect 21404 23536 21410 23588
rect 23186 23576 23192 23588
rect 23147 23548 23192 23576
rect 23186 23536 23192 23548
rect 23244 23536 23250 23588
rect 20208 23480 20840 23508
rect 20208 23468 20214 23480
rect 24474 23468 24480 23520
rect 24532 23508 24538 23520
rect 24891 23511 24949 23517
rect 24891 23508 24903 23511
rect 24532 23480 24903 23508
rect 24532 23468 24538 23480
rect 24891 23477 24903 23480
rect 24937 23477 24949 23511
rect 24891 23471 24949 23477
rect 632 23418 26392 23440
rect 632 23366 9843 23418
rect 9895 23366 9907 23418
rect 9959 23366 9971 23418
rect 10023 23366 10035 23418
rect 10087 23366 19176 23418
rect 19228 23366 19240 23418
rect 19292 23366 19304 23418
rect 19356 23366 19368 23418
rect 19420 23366 26392 23418
rect 632 23344 26392 23366
rect 20610 23264 20616 23316
rect 20668 23304 20674 23316
rect 20981 23307 21039 23313
rect 20981 23304 20993 23307
rect 20668 23276 20993 23304
rect 20668 23264 20674 23276
rect 20981 23273 20993 23276
rect 21027 23273 21039 23307
rect 20981 23267 21039 23273
rect 22910 23264 22916 23316
rect 22968 23264 22974 23316
rect 24198 23304 24204 23316
rect 23020 23276 24204 23304
rect 10858 23236 10864 23248
rect 10819 23208 10864 23236
rect 10858 23196 10864 23208
rect 10916 23196 10922 23248
rect 10953 23239 11011 23245
rect 10953 23205 10965 23239
rect 10999 23236 11011 23239
rect 11318 23236 11324 23248
rect 10999 23208 11324 23236
rect 10999 23205 11011 23208
rect 10953 23199 11011 23205
rect 11318 23196 11324 23208
rect 11376 23196 11382 23248
rect 12241 23239 12299 23245
rect 12241 23205 12253 23239
rect 12287 23236 12299 23239
rect 12517 23239 12575 23245
rect 12517 23236 12529 23239
rect 12287 23208 12529 23236
rect 12287 23205 12299 23208
rect 12241 23199 12299 23205
rect 12517 23205 12529 23208
rect 12563 23236 12575 23239
rect 12882 23236 12888 23248
rect 12563 23208 12888 23236
rect 12563 23205 12575 23208
rect 12517 23199 12575 23205
rect 12882 23196 12888 23208
rect 12940 23196 12946 23248
rect 13066 23236 13072 23248
rect 13027 23208 13072 23236
rect 13066 23196 13072 23208
rect 13124 23236 13130 23248
rect 13897 23239 13955 23245
rect 13897 23236 13909 23239
rect 13124 23208 13909 23236
rect 13124 23196 13130 23208
rect 13897 23205 13909 23208
rect 13943 23205 13955 23239
rect 15182 23236 15188 23248
rect 15143 23208 15188 23236
rect 13897 23199 13955 23205
rect 15182 23196 15188 23208
rect 15240 23196 15246 23248
rect 16746 23236 16752 23248
rect 16707 23208 16752 23236
rect 16746 23196 16752 23208
rect 16804 23196 16810 23248
rect 18218 23196 18224 23248
rect 18276 23236 18282 23248
rect 18313 23239 18371 23245
rect 18313 23236 18325 23239
rect 18276 23208 18325 23236
rect 18276 23196 18282 23208
rect 18313 23205 18325 23208
rect 18359 23205 18371 23239
rect 21438 23236 21444 23248
rect 21399 23208 21444 23236
rect 18313 23199 18371 23205
rect 21438 23196 21444 23208
rect 21496 23196 21502 23248
rect 21533 23239 21591 23245
rect 21533 23205 21545 23239
rect 21579 23236 21591 23239
rect 21622 23236 21628 23248
rect 21579 23208 21628 23236
rect 21579 23205 21591 23208
rect 21533 23199 21591 23205
rect 21622 23196 21628 23208
rect 21680 23236 21686 23248
rect 22928 23236 22956 23264
rect 23020 23245 23048 23276
rect 24198 23264 24204 23276
rect 24256 23264 24262 23316
rect 24382 23264 24388 23316
rect 24440 23304 24446 23316
rect 24615 23307 24673 23313
rect 24615 23304 24627 23307
rect 24440 23276 24627 23304
rect 24440 23264 24446 23276
rect 24615 23273 24627 23276
rect 24661 23273 24673 23307
rect 24615 23267 24673 23273
rect 21680 23208 22956 23236
rect 23005 23239 23063 23245
rect 21680 23196 21686 23208
rect 23005 23205 23017 23239
rect 23051 23205 23063 23239
rect 23005 23199 23063 23205
rect 23097 23239 23155 23245
rect 23097 23205 23109 23239
rect 23143 23236 23155 23239
rect 23186 23236 23192 23248
rect 23143 23208 23192 23236
rect 23143 23205 23155 23208
rect 23097 23199 23155 23205
rect 23186 23196 23192 23208
rect 23244 23196 23250 23248
rect 9846 23168 9852 23180
rect 9807 23140 9852 23168
rect 9846 23128 9852 23140
rect 9904 23128 9910 23180
rect 24566 23177 24572 23180
rect 24544 23171 24572 23177
rect 24544 23137 24556 23171
rect 24544 23131 24572 23137
rect 24566 23128 24572 23131
rect 24624 23128 24630 23180
rect 9202 23100 9208 23112
rect 9163 23072 9208 23100
rect 9202 23060 9208 23072
rect 9260 23060 9266 23112
rect 11505 23103 11563 23109
rect 11505 23069 11517 23103
rect 11551 23100 11563 23103
rect 12422 23100 12428 23112
rect 11551 23072 12428 23100
rect 11551 23069 11563 23072
rect 11505 23063 11563 23069
rect 12422 23060 12428 23072
rect 12480 23060 12486 23112
rect 15090 23100 15096 23112
rect 15051 23072 15096 23100
rect 15090 23060 15096 23072
rect 15148 23060 15154 23112
rect 15737 23103 15795 23109
rect 15737 23069 15749 23103
rect 15783 23100 15795 23103
rect 15918 23100 15924 23112
rect 15783 23072 15924 23100
rect 15783 23069 15795 23072
rect 15737 23063 15795 23069
rect 15918 23060 15924 23072
rect 15976 23100 15982 23112
rect 16286 23100 16292 23112
rect 15976 23072 16292 23100
rect 15976 23060 15982 23072
rect 16286 23060 16292 23072
rect 16344 23060 16350 23112
rect 16654 23100 16660 23112
rect 16615 23072 16660 23100
rect 16654 23060 16660 23072
rect 16712 23060 16718 23112
rect 17298 23100 17304 23112
rect 17259 23072 17304 23100
rect 17298 23060 17304 23072
rect 17356 23100 17362 23112
rect 17758 23100 17764 23112
rect 17356 23072 17764 23100
rect 17356 23060 17362 23072
rect 17758 23060 17764 23072
rect 17816 23060 17822 23112
rect 18034 23060 18040 23112
rect 18092 23100 18098 23112
rect 18221 23103 18279 23109
rect 18221 23100 18233 23103
rect 18092 23072 18233 23100
rect 18092 23060 18098 23072
rect 18221 23069 18233 23072
rect 18267 23069 18279 23103
rect 18494 23100 18500 23112
rect 18455 23072 18500 23100
rect 18221 23063 18279 23069
rect 18494 23060 18500 23072
rect 18552 23060 18558 23112
rect 22085 23103 22143 23109
rect 22085 23069 22097 23103
rect 22131 23100 22143 23103
rect 23278 23100 23284 23112
rect 22131 23072 23284 23100
rect 22131 23069 22143 23072
rect 22085 23063 22143 23069
rect 23278 23060 23284 23072
rect 23336 23060 23342 23112
rect 17666 23032 17672 23044
rect 17627 23004 17672 23032
rect 17666 22992 17672 23004
rect 17724 22992 17730 23044
rect 15642 22924 15648 22976
rect 15700 22964 15706 22976
rect 16013 22967 16071 22973
rect 16013 22964 16025 22967
rect 15700 22936 16025 22964
rect 15700 22924 15706 22936
rect 16013 22933 16025 22936
rect 16059 22933 16071 22967
rect 20702 22964 20708 22976
rect 20663 22936 20708 22964
rect 16013 22927 16071 22933
rect 20702 22924 20708 22936
rect 20760 22924 20766 22976
rect 632 22874 26392 22896
rect 632 22822 5176 22874
rect 5228 22822 5240 22874
rect 5292 22822 5304 22874
rect 5356 22822 5368 22874
rect 5420 22822 14510 22874
rect 14562 22822 14574 22874
rect 14626 22822 14638 22874
rect 14690 22822 14702 22874
rect 14754 22822 23843 22874
rect 23895 22822 23907 22874
rect 23959 22822 23971 22874
rect 24023 22822 24035 22874
rect 24087 22822 26392 22874
rect 632 22800 26392 22822
rect 9202 22760 9208 22772
rect 9163 22732 9208 22760
rect 9202 22720 9208 22732
rect 9260 22720 9266 22772
rect 9570 22720 9576 22772
rect 9628 22760 9634 22772
rect 9846 22760 9852 22772
rect 9628 22732 9852 22760
rect 9628 22720 9634 22732
rect 9846 22720 9852 22732
rect 9904 22760 9910 22772
rect 10309 22763 10367 22769
rect 10309 22760 10321 22763
rect 9904 22732 10321 22760
rect 9904 22720 9910 22732
rect 10309 22729 10321 22732
rect 10355 22729 10367 22763
rect 10309 22723 10367 22729
rect 10950 22720 10956 22772
rect 11008 22769 11014 22772
rect 11008 22763 11057 22769
rect 11008 22729 11011 22763
rect 11045 22729 11057 22763
rect 11318 22760 11324 22772
rect 11279 22732 11324 22760
rect 11008 22723 11057 22729
rect 11008 22720 11014 22723
rect 11318 22720 11324 22732
rect 11376 22720 11382 22772
rect 15090 22720 15096 22772
rect 15148 22760 15154 22772
rect 15369 22763 15427 22769
rect 15369 22760 15381 22763
rect 15148 22732 15381 22760
rect 15148 22720 15154 22732
rect 15369 22729 15381 22732
rect 15415 22729 15427 22763
rect 15369 22723 15427 22729
rect 16654 22720 16660 22772
rect 16712 22760 16718 22772
rect 16933 22763 16991 22769
rect 16933 22760 16945 22763
rect 16712 22732 16945 22760
rect 16712 22720 16718 22732
rect 16933 22729 16945 22732
rect 16979 22729 16991 22763
rect 16933 22723 16991 22729
rect 17206 22720 17212 22772
rect 17264 22760 17270 22772
rect 17301 22763 17359 22769
rect 17301 22760 17313 22763
rect 17264 22732 17313 22760
rect 17264 22720 17270 22732
rect 17301 22729 17313 22732
rect 17347 22729 17359 22763
rect 17301 22723 17359 22729
rect 18034 22720 18040 22772
rect 18092 22760 18098 22772
rect 18957 22763 19015 22769
rect 18957 22760 18969 22763
rect 18092 22732 18969 22760
rect 18092 22720 18098 22732
rect 18957 22729 18969 22732
rect 19003 22729 19015 22763
rect 18957 22723 19015 22729
rect 19279 22763 19337 22769
rect 19279 22729 19291 22763
rect 19325 22760 19337 22763
rect 19506 22760 19512 22772
rect 19325 22732 19512 22760
rect 19325 22729 19337 22732
rect 19279 22723 19337 22729
rect 19506 22720 19512 22732
rect 19564 22720 19570 22772
rect 21622 22760 21628 22772
rect 21583 22732 21628 22760
rect 21622 22720 21628 22732
rect 21680 22720 21686 22772
rect 23005 22763 23063 22769
rect 23005 22729 23017 22763
rect 23051 22760 23063 22763
rect 23186 22760 23192 22772
rect 23051 22732 23192 22760
rect 23051 22729 23063 22732
rect 23005 22723 23063 22729
rect 23186 22720 23192 22732
rect 23244 22720 23250 22772
rect 24198 22760 24204 22772
rect 24159 22732 24204 22760
rect 24198 22720 24204 22732
rect 24256 22720 24262 22772
rect 21438 22652 21444 22704
rect 21496 22692 21502 22704
rect 21993 22695 22051 22701
rect 21993 22692 22005 22695
rect 21496 22664 22005 22692
rect 21496 22652 21502 22664
rect 21993 22661 22005 22664
rect 22039 22661 22051 22695
rect 21993 22655 22051 22661
rect 12422 22624 12428 22636
rect 12383 22596 12428 22624
rect 12422 22584 12428 22596
rect 12480 22624 12486 22636
rect 13345 22627 13403 22633
rect 13345 22624 13357 22627
rect 12480 22596 13357 22624
rect 12480 22584 12486 22596
rect 13345 22593 13357 22596
rect 13391 22593 13403 22627
rect 14078 22624 14084 22636
rect 14039 22596 14084 22624
rect 13345 22587 13403 22593
rect 14078 22584 14084 22596
rect 14136 22584 14142 22636
rect 15093 22627 15151 22633
rect 15093 22593 15105 22627
rect 15139 22624 15151 22627
rect 15182 22624 15188 22636
rect 15139 22596 15188 22624
rect 15139 22593 15151 22596
rect 15093 22587 15151 22593
rect 15182 22584 15188 22596
rect 15240 22584 15246 22636
rect 15642 22624 15648 22636
rect 15476 22596 15648 22624
rect 10896 22559 10954 22565
rect 10896 22556 10908 22559
rect 10692 22528 10908 22556
rect 8285 22491 8343 22497
rect 8285 22457 8297 22491
rect 8331 22488 8343 22491
rect 8837 22491 8895 22497
rect 8837 22488 8849 22491
rect 8331 22460 8849 22488
rect 8331 22457 8343 22460
rect 8285 22451 8343 22457
rect 8837 22457 8849 22460
rect 8883 22488 8895 22491
rect 9389 22491 9447 22497
rect 9389 22488 9401 22491
rect 8883 22460 9401 22488
rect 8883 22457 8895 22460
rect 8837 22451 8895 22457
rect 9389 22457 9401 22460
rect 9435 22457 9447 22491
rect 9389 22451 9447 22457
rect 9481 22491 9539 22497
rect 9481 22457 9493 22491
rect 9527 22457 9539 22491
rect 9481 22451 9539 22457
rect 10033 22491 10091 22497
rect 10033 22457 10045 22491
rect 10079 22488 10091 22491
rect 10214 22488 10220 22500
rect 10079 22460 10220 22488
rect 10079 22457 10091 22460
rect 10033 22451 10091 22457
rect 9202 22380 9208 22432
rect 9260 22420 9266 22432
rect 9496 22420 9524 22451
rect 10214 22448 10220 22460
rect 10272 22488 10278 22500
rect 10692 22497 10720 22528
rect 10896 22525 10908 22528
rect 10942 22525 10954 22559
rect 10896 22519 10954 22525
rect 14725 22559 14783 22565
rect 14725 22525 14737 22559
rect 14771 22556 14783 22559
rect 15476 22556 15504 22596
rect 15642 22584 15648 22596
rect 15700 22584 15706 22636
rect 15918 22624 15924 22636
rect 15879 22596 15924 22624
rect 15918 22584 15924 22596
rect 15976 22584 15982 22636
rect 17298 22584 17304 22636
rect 17356 22624 17362 22636
rect 17945 22627 18003 22633
rect 17945 22624 17957 22627
rect 17356 22596 17957 22624
rect 17356 22584 17362 22596
rect 17945 22593 17957 22596
rect 17991 22593 18003 22627
rect 21346 22624 21352 22636
rect 21307 22596 21352 22624
rect 17945 22587 18003 22593
rect 21346 22584 21352 22596
rect 21404 22584 21410 22636
rect 23278 22624 23284 22636
rect 23239 22596 23284 22624
rect 23278 22584 23284 22596
rect 23336 22584 23342 22636
rect 23554 22624 23560 22636
rect 23515 22596 23560 22624
rect 23554 22584 23560 22596
rect 23612 22624 23618 22636
rect 24566 22624 24572 22636
rect 23612 22596 24572 22624
rect 23612 22584 23618 22596
rect 24566 22584 24572 22596
rect 24624 22584 24630 22636
rect 14771 22528 15504 22556
rect 14771 22525 14783 22528
rect 14725 22519 14783 22525
rect 18494 22516 18500 22568
rect 18552 22556 18558 22568
rect 19176 22559 19234 22565
rect 19176 22556 19188 22559
rect 18552 22528 19188 22556
rect 18552 22516 18558 22528
rect 19176 22525 19188 22528
rect 19222 22556 19234 22559
rect 19601 22559 19659 22565
rect 19601 22556 19613 22559
rect 19222 22528 19613 22556
rect 19222 22525 19234 22528
rect 19176 22519 19234 22525
rect 19601 22525 19613 22528
rect 19647 22525 19659 22559
rect 19601 22519 19659 22525
rect 10677 22491 10735 22497
rect 10677 22488 10689 22491
rect 10272 22460 10689 22488
rect 10272 22448 10278 22460
rect 10677 22457 10689 22460
rect 10723 22457 10735 22491
rect 12054 22488 12060 22500
rect 12015 22460 12060 22488
rect 10677 22451 10735 22457
rect 12054 22448 12060 22460
rect 12112 22448 12118 22500
rect 12149 22491 12207 22497
rect 12149 22457 12161 22491
rect 12195 22457 12207 22491
rect 12149 22451 12207 22457
rect 14173 22491 14231 22497
rect 14173 22457 14185 22491
rect 14219 22457 14231 22491
rect 14173 22451 14231 22457
rect 15737 22491 15795 22497
rect 15737 22457 15749 22491
rect 15783 22488 15795 22491
rect 15826 22488 15832 22500
rect 15783 22460 15832 22488
rect 15783 22457 15795 22460
rect 15737 22451 15795 22457
rect 9260 22392 9524 22420
rect 11781 22423 11839 22429
rect 9260 22380 9266 22392
rect 11781 22389 11793 22423
rect 11827 22420 11839 22423
rect 11870 22420 11876 22432
rect 11827 22392 11876 22420
rect 11827 22389 11839 22392
rect 11781 22383 11839 22389
rect 11870 22380 11876 22392
rect 11928 22420 11934 22432
rect 12164 22420 12192 22451
rect 11928 22392 12192 22420
rect 11928 22380 11934 22392
rect 12882 22380 12888 22432
rect 12940 22420 12946 22432
rect 12977 22423 13035 22429
rect 12977 22420 12989 22423
rect 12940 22392 12989 22420
rect 12940 22380 12946 22392
rect 12977 22389 12989 22392
rect 13023 22389 13035 22423
rect 12977 22383 13035 22389
rect 13342 22380 13348 22432
rect 13400 22420 13406 22432
rect 13805 22423 13863 22429
rect 13805 22420 13817 22423
rect 13400 22392 13817 22420
rect 13400 22380 13406 22392
rect 13805 22389 13817 22392
rect 13851 22420 13863 22423
rect 14188 22420 14216 22451
rect 15826 22448 15832 22460
rect 15884 22448 15890 22500
rect 17666 22488 17672 22500
rect 17627 22460 17672 22488
rect 17666 22448 17672 22460
rect 17724 22448 17730 22500
rect 17761 22491 17819 22497
rect 17761 22457 17773 22491
rect 17807 22457 17819 22491
rect 20702 22488 20708 22500
rect 20663 22460 20708 22488
rect 17761 22451 17819 22457
rect 16654 22420 16660 22432
rect 13851 22392 14216 22420
rect 16615 22392 16660 22420
rect 13851 22389 13863 22392
rect 13805 22383 13863 22389
rect 16654 22380 16660 22392
rect 16712 22380 16718 22432
rect 17206 22380 17212 22432
rect 17264 22420 17270 22432
rect 17776 22420 17804 22451
rect 20702 22448 20708 22460
rect 20760 22448 20766 22500
rect 20797 22491 20855 22497
rect 20797 22457 20809 22491
rect 20843 22457 20855 22491
rect 20797 22451 20855 22457
rect 23373 22491 23431 22497
rect 23373 22457 23385 22491
rect 23419 22457 23431 22491
rect 23373 22451 23431 22457
rect 17264 22392 17804 22420
rect 17264 22380 17270 22392
rect 18126 22380 18132 22432
rect 18184 22420 18190 22432
rect 18589 22423 18647 22429
rect 18589 22420 18601 22423
rect 18184 22392 18601 22420
rect 18184 22380 18190 22392
rect 18589 22389 18601 22392
rect 18635 22389 18647 22423
rect 18589 22383 18647 22389
rect 20521 22423 20579 22429
rect 20521 22389 20533 22423
rect 20567 22420 20579 22423
rect 20610 22420 20616 22432
rect 20567 22392 20616 22420
rect 20567 22389 20579 22392
rect 20521 22383 20579 22389
rect 20610 22380 20616 22392
rect 20668 22420 20674 22432
rect 20812 22420 20840 22451
rect 20668 22392 20840 22420
rect 22637 22423 22695 22429
rect 20668 22380 20674 22392
rect 22637 22389 22649 22423
rect 22683 22420 22695 22423
rect 23186 22420 23192 22432
rect 22683 22392 23192 22420
rect 22683 22389 22695 22392
rect 22637 22383 22695 22389
rect 23186 22380 23192 22392
rect 23244 22420 23250 22432
rect 23388 22420 23416 22451
rect 23244 22392 23416 22420
rect 23244 22380 23250 22392
rect 632 22330 26392 22352
rect 632 22278 9843 22330
rect 9895 22278 9907 22330
rect 9959 22278 9971 22330
rect 10023 22278 10035 22330
rect 10087 22278 19176 22330
rect 19228 22278 19240 22330
rect 19292 22278 19304 22330
rect 19356 22278 19368 22330
rect 19420 22278 26392 22330
rect 632 22256 26392 22278
rect 10858 22216 10864 22228
rect 10819 22188 10864 22216
rect 10858 22176 10864 22188
rect 10916 22176 10922 22228
rect 11870 22216 11876 22228
rect 11831 22188 11876 22216
rect 11870 22176 11876 22188
rect 11928 22176 11934 22228
rect 14078 22176 14084 22228
rect 14136 22216 14142 22228
rect 14173 22219 14231 22225
rect 14173 22216 14185 22219
rect 14136 22188 14185 22216
rect 14136 22176 14142 22188
rect 14173 22185 14185 22188
rect 14219 22185 14231 22219
rect 14173 22179 14231 22185
rect 19325 22219 19383 22225
rect 19325 22185 19337 22219
rect 19371 22216 19383 22219
rect 20702 22216 20708 22228
rect 19371 22188 20708 22216
rect 19371 22185 19383 22188
rect 19325 22179 19383 22185
rect 20702 22176 20708 22188
rect 20760 22176 20766 22228
rect 23278 22176 23284 22228
rect 23336 22216 23342 22228
rect 23833 22219 23891 22225
rect 23833 22216 23845 22219
rect 23336 22188 23845 22216
rect 23336 22176 23342 22188
rect 23833 22185 23845 22188
rect 23879 22185 23891 22219
rect 23833 22179 23891 22185
rect 9570 22148 9576 22160
rect 9531 22120 9576 22148
rect 9570 22108 9576 22120
rect 9628 22108 9634 22160
rect 10125 22151 10183 22157
rect 10125 22117 10137 22151
rect 10171 22148 10183 22151
rect 10214 22148 10220 22160
rect 10171 22120 10220 22148
rect 10171 22117 10183 22120
rect 10125 22111 10183 22117
rect 10214 22108 10220 22120
rect 10272 22108 10278 22160
rect 14906 22148 14912 22160
rect 14740 22120 14912 22148
rect 1014 22089 1020 22092
rect 992 22083 1020 22089
rect 992 22049 1004 22083
rect 992 22043 1020 22049
rect 1014 22040 1020 22043
rect 1072 22040 1078 22092
rect 11318 22040 11324 22092
rect 11376 22080 11382 22092
rect 11689 22083 11747 22089
rect 11689 22080 11701 22083
rect 11376 22052 11701 22080
rect 11376 22040 11382 22052
rect 11689 22049 11701 22052
rect 11735 22049 11747 22083
rect 11689 22043 11747 22049
rect 13250 22040 13256 22092
rect 13308 22080 13314 22092
rect 13802 22080 13808 22092
rect 13308 22052 13808 22080
rect 13308 22040 13314 22052
rect 13802 22040 13808 22052
rect 13860 22040 13866 22092
rect 13897 22083 13955 22089
rect 13897 22049 13909 22083
rect 13943 22080 13955 22083
rect 14740 22080 14768 22120
rect 14906 22108 14912 22120
rect 14964 22148 14970 22160
rect 15001 22151 15059 22157
rect 15001 22148 15013 22151
rect 14964 22120 15013 22148
rect 14964 22108 14970 22120
rect 15001 22117 15013 22120
rect 15047 22117 15059 22151
rect 15001 22111 15059 22117
rect 15553 22151 15611 22157
rect 15553 22117 15565 22151
rect 15599 22148 15611 22151
rect 15642 22148 15648 22160
rect 15599 22120 15648 22148
rect 15599 22117 15611 22120
rect 15553 22111 15611 22117
rect 15642 22108 15648 22120
rect 15700 22108 15706 22160
rect 18126 22148 18132 22160
rect 18087 22120 18132 22148
rect 18126 22108 18132 22120
rect 18184 22108 18190 22160
rect 20242 22108 20248 22160
rect 20300 22148 20306 22160
rect 20613 22151 20671 22157
rect 20613 22148 20625 22151
rect 20300 22120 20625 22148
rect 20300 22108 20306 22120
rect 20613 22117 20625 22120
rect 20659 22117 20671 22151
rect 23002 22148 23008 22160
rect 22963 22120 23008 22148
rect 20613 22111 20671 22117
rect 23002 22108 23008 22120
rect 23060 22108 23066 22160
rect 23554 22148 23560 22160
rect 23515 22120 23560 22148
rect 23554 22108 23560 22120
rect 23612 22108 23618 22160
rect 13943 22052 14768 22080
rect 13943 22049 13955 22052
rect 13897 22043 13955 22049
rect 17390 22040 17396 22092
rect 17448 22080 17454 22092
rect 17758 22080 17764 22092
rect 17448 22052 17764 22080
rect 17448 22040 17454 22052
rect 17758 22040 17764 22052
rect 17816 22040 17822 22092
rect 24474 22089 24480 22092
rect 24452 22083 24480 22089
rect 24452 22049 24464 22083
rect 24452 22043 24480 22049
rect 24474 22040 24480 22043
rect 24532 22040 24538 22092
rect 9478 22012 9484 22024
rect 9439 21984 9484 22012
rect 9478 21972 9484 21984
rect 9536 21972 9542 22024
rect 14909 22015 14967 22021
rect 14909 21981 14921 22015
rect 14955 22012 14967 22015
rect 15918 22012 15924 22024
rect 14955 21984 15924 22012
rect 14955 21981 14967 21984
rect 14909 21975 14967 21981
rect 15918 21972 15924 21984
rect 15976 21972 15982 22024
rect 20518 22012 20524 22024
rect 20479 21984 20524 22012
rect 20518 21972 20524 21984
rect 20576 21972 20582 22024
rect 20794 22012 20800 22024
rect 20755 21984 20800 22012
rect 20794 21972 20800 21984
rect 20852 21972 20858 22024
rect 22542 21972 22548 22024
rect 22600 22012 22606 22024
rect 22913 22015 22971 22021
rect 22913 22012 22925 22015
rect 22600 21984 22925 22012
rect 22600 21972 22606 21984
rect 22913 21981 22925 21984
rect 22959 21981 22971 22015
rect 22913 21975 22971 21981
rect 1063 21879 1121 21885
rect 1063 21845 1075 21879
rect 1109 21876 1121 21879
rect 2210 21876 2216 21888
rect 1109 21848 2216 21876
rect 1109 21845 1121 21848
rect 1063 21839 1121 21845
rect 2210 21836 2216 21848
rect 2268 21836 2274 21888
rect 12054 21836 12060 21888
rect 12112 21876 12118 21888
rect 12698 21876 12704 21888
rect 12112 21848 12704 21876
rect 12112 21836 12118 21848
rect 12698 21836 12704 21848
rect 12756 21836 12762 21888
rect 15826 21876 15832 21888
rect 15787 21848 15832 21876
rect 15826 21836 15832 21848
rect 15884 21836 15890 21888
rect 18494 21876 18500 21888
rect 18455 21848 18500 21876
rect 18494 21836 18500 21848
rect 18552 21836 18558 21888
rect 24382 21836 24388 21888
rect 24440 21876 24446 21888
rect 24523 21879 24581 21885
rect 24523 21876 24535 21879
rect 24440 21848 24535 21876
rect 24440 21836 24446 21848
rect 24523 21845 24535 21848
rect 24569 21845 24581 21879
rect 24523 21839 24581 21845
rect 632 21786 26392 21808
rect 632 21734 5176 21786
rect 5228 21734 5240 21786
rect 5292 21734 5304 21786
rect 5356 21734 5368 21786
rect 5420 21734 14510 21786
rect 14562 21734 14574 21786
rect 14626 21734 14638 21786
rect 14690 21734 14702 21786
rect 14754 21734 23843 21786
rect 23895 21734 23907 21786
rect 23959 21734 23971 21786
rect 24023 21734 24035 21786
rect 24087 21734 26392 21786
rect 632 21712 26392 21734
rect 1014 21632 1020 21684
rect 1072 21672 1078 21684
rect 1109 21675 1167 21681
rect 1109 21672 1121 21675
rect 1072 21644 1121 21672
rect 1072 21632 1078 21644
rect 1109 21641 1121 21644
rect 1155 21641 1167 21675
rect 1109 21635 1167 21641
rect 4142 21632 4148 21684
rect 4200 21672 4206 21684
rect 4237 21675 4295 21681
rect 4237 21672 4249 21675
rect 4200 21644 4249 21672
rect 4200 21632 4206 21644
rect 4237 21641 4249 21644
rect 4283 21641 4295 21675
rect 4237 21635 4295 21641
rect 9570 21632 9576 21684
rect 9628 21672 9634 21684
rect 9941 21675 9999 21681
rect 9941 21672 9953 21675
rect 9628 21644 9953 21672
rect 9628 21632 9634 21644
rect 9941 21641 9953 21644
rect 9987 21672 9999 21675
rect 10214 21672 10220 21684
rect 9987 21644 10220 21672
rect 9987 21641 9999 21644
rect 9941 21635 9999 21641
rect 10214 21632 10220 21644
rect 10272 21632 10278 21684
rect 11318 21632 11324 21684
rect 11376 21672 11382 21684
rect 11597 21675 11655 21681
rect 11597 21672 11609 21675
rect 11376 21644 11609 21672
rect 11376 21632 11382 21644
rect 11597 21641 11609 21644
rect 11643 21641 11655 21675
rect 12514 21672 12520 21684
rect 12475 21644 12520 21672
rect 11597 21635 11655 21641
rect 12514 21632 12520 21644
rect 12572 21632 12578 21684
rect 13069 21675 13127 21681
rect 13069 21641 13081 21675
rect 13115 21672 13127 21675
rect 13802 21672 13808 21684
rect 13115 21644 13808 21672
rect 13115 21641 13127 21644
rect 13069 21635 13127 21641
rect 13802 21632 13808 21644
rect 13860 21672 13866 21684
rect 14449 21675 14507 21681
rect 14449 21672 14461 21675
rect 13860 21644 14461 21672
rect 13860 21632 13866 21644
rect 14449 21641 14461 21644
rect 14495 21641 14507 21675
rect 14906 21672 14912 21684
rect 14867 21644 14912 21672
rect 14449 21635 14507 21641
rect 14906 21632 14912 21644
rect 14964 21632 14970 21684
rect 17758 21672 17764 21684
rect 17719 21644 17764 21672
rect 17758 21632 17764 21644
rect 17816 21632 17822 21684
rect 20610 21672 20616 21684
rect 20571 21644 20616 21672
rect 20610 21632 20616 21644
rect 20668 21632 20674 21684
rect 21714 21632 21720 21684
rect 21772 21672 21778 21684
rect 22085 21675 22143 21681
rect 22085 21672 22097 21675
rect 21772 21644 22097 21672
rect 21772 21632 21778 21644
rect 22085 21641 22097 21644
rect 22131 21641 22143 21675
rect 22542 21672 22548 21684
rect 22503 21644 22548 21672
rect 22085 21635 22143 21641
rect 22542 21632 22548 21644
rect 22600 21632 22606 21684
rect 24474 21672 24480 21684
rect 24435 21644 24480 21672
rect 24474 21632 24480 21644
rect 24532 21632 24538 21684
rect 25302 21672 25308 21684
rect 25263 21644 25308 21672
rect 25302 21632 25308 21644
rect 25360 21632 25366 21684
rect 15829 21607 15887 21613
rect 15829 21573 15841 21607
rect 15875 21604 15887 21607
rect 15918 21604 15924 21616
rect 15875 21576 15924 21604
rect 15875 21573 15887 21576
rect 15829 21567 15887 21573
rect 15918 21564 15924 21576
rect 15976 21564 15982 21616
rect 20518 21564 20524 21616
rect 20576 21604 20582 21616
rect 21349 21607 21407 21613
rect 21349 21604 21361 21607
rect 20576 21576 21361 21604
rect 20576 21564 20582 21576
rect 21349 21573 21361 21576
rect 21395 21573 21407 21607
rect 21349 21567 21407 21573
rect 7454 21536 7460 21548
rect 7415 21508 7460 21536
rect 7454 21496 7460 21508
rect 7512 21496 7518 21548
rect 8101 21539 8159 21545
rect 8101 21505 8113 21539
rect 8147 21536 8159 21539
rect 9297 21539 9355 21545
rect 9297 21536 9309 21539
rect 8147 21508 9309 21536
rect 8147 21505 8159 21508
rect 8101 21499 8159 21505
rect 9297 21505 9309 21508
rect 9343 21536 9355 21539
rect 9478 21536 9484 21548
rect 9343 21508 9484 21536
rect 9343 21505 9355 21508
rect 9297 21499 9355 21505
rect 9478 21496 9484 21508
rect 9536 21536 9542 21548
rect 10309 21539 10367 21545
rect 10309 21536 10321 21539
rect 9536 21508 10321 21536
rect 9536 21496 9542 21508
rect 10309 21505 10321 21508
rect 10355 21505 10367 21539
rect 10309 21499 10367 21505
rect 15090 21496 15096 21548
rect 15148 21536 15154 21548
rect 15277 21539 15335 21545
rect 15277 21536 15289 21539
rect 15148 21508 15289 21536
rect 15148 21496 15154 21508
rect 15277 21505 15289 21508
rect 15323 21505 15335 21539
rect 18954 21536 18960 21548
rect 18915 21508 18960 21536
rect 15277 21499 15335 21505
rect 18954 21496 18960 21508
rect 19012 21496 19018 21548
rect 22913 21539 22971 21545
rect 22913 21505 22925 21539
rect 22959 21536 22971 21539
rect 23002 21536 23008 21548
rect 22959 21508 23008 21536
rect 22959 21505 22971 21508
rect 22913 21499 22971 21505
rect 23002 21496 23008 21508
rect 23060 21536 23066 21548
rect 23189 21539 23247 21545
rect 23189 21536 23201 21539
rect 23060 21508 23201 21536
rect 23060 21496 23066 21508
rect 23189 21505 23201 21508
rect 23235 21505 23247 21539
rect 23189 21499 23247 21505
rect 3844 21471 3902 21477
rect 3844 21437 3856 21471
rect 3890 21468 3902 21471
rect 4142 21468 4148 21480
rect 3890 21440 4148 21468
rect 3890 21437 3902 21440
rect 3844 21431 3902 21437
rect 4142 21428 4148 21440
rect 4200 21428 4206 21480
rect 12124 21471 12182 21477
rect 12124 21437 12136 21471
rect 12170 21468 12182 21471
rect 12514 21468 12520 21480
rect 12170 21440 12520 21468
rect 12170 21437 12182 21440
rect 12124 21431 12182 21437
rect 12514 21428 12520 21440
rect 12572 21428 12578 21480
rect 13529 21471 13587 21477
rect 13529 21437 13541 21471
rect 13575 21468 13587 21471
rect 13618 21468 13624 21480
rect 13575 21440 13624 21468
rect 13575 21437 13587 21440
rect 13529 21431 13587 21437
rect 13618 21428 13624 21440
rect 13676 21428 13682 21480
rect 19877 21471 19935 21477
rect 19877 21437 19889 21471
rect 19923 21468 19935 21471
rect 20150 21468 20156 21480
rect 19923 21440 20156 21468
rect 19923 21437 19935 21440
rect 19877 21431 19935 21437
rect 20150 21428 20156 21440
rect 20208 21468 20214 21480
rect 20702 21468 20708 21480
rect 20208 21440 20708 21468
rect 20208 21428 20214 21440
rect 20702 21428 20708 21440
rect 20760 21428 20766 21480
rect 21901 21471 21959 21477
rect 21901 21468 21913 21471
rect 21732 21440 21913 21468
rect 7273 21403 7331 21409
rect 7273 21369 7285 21403
rect 7319 21400 7331 21403
rect 7549 21403 7607 21409
rect 7549 21400 7561 21403
rect 7319 21372 7561 21400
rect 7319 21369 7331 21372
rect 7273 21363 7331 21369
rect 7549 21369 7561 21372
rect 7595 21400 7607 21403
rect 7638 21400 7644 21412
rect 7595 21372 7644 21400
rect 7595 21369 7607 21372
rect 7549 21363 7607 21369
rect 7638 21360 7644 21372
rect 7696 21360 7702 21412
rect 9018 21400 9024 21412
rect 8979 21372 9024 21400
rect 9018 21360 9024 21372
rect 9076 21360 9082 21412
rect 9113 21403 9171 21409
rect 9113 21369 9125 21403
rect 9159 21369 9171 21403
rect 9113 21363 9171 21369
rect 3915 21335 3973 21341
rect 3915 21301 3927 21335
rect 3961 21332 3973 21335
rect 4970 21332 4976 21344
rect 3961 21304 4976 21332
rect 3961 21301 3973 21304
rect 3915 21295 3973 21301
rect 4970 21292 4976 21304
rect 5028 21292 5034 21344
rect 8742 21332 8748 21344
rect 8703 21304 8748 21332
rect 8742 21292 8748 21304
rect 8800 21332 8806 21344
rect 9128 21332 9156 21363
rect 11686 21360 11692 21412
rect 11744 21400 11750 21412
rect 13345 21403 13403 21409
rect 13345 21400 13357 21403
rect 11744 21372 13357 21400
rect 11744 21360 11750 21372
rect 13345 21369 13357 21372
rect 13391 21400 13403 21403
rect 13850 21403 13908 21409
rect 13850 21400 13862 21403
rect 13391 21372 13862 21400
rect 13391 21369 13403 21372
rect 13345 21363 13403 21369
rect 13850 21369 13862 21372
rect 13896 21369 13908 21403
rect 18494 21400 18500 21412
rect 18455 21372 18500 21400
rect 13850 21363 13908 21369
rect 18494 21360 18500 21372
rect 18552 21360 18558 21412
rect 18586 21360 18592 21412
rect 18644 21400 18650 21412
rect 18644 21372 18689 21400
rect 18644 21360 18650 21372
rect 12238 21341 12244 21344
rect 8800 21304 9156 21332
rect 12195 21335 12244 21341
rect 8800 21292 8806 21304
rect 12195 21301 12207 21335
rect 12241 21301 12244 21335
rect 12195 21295 12244 21301
rect 12238 21292 12244 21295
rect 12296 21292 12302 21344
rect 18313 21335 18371 21341
rect 18313 21301 18325 21335
rect 18359 21332 18371 21335
rect 18604 21332 18632 21360
rect 20242 21332 20248 21344
rect 18359 21304 18632 21332
rect 20203 21304 20248 21332
rect 18359 21301 18371 21304
rect 18313 21295 18371 21301
rect 20242 21292 20248 21304
rect 20300 21292 20306 21344
rect 21622 21292 21628 21344
rect 21680 21332 21686 21344
rect 21732 21341 21760 21440
rect 21901 21437 21913 21440
rect 21947 21437 21959 21471
rect 23278 21468 23284 21480
rect 23239 21440 23284 21468
rect 21901 21431 21959 21437
rect 23278 21428 23284 21440
rect 23336 21428 23342 21480
rect 24820 21471 24878 21477
rect 24820 21437 24832 21471
rect 24866 21468 24878 21471
rect 25302 21468 25308 21480
rect 24866 21440 25308 21468
rect 24866 21437 24878 21440
rect 24820 21431 24878 21437
rect 25302 21428 25308 21440
rect 25360 21428 25366 21480
rect 21717 21335 21775 21341
rect 21717 21332 21729 21335
rect 21680 21304 21729 21332
rect 21680 21292 21686 21304
rect 21717 21301 21729 21304
rect 21763 21301 21775 21335
rect 21717 21295 21775 21301
rect 24474 21292 24480 21344
rect 24532 21332 24538 21344
rect 24891 21335 24949 21341
rect 24891 21332 24903 21335
rect 24532 21304 24903 21332
rect 24532 21292 24538 21304
rect 24891 21301 24903 21304
rect 24937 21301 24949 21335
rect 24891 21295 24949 21301
rect 632 21242 26392 21264
rect 632 21190 9843 21242
rect 9895 21190 9907 21242
rect 9959 21190 9971 21242
rect 10023 21190 10035 21242
rect 10087 21190 19176 21242
rect 19228 21190 19240 21242
rect 19292 21190 19304 21242
rect 19356 21190 19368 21242
rect 19420 21190 26392 21242
rect 632 21168 26392 21190
rect 7454 21128 7460 21140
rect 7415 21100 7460 21128
rect 7454 21088 7460 21100
rect 7512 21088 7518 21140
rect 10214 21128 10220 21140
rect 10175 21100 10220 21128
rect 10214 21088 10220 21100
rect 10272 21088 10278 21140
rect 11318 21088 11324 21140
rect 11376 21128 11382 21140
rect 12241 21131 12299 21137
rect 12241 21128 12253 21131
rect 11376 21100 12253 21128
rect 11376 21088 11382 21100
rect 12241 21097 12253 21100
rect 12287 21097 12299 21131
rect 12241 21091 12299 21097
rect 17301 21131 17359 21137
rect 17301 21097 17313 21131
rect 17347 21128 17359 21131
rect 17758 21128 17764 21140
rect 17347 21100 17764 21128
rect 17347 21097 17359 21100
rect 17301 21091 17359 21097
rect 17758 21088 17764 21100
rect 17816 21088 17822 21140
rect 22542 21088 22548 21140
rect 22600 21128 22606 21140
rect 22913 21131 22971 21137
rect 22913 21128 22925 21131
rect 22600 21100 22925 21128
rect 22600 21088 22606 21100
rect 22913 21097 22925 21100
rect 22959 21097 22971 21131
rect 22913 21091 22971 21097
rect 24198 21088 24204 21140
rect 24256 21128 24262 21140
rect 24293 21131 24351 21137
rect 24293 21128 24305 21131
rect 24256 21100 24305 21128
rect 24256 21088 24262 21100
rect 24293 21097 24305 21100
rect 24339 21097 24351 21131
rect 24293 21091 24351 21097
rect 8285 21063 8343 21069
rect 8285 21029 8297 21063
rect 8331 21060 8343 21063
rect 8742 21060 8748 21072
rect 8331 21032 8748 21060
rect 8331 21029 8343 21032
rect 8285 21023 8343 21029
rect 8742 21020 8748 21032
rect 8800 21020 8806 21072
rect 9662 21069 9668 21072
rect 9659 21060 9668 21069
rect 9623 21032 9668 21060
rect 9659 21023 9668 21032
rect 9662 21020 9668 21023
rect 9720 21020 9726 21072
rect 11686 21069 11692 21072
rect 11683 21060 11692 21069
rect 11647 21032 11692 21060
rect 11683 21023 11692 21032
rect 11686 21020 11692 21023
rect 11744 21020 11750 21072
rect 16746 21069 16752 21072
rect 16743 21060 16752 21069
rect 16707 21032 16752 21060
rect 16743 21023 16752 21032
rect 16746 21020 16752 21023
rect 16804 21020 16810 21072
rect 18681 21063 18739 21069
rect 18681 21029 18693 21063
rect 18727 21060 18739 21063
rect 18862 21060 18868 21072
rect 18727 21032 18868 21060
rect 18727 21029 18739 21032
rect 18681 21023 18739 21029
rect 18862 21020 18868 21032
rect 18920 21060 18926 21072
rect 18957 21063 19015 21069
rect 18957 21060 18969 21063
rect 18920 21032 18969 21060
rect 18920 21020 18926 21032
rect 18957 21029 18969 21032
rect 19003 21029 19015 21063
rect 20426 21060 20432 21072
rect 20387 21032 20432 21060
rect 18957 21023 19015 21029
rect 20426 21020 20432 21032
rect 20484 21020 20490 21072
rect 7638 20952 7644 21004
rect 7696 20992 7702 21004
rect 8193 20995 8251 21001
rect 8193 20992 8205 20995
rect 7696 20964 8205 20992
rect 7696 20952 7702 20964
rect 8193 20961 8205 20964
rect 8239 20992 8251 20995
rect 9110 20992 9116 21004
rect 8239 20964 9116 20992
rect 8239 20961 8251 20964
rect 8193 20955 8251 20961
rect 9110 20952 9116 20964
rect 9168 20952 9174 21004
rect 15093 20995 15151 21001
rect 15093 20961 15105 20995
rect 15139 20961 15151 20995
rect 15366 20992 15372 21004
rect 15327 20964 15372 20992
rect 15093 20955 15151 20961
rect 9294 20924 9300 20936
rect 9255 20896 9300 20924
rect 9294 20884 9300 20896
rect 9352 20884 9358 20936
rect 11226 20884 11232 20936
rect 11284 20924 11290 20936
rect 11321 20927 11379 20933
rect 11321 20924 11333 20927
rect 11284 20896 11333 20924
rect 11284 20884 11290 20896
rect 11321 20893 11333 20896
rect 11367 20893 11379 20927
rect 15108 20924 15136 20955
rect 15366 20952 15372 20964
rect 15424 20952 15430 21004
rect 20518 20992 20524 21004
rect 20479 20964 20524 20992
rect 20518 20952 20524 20964
rect 20576 20952 20582 21004
rect 24109 20995 24167 21001
rect 24109 20961 24121 20995
rect 24155 20992 24167 20995
rect 24382 20992 24388 21004
rect 24155 20964 24388 20992
rect 24155 20961 24167 20964
rect 24109 20955 24167 20961
rect 24382 20952 24388 20964
rect 24440 20952 24446 21004
rect 15274 20924 15280 20936
rect 15108 20896 15280 20924
rect 11321 20887 11379 20893
rect 15274 20884 15280 20896
rect 15332 20884 15338 20936
rect 15553 20927 15611 20933
rect 15553 20893 15565 20927
rect 15599 20924 15611 20927
rect 15734 20924 15740 20936
rect 15599 20896 15740 20924
rect 15599 20893 15611 20896
rect 15553 20887 15611 20893
rect 15734 20884 15740 20896
rect 15792 20924 15798 20936
rect 15829 20927 15887 20933
rect 15829 20924 15841 20927
rect 15792 20896 15841 20924
rect 15792 20884 15798 20896
rect 15829 20893 15841 20896
rect 15875 20893 15887 20927
rect 16378 20924 16384 20936
rect 16339 20896 16384 20924
rect 15829 20887 15887 20893
rect 16378 20884 16384 20896
rect 16436 20884 16442 20936
rect 18865 20927 18923 20933
rect 18865 20893 18877 20927
rect 18911 20924 18923 20927
rect 18954 20924 18960 20936
rect 18911 20896 18960 20924
rect 18911 20893 18923 20896
rect 18865 20887 18923 20893
rect 18954 20884 18960 20896
rect 19012 20884 19018 20936
rect 19506 20924 19512 20936
rect 19467 20896 19512 20924
rect 19506 20884 19512 20896
rect 19564 20884 19570 20936
rect 9018 20788 9024 20800
rect 8979 20760 9024 20788
rect 9018 20748 9024 20760
rect 9076 20748 9082 20800
rect 13618 20788 13624 20800
rect 13579 20760 13624 20788
rect 13618 20748 13624 20760
rect 13676 20748 13682 20800
rect 13894 20748 13900 20800
rect 13952 20788 13958 20800
rect 13989 20791 14047 20797
rect 13989 20788 14001 20791
rect 13952 20760 14001 20788
rect 13952 20748 13958 20760
rect 13989 20757 14001 20760
rect 14035 20757 14047 20791
rect 17666 20788 17672 20800
rect 17627 20760 17672 20788
rect 13989 20751 14047 20757
rect 17666 20748 17672 20760
rect 17724 20748 17730 20800
rect 23002 20748 23008 20800
rect 23060 20788 23066 20800
rect 23278 20788 23284 20800
rect 23060 20760 23284 20788
rect 23060 20748 23066 20760
rect 23278 20748 23284 20760
rect 23336 20788 23342 20800
rect 23373 20791 23431 20797
rect 23373 20788 23385 20791
rect 23336 20760 23385 20788
rect 23336 20748 23342 20760
rect 23373 20757 23385 20760
rect 23419 20757 23431 20791
rect 23373 20751 23431 20757
rect 632 20698 26392 20720
rect 632 20646 5176 20698
rect 5228 20646 5240 20698
rect 5292 20646 5304 20698
rect 5356 20646 5368 20698
rect 5420 20646 14510 20698
rect 14562 20646 14574 20698
rect 14626 20646 14638 20698
rect 14690 20646 14702 20698
rect 14754 20646 23843 20698
rect 23895 20646 23907 20698
rect 23959 20646 23971 20698
rect 24023 20646 24035 20698
rect 24087 20646 26392 20698
rect 632 20624 26392 20646
rect 7638 20584 7644 20596
rect 7599 20556 7644 20584
rect 7638 20544 7644 20556
rect 7696 20544 7702 20596
rect 9202 20544 9208 20596
rect 9260 20584 9266 20596
rect 9941 20587 9999 20593
rect 9941 20584 9953 20587
rect 9260 20556 9953 20584
rect 9260 20544 9266 20556
rect 9941 20553 9953 20556
rect 9987 20553 9999 20587
rect 12882 20584 12888 20596
rect 12843 20556 12888 20584
rect 9941 20547 9999 20553
rect 12882 20544 12888 20556
rect 12940 20544 12946 20596
rect 14909 20587 14967 20593
rect 14909 20553 14921 20587
rect 14955 20584 14967 20587
rect 15826 20584 15832 20596
rect 14955 20556 15832 20584
rect 14955 20553 14967 20556
rect 14909 20547 14967 20553
rect 15826 20544 15832 20556
rect 15884 20544 15890 20596
rect 16654 20584 16660 20596
rect 16615 20556 16660 20584
rect 16654 20544 16660 20556
rect 16712 20544 16718 20596
rect 20518 20584 20524 20596
rect 20479 20556 20524 20584
rect 20518 20544 20524 20556
rect 20576 20544 20582 20596
rect 21714 20544 21720 20596
rect 21772 20584 21778 20596
rect 22177 20587 22235 20593
rect 22177 20584 22189 20587
rect 21772 20556 22189 20584
rect 21772 20544 21778 20556
rect 22177 20553 22189 20556
rect 22223 20553 22235 20587
rect 22177 20547 22235 20553
rect 24382 20544 24388 20596
rect 24440 20584 24446 20596
rect 24937 20587 24995 20593
rect 24937 20584 24949 20587
rect 24440 20556 24949 20584
rect 24440 20544 24446 20556
rect 24937 20553 24949 20556
rect 24983 20584 24995 20587
rect 25259 20587 25317 20593
rect 25259 20584 25271 20587
rect 24983 20556 25271 20584
rect 24983 20553 24995 20556
rect 24937 20547 24995 20553
rect 25259 20553 25271 20556
rect 25305 20553 25317 20587
rect 25259 20547 25317 20553
rect 24290 20476 24296 20528
rect 24348 20516 24354 20528
rect 24569 20519 24627 20525
rect 24569 20516 24581 20519
rect 24348 20488 24581 20516
rect 24348 20476 24354 20488
rect 24569 20485 24581 20488
rect 24615 20485 24627 20519
rect 24569 20479 24627 20485
rect 9294 20408 9300 20460
rect 9352 20448 9358 20460
rect 10217 20451 10275 20457
rect 10217 20448 10229 20451
rect 9352 20420 10229 20448
rect 9352 20408 9358 20420
rect 10217 20417 10229 20420
rect 10263 20417 10275 20451
rect 15734 20448 15740 20460
rect 15695 20420 15740 20448
rect 10217 20411 10275 20417
rect 15734 20408 15740 20420
rect 15792 20408 15798 20460
rect 18313 20451 18371 20457
rect 18313 20417 18325 20451
rect 18359 20448 18371 20451
rect 18586 20448 18592 20460
rect 18359 20420 18592 20448
rect 18359 20417 18371 20420
rect 18313 20411 18371 20417
rect 18586 20408 18592 20420
rect 18644 20448 18650 20460
rect 18954 20448 18960 20460
rect 18644 20420 18960 20448
rect 18644 20408 18650 20420
rect 18954 20408 18960 20420
rect 19012 20408 19018 20460
rect 19506 20448 19512 20460
rect 19467 20420 19512 20448
rect 19506 20408 19512 20420
rect 19564 20408 19570 20460
rect 8193 20383 8251 20389
rect 8193 20349 8205 20383
rect 8239 20380 8251 20383
rect 9021 20383 9079 20389
rect 9021 20380 9033 20383
rect 8239 20352 9033 20380
rect 8239 20349 8251 20352
rect 8193 20343 8251 20349
rect 9021 20349 9033 20352
rect 9067 20380 9079 20383
rect 9110 20380 9116 20392
rect 9067 20352 9116 20380
rect 9067 20349 9079 20352
rect 9021 20343 9079 20349
rect 9110 20340 9116 20352
rect 9168 20340 9174 20392
rect 11965 20383 12023 20389
rect 11965 20349 11977 20383
rect 12011 20380 12023 20383
rect 12054 20380 12060 20392
rect 12011 20352 12060 20380
rect 12011 20349 12023 20352
rect 11965 20343 12023 20349
rect 12054 20340 12060 20352
rect 12112 20340 12118 20392
rect 12210 20352 12376 20380
rect 8561 20315 8619 20321
rect 8561 20281 8573 20315
rect 8607 20312 8619 20315
rect 8929 20315 8987 20321
rect 8929 20312 8941 20315
rect 8607 20284 8941 20312
rect 8607 20281 8619 20284
rect 8561 20275 8619 20281
rect 8929 20281 8941 20284
rect 8975 20312 8987 20315
rect 9383 20315 9441 20321
rect 9383 20312 9395 20315
rect 8975 20284 9395 20312
rect 8975 20281 8987 20284
rect 8929 20275 8987 20281
rect 9383 20281 9395 20284
rect 9429 20312 9441 20315
rect 9662 20312 9668 20324
rect 9429 20284 9668 20312
rect 9429 20281 9441 20284
rect 9383 20275 9441 20281
rect 9662 20272 9668 20284
rect 9720 20272 9726 20324
rect 11045 20315 11103 20321
rect 11045 20281 11057 20315
rect 11091 20312 11103 20315
rect 11226 20312 11232 20324
rect 11091 20284 11232 20312
rect 11091 20281 11103 20284
rect 11045 20275 11103 20281
rect 11226 20272 11232 20284
rect 11284 20312 11290 20324
rect 11870 20312 11876 20324
rect 11284 20284 11876 20312
rect 11284 20272 11290 20284
rect 11870 20272 11876 20284
rect 11928 20272 11934 20324
rect 9680 20244 9708 20272
rect 11321 20247 11379 20253
rect 11321 20244 11333 20247
rect 9680 20216 11333 20244
rect 11321 20213 11333 20216
rect 11367 20244 11379 20247
rect 11686 20244 11692 20256
rect 11367 20216 11692 20244
rect 11367 20213 11379 20216
rect 11321 20207 11379 20213
rect 11686 20204 11692 20216
rect 11744 20244 11750 20256
rect 12210 20244 12238 20352
rect 12348 20321 12376 20352
rect 13894 20340 13900 20392
rect 13952 20380 13958 20392
rect 13989 20383 14047 20389
rect 13989 20380 14001 20383
rect 13952 20352 14001 20380
rect 13952 20340 13958 20352
rect 13989 20349 14001 20352
rect 14035 20349 14047 20383
rect 16746 20380 16752 20392
rect 13989 20343 14047 20349
rect 16212 20352 16752 20380
rect 16212 20324 16240 20352
rect 16746 20340 16752 20352
rect 16804 20380 16810 20392
rect 16933 20383 16991 20389
rect 16933 20380 16945 20383
rect 16804 20352 16945 20380
rect 16804 20340 16810 20352
rect 16933 20349 16945 20352
rect 16979 20349 16991 20383
rect 16933 20343 16991 20349
rect 21162 20340 21168 20392
rect 21220 20380 21226 20392
rect 21257 20383 21315 20389
rect 21257 20380 21269 20383
rect 21220 20352 21269 20380
rect 21220 20340 21226 20352
rect 21257 20349 21269 20352
rect 21303 20349 21315 20383
rect 21257 20343 21315 20349
rect 24176 20383 24234 20389
rect 24176 20349 24188 20383
rect 24222 20380 24234 20383
rect 24308 20380 24336 20476
rect 24222 20352 24336 20380
rect 24222 20349 24234 20352
rect 24176 20343 24234 20349
rect 24474 20340 24480 20392
rect 24532 20380 24538 20392
rect 25188 20383 25246 20389
rect 25188 20380 25200 20383
rect 24532 20352 25200 20380
rect 24532 20340 24538 20352
rect 25188 20349 25200 20352
rect 25234 20380 25246 20383
rect 25581 20383 25639 20389
rect 25581 20380 25593 20383
rect 25234 20352 25593 20380
rect 25234 20349 25246 20352
rect 25188 20343 25246 20349
rect 25581 20349 25593 20352
rect 25627 20349 25639 20383
rect 25581 20343 25639 20349
rect 12327 20315 12385 20321
rect 12327 20281 12339 20315
rect 12373 20312 12385 20315
rect 13805 20315 13863 20321
rect 13805 20312 13817 20315
rect 12373 20284 13817 20312
rect 12373 20281 12385 20284
rect 12327 20275 12385 20281
rect 13805 20281 13817 20284
rect 13851 20312 13863 20315
rect 14310 20315 14368 20321
rect 14310 20312 14322 20315
rect 13851 20284 14322 20312
rect 13851 20281 13863 20284
rect 13805 20275 13863 20281
rect 14310 20281 14322 20284
rect 14356 20312 14368 20315
rect 15553 20315 15611 20321
rect 15553 20312 15565 20315
rect 14356 20284 15565 20312
rect 14356 20281 14368 20284
rect 14310 20275 14368 20281
rect 15553 20281 15565 20284
rect 15599 20312 15611 20315
rect 16058 20315 16116 20321
rect 16058 20312 16070 20315
rect 15599 20284 16070 20312
rect 15599 20281 15611 20284
rect 15553 20275 15611 20281
rect 16058 20281 16070 20284
rect 16104 20312 16116 20315
rect 16194 20312 16200 20324
rect 16104 20284 16200 20312
rect 16104 20281 16116 20284
rect 16058 20275 16116 20281
rect 16194 20272 16200 20284
rect 16252 20272 16258 20324
rect 16378 20272 16384 20324
rect 16436 20312 16442 20324
rect 17301 20315 17359 20321
rect 17301 20312 17313 20315
rect 16436 20284 17313 20312
rect 16436 20272 16442 20284
rect 17301 20281 17313 20284
rect 17347 20281 17359 20315
rect 17301 20275 17359 20281
rect 17669 20315 17727 20321
rect 17669 20281 17681 20315
rect 17715 20281 17727 20315
rect 17669 20275 17727 20281
rect 15274 20244 15280 20256
rect 11744 20216 12238 20244
rect 15235 20216 15280 20244
rect 11744 20204 11750 20216
rect 15274 20204 15280 20216
rect 15332 20204 15338 20256
rect 17574 20204 17580 20256
rect 17632 20244 17638 20256
rect 17684 20244 17712 20275
rect 17758 20272 17764 20324
rect 17816 20312 17822 20324
rect 19233 20315 19291 20321
rect 19233 20312 19245 20315
rect 17816 20284 17861 20312
rect 18604 20284 19245 20312
rect 17816 20272 17822 20284
rect 17632 20216 17712 20244
rect 17632 20204 17638 20216
rect 18494 20204 18500 20256
rect 18552 20244 18558 20256
rect 18604 20253 18632 20284
rect 19233 20281 19245 20284
rect 19279 20281 19291 20315
rect 19233 20275 19291 20281
rect 19325 20315 19383 20321
rect 19325 20281 19337 20315
rect 19371 20281 19383 20315
rect 21578 20315 21636 20321
rect 21578 20312 21590 20315
rect 19325 20275 19383 20281
rect 21088 20284 21590 20312
rect 18589 20247 18647 20253
rect 18589 20244 18601 20247
rect 18552 20216 18601 20244
rect 18552 20204 18558 20216
rect 18589 20213 18601 20216
rect 18635 20213 18647 20247
rect 18954 20244 18960 20256
rect 18915 20216 18960 20244
rect 18589 20207 18647 20213
rect 18954 20204 18960 20216
rect 19012 20244 19018 20256
rect 19340 20244 19368 20275
rect 21088 20256 21116 20284
rect 21578 20281 21590 20284
rect 21624 20281 21636 20315
rect 21578 20275 21636 20281
rect 21070 20244 21076 20256
rect 19012 20216 19368 20244
rect 21031 20216 21076 20244
rect 19012 20204 19018 20216
rect 21070 20204 21076 20216
rect 21128 20204 21134 20256
rect 23002 20204 23008 20256
rect 23060 20244 23066 20256
rect 24247 20247 24305 20253
rect 24247 20244 24259 20247
rect 23060 20216 24259 20244
rect 23060 20204 23066 20216
rect 24247 20213 24259 20216
rect 24293 20213 24305 20247
rect 24247 20207 24305 20213
rect 632 20154 26392 20176
rect 632 20102 9843 20154
rect 9895 20102 9907 20154
rect 9959 20102 9971 20154
rect 10023 20102 10035 20154
rect 10087 20102 19176 20154
rect 19228 20102 19240 20154
rect 19292 20102 19304 20154
rect 19356 20102 19368 20154
rect 19420 20102 26392 20154
rect 632 20080 26392 20102
rect 9294 20000 9300 20052
rect 9352 20040 9358 20052
rect 9573 20043 9631 20049
rect 9573 20040 9585 20043
rect 9352 20012 9585 20040
rect 9352 20000 9358 20012
rect 9573 20009 9585 20012
rect 9619 20009 9631 20043
rect 9573 20003 9631 20009
rect 17393 20043 17451 20049
rect 17393 20009 17405 20043
rect 17439 20040 17451 20043
rect 17666 20040 17672 20052
rect 17439 20012 17672 20040
rect 17439 20009 17451 20012
rect 17393 20003 17451 20009
rect 17666 20000 17672 20012
rect 17724 20000 17730 20052
rect 18586 20040 18592 20052
rect 18547 20012 18592 20040
rect 18586 20000 18592 20012
rect 18644 20000 18650 20052
rect 18954 20040 18960 20052
rect 18915 20012 18960 20040
rect 18954 20000 18960 20012
rect 19012 20000 19018 20052
rect 20567 20043 20625 20049
rect 20567 20009 20579 20043
rect 20613 20040 20625 20043
rect 21530 20040 21536 20052
rect 20613 20012 21536 20040
rect 20613 20009 20625 20012
rect 20567 20003 20625 20009
rect 21530 20000 21536 20012
rect 21588 20000 21594 20052
rect 22453 20043 22511 20049
rect 22453 20009 22465 20043
rect 22499 20040 22511 20043
rect 22910 20040 22916 20052
rect 22499 20012 22916 20040
rect 22499 20009 22511 20012
rect 22453 20003 22511 20009
rect 22910 20000 22916 20012
rect 22968 20000 22974 20052
rect 13894 19972 13900 19984
rect 13855 19944 13900 19972
rect 13894 19932 13900 19944
rect 13952 19932 13958 19984
rect 15645 19975 15703 19981
rect 15645 19941 15657 19975
rect 15691 19972 15703 19975
rect 16378 19972 16384 19984
rect 15691 19944 16384 19972
rect 15691 19941 15703 19944
rect 15645 19935 15703 19941
rect 16378 19932 16384 19944
rect 16436 19932 16442 19984
rect 16746 19932 16752 19984
rect 16804 19981 16810 19984
rect 16804 19975 16852 19981
rect 16804 19941 16806 19975
rect 16840 19941 16852 19975
rect 16804 19935 16852 19941
rect 16804 19932 16810 19935
rect 21070 19932 21076 19984
rect 21128 19972 21134 19984
rect 21854 19975 21912 19981
rect 21854 19972 21866 19975
rect 21128 19944 21866 19972
rect 21128 19932 21134 19944
rect 21854 19941 21866 19944
rect 21900 19941 21912 19975
rect 21854 19935 21912 19941
rect 9481 19907 9539 19913
rect 9481 19873 9493 19907
rect 9527 19873 9539 19907
rect 9481 19867 9539 19873
rect 9496 19836 9524 19867
rect 9570 19864 9576 19916
rect 9628 19904 9634 19916
rect 9941 19907 9999 19913
rect 9941 19904 9953 19907
rect 9628 19876 9953 19904
rect 9628 19864 9634 19876
rect 9941 19873 9953 19876
rect 9987 19873 9999 19907
rect 11502 19904 11508 19916
rect 11463 19876 11508 19904
rect 9941 19867 9999 19873
rect 11502 19864 11508 19876
rect 11560 19864 11566 19916
rect 11965 19907 12023 19913
rect 11965 19873 11977 19907
rect 12011 19904 12023 19907
rect 12146 19904 12152 19916
rect 12011 19876 12152 19904
rect 12011 19873 12023 19876
rect 11965 19867 12023 19873
rect 12146 19864 12152 19876
rect 12204 19864 12210 19916
rect 13342 19904 13348 19916
rect 13303 19876 13348 19904
rect 13342 19864 13348 19876
rect 13400 19864 13406 19916
rect 13713 19907 13771 19913
rect 13713 19873 13725 19907
rect 13759 19904 13771 19907
rect 13986 19904 13992 19916
rect 13759 19876 13992 19904
rect 13759 19873 13771 19876
rect 13713 19867 13771 19873
rect 13986 19864 13992 19876
rect 14044 19864 14050 19916
rect 14906 19904 14912 19916
rect 14867 19876 14912 19904
rect 14906 19864 14912 19876
rect 14964 19864 14970 19916
rect 15366 19904 15372 19916
rect 15279 19876 15372 19904
rect 15366 19864 15372 19876
rect 15424 19864 15430 19916
rect 17666 19904 17672 19916
rect 17627 19876 17672 19904
rect 17666 19864 17672 19876
rect 17724 19864 17730 19916
rect 18862 19904 18868 19916
rect 18823 19876 18868 19904
rect 18862 19864 18868 19876
rect 18920 19864 18926 19916
rect 19506 19864 19512 19916
rect 19564 19904 19570 19916
rect 20464 19907 20522 19913
rect 20464 19904 20476 19907
rect 19564 19876 20476 19904
rect 19564 19864 19570 19876
rect 20464 19873 20476 19876
rect 20510 19904 20522 19907
rect 20978 19904 20984 19916
rect 20510 19876 20984 19904
rect 20510 19873 20522 19876
rect 20464 19867 20522 19873
rect 20978 19864 20984 19876
rect 21036 19864 21042 19916
rect 23646 19904 23652 19916
rect 23607 19876 23652 19904
rect 23646 19864 23652 19876
rect 23704 19864 23710 19916
rect 24912 19907 24970 19913
rect 24912 19873 24924 19907
rect 24958 19904 24970 19907
rect 25394 19904 25400 19916
rect 24958 19876 25400 19904
rect 24958 19873 24970 19876
rect 24912 19867 24970 19873
rect 25394 19864 25400 19876
rect 25452 19864 25458 19916
rect 10306 19836 10312 19848
rect 9496 19808 10312 19836
rect 10306 19796 10312 19808
rect 10364 19796 10370 19848
rect 12054 19836 12060 19848
rect 12015 19808 12060 19836
rect 12054 19796 12060 19808
rect 12112 19836 12118 19848
rect 12517 19839 12575 19845
rect 12517 19836 12529 19839
rect 12112 19808 12529 19836
rect 12112 19796 12118 19808
rect 12517 19805 12529 19808
rect 12563 19805 12575 19839
rect 15384 19836 15412 19864
rect 16470 19836 16476 19848
rect 12517 19799 12575 19805
rect 14832 19808 15412 19836
rect 16431 19808 16476 19836
rect 14832 19712 14860 19808
rect 16470 19796 16476 19808
rect 16528 19796 16534 19848
rect 21530 19836 21536 19848
rect 21491 19808 21536 19836
rect 21530 19796 21536 19808
rect 21588 19796 21594 19848
rect 24382 19728 24388 19780
rect 24440 19768 24446 19780
rect 24983 19771 25041 19777
rect 24983 19768 24995 19771
rect 24440 19740 24995 19768
rect 24440 19728 24446 19740
rect 24983 19737 24995 19740
rect 25029 19737 25041 19771
rect 24983 19731 25041 19737
rect 14633 19703 14691 19709
rect 14633 19669 14645 19703
rect 14679 19700 14691 19703
rect 14814 19700 14820 19712
rect 14679 19672 14820 19700
rect 14679 19669 14691 19672
rect 14633 19663 14691 19669
rect 14814 19660 14820 19672
rect 14872 19660 14878 19712
rect 21162 19660 21168 19712
rect 21220 19700 21226 19712
rect 21257 19703 21315 19709
rect 21257 19700 21269 19703
rect 21220 19672 21269 19700
rect 21220 19660 21226 19672
rect 21257 19669 21269 19672
rect 21303 19669 21315 19703
rect 23554 19700 23560 19712
rect 23515 19672 23560 19700
rect 21257 19663 21315 19669
rect 23554 19660 23560 19672
rect 23612 19660 23618 19712
rect 632 19610 26392 19632
rect 632 19558 5176 19610
rect 5228 19558 5240 19610
rect 5292 19558 5304 19610
rect 5356 19558 5368 19610
rect 5420 19558 14510 19610
rect 14562 19558 14574 19610
rect 14626 19558 14638 19610
rect 14690 19558 14702 19610
rect 14754 19558 23843 19610
rect 23895 19558 23907 19610
rect 23959 19558 23971 19610
rect 24023 19558 24035 19610
rect 24087 19558 26392 19610
rect 632 19536 26392 19558
rect 16194 19456 16200 19508
rect 16252 19496 16258 19508
rect 16473 19499 16531 19505
rect 16473 19496 16485 19499
rect 16252 19468 16485 19496
rect 16252 19456 16258 19468
rect 16473 19465 16485 19468
rect 16519 19496 16531 19499
rect 16746 19496 16752 19508
rect 16519 19468 16752 19496
rect 16519 19465 16531 19468
rect 16473 19459 16531 19465
rect 16746 19456 16752 19468
rect 16804 19456 16810 19508
rect 18862 19496 18868 19508
rect 18823 19468 18868 19496
rect 18862 19456 18868 19468
rect 18920 19456 18926 19508
rect 20978 19496 20984 19508
rect 20939 19468 20984 19496
rect 20978 19456 20984 19468
rect 21036 19456 21042 19508
rect 25394 19496 25400 19508
rect 25355 19468 25400 19496
rect 25394 19456 25400 19468
rect 25452 19456 25458 19508
rect 13342 19388 13348 19440
rect 13400 19428 13406 19440
rect 14906 19428 14912 19440
rect 13400 19400 14912 19428
rect 13400 19388 13406 19400
rect 14906 19388 14912 19400
rect 14964 19388 14970 19440
rect 16746 19320 16752 19372
rect 16804 19360 16810 19372
rect 17301 19363 17359 19369
rect 17301 19360 17313 19363
rect 16804 19332 17313 19360
rect 16804 19320 16810 19332
rect 17301 19329 17313 19332
rect 17347 19329 17359 19363
rect 23646 19360 23652 19372
rect 17301 19323 17359 19329
rect 23112 19332 23652 19360
rect 9205 19295 9263 19301
rect 9205 19261 9217 19295
rect 9251 19292 9263 19295
rect 9478 19292 9484 19304
rect 9251 19264 9484 19292
rect 9251 19261 9263 19264
rect 9205 19255 9263 19261
rect 9478 19252 9484 19264
rect 9536 19252 9542 19304
rect 9570 19252 9576 19304
rect 9628 19292 9634 19304
rect 9757 19295 9815 19301
rect 9757 19292 9769 19295
rect 9628 19264 9769 19292
rect 9628 19252 9634 19264
rect 9757 19261 9769 19264
rect 9803 19261 9815 19295
rect 11502 19292 11508 19304
rect 9757 19255 9815 19261
rect 10324 19264 11508 19292
rect 8837 19227 8895 19233
rect 8837 19193 8849 19227
rect 8883 19224 8895 19227
rect 9588 19224 9616 19252
rect 8883 19196 9616 19224
rect 8883 19193 8895 19196
rect 8837 19187 8895 19193
rect 10324 19168 10352 19264
rect 11502 19252 11508 19264
rect 11560 19252 11566 19304
rect 12054 19292 12060 19304
rect 12015 19264 12060 19292
rect 12054 19252 12060 19264
rect 12112 19252 12118 19304
rect 12517 19295 12575 19301
rect 12517 19261 12529 19295
rect 12563 19292 12575 19295
rect 13250 19292 13256 19304
rect 12563 19264 13256 19292
rect 12563 19261 12575 19264
rect 12517 19255 12575 19261
rect 12146 19224 12152 19236
rect 11152 19196 12152 19224
rect 9202 19116 9208 19168
rect 9260 19156 9266 19168
rect 9389 19159 9447 19165
rect 9389 19156 9401 19159
rect 9260 19128 9401 19156
rect 9260 19116 9266 19128
rect 9389 19125 9401 19128
rect 9435 19125 9447 19159
rect 10306 19156 10312 19168
rect 10267 19128 10312 19156
rect 9389 19119 9447 19125
rect 10306 19116 10312 19128
rect 10364 19116 10370 19168
rect 11152 19165 11180 19196
rect 12146 19184 12152 19196
rect 12204 19224 12210 19236
rect 12532 19224 12560 19255
rect 13250 19252 13256 19264
rect 13308 19252 13314 19304
rect 13710 19292 13716 19304
rect 13671 19264 13716 19292
rect 13710 19252 13716 19264
rect 13768 19252 13774 19304
rect 13986 19292 13992 19304
rect 13947 19264 13992 19292
rect 13986 19252 13992 19264
rect 14044 19292 14050 19304
rect 14541 19295 14599 19301
rect 14541 19292 14553 19295
rect 14044 19264 14553 19292
rect 14044 19252 14050 19264
rect 14541 19261 14553 19264
rect 14587 19261 14599 19295
rect 15274 19292 15280 19304
rect 15235 19264 15280 19292
rect 14541 19255 14599 19261
rect 15274 19252 15280 19264
rect 15332 19252 15338 19304
rect 15550 19252 15556 19304
rect 15608 19292 15614 19304
rect 15737 19295 15795 19301
rect 15737 19292 15749 19295
rect 15608 19264 15749 19292
rect 15608 19252 15614 19264
rect 15737 19261 15749 19264
rect 15783 19261 15795 19295
rect 15737 19255 15795 19261
rect 16013 19295 16071 19301
rect 16013 19261 16025 19295
rect 16059 19292 16071 19295
rect 16470 19292 16476 19304
rect 16059 19264 16476 19292
rect 16059 19261 16071 19264
rect 16013 19255 16071 19261
rect 16470 19252 16476 19264
rect 16528 19292 16534 19304
rect 16841 19295 16899 19301
rect 16841 19292 16853 19295
rect 16528 19264 16853 19292
rect 16528 19252 16534 19264
rect 16841 19261 16853 19264
rect 16887 19261 16899 19295
rect 16841 19255 16899 19261
rect 13158 19224 13164 19236
rect 12204 19196 12560 19224
rect 13119 19196 13164 19224
rect 12204 19184 12210 19196
rect 13158 19184 13164 19196
rect 13216 19184 13222 19236
rect 17316 19224 17344 19323
rect 17574 19292 17580 19304
rect 17535 19264 17580 19292
rect 17574 19252 17580 19264
rect 17632 19252 17638 19304
rect 18497 19295 18555 19301
rect 18497 19261 18509 19295
rect 18543 19292 18555 19295
rect 18862 19292 18868 19304
rect 18543 19264 18868 19292
rect 18543 19261 18555 19264
rect 18497 19255 18555 19261
rect 18862 19252 18868 19264
rect 18920 19252 18926 19304
rect 19782 19292 19788 19304
rect 19743 19264 19788 19292
rect 19782 19252 19788 19264
rect 19840 19252 19846 19304
rect 20702 19292 20708 19304
rect 20663 19264 20708 19292
rect 20702 19252 20708 19264
rect 20760 19252 20766 19304
rect 22266 19252 22272 19304
rect 22324 19292 22330 19304
rect 22637 19295 22695 19301
rect 22637 19292 22649 19295
rect 22324 19264 22649 19292
rect 22324 19252 22330 19264
rect 22637 19261 22649 19264
rect 22683 19292 22695 19295
rect 23112 19292 23140 19332
rect 23646 19320 23652 19332
rect 23704 19320 23710 19372
rect 24017 19363 24075 19369
rect 24017 19329 24029 19363
rect 24063 19360 24075 19363
rect 24198 19360 24204 19372
rect 24063 19332 24204 19360
rect 24063 19329 24075 19332
rect 24017 19323 24075 19329
rect 24198 19320 24204 19332
rect 24256 19360 24262 19372
rect 24474 19360 24480 19372
rect 24256 19332 24480 19360
rect 24256 19320 24262 19332
rect 24474 19320 24480 19332
rect 24532 19320 24538 19372
rect 22683 19264 23140 19292
rect 24912 19295 24970 19301
rect 22683 19261 22695 19264
rect 22637 19255 22695 19261
rect 24912 19261 24924 19295
rect 24958 19292 24970 19295
rect 25765 19295 25823 19301
rect 25765 19292 25777 19295
rect 24958 19264 25777 19292
rect 24958 19261 24970 19264
rect 24912 19255 24970 19261
rect 25765 19261 25777 19264
rect 25811 19292 25823 19295
rect 26866 19292 26872 19304
rect 25811 19264 26872 19292
rect 25811 19261 25823 19264
rect 25765 19255 25823 19261
rect 26866 19252 26872 19264
rect 26924 19252 26930 19304
rect 17898 19227 17956 19233
rect 17898 19224 17910 19227
rect 17316 19196 17910 19224
rect 17898 19193 17910 19196
rect 17944 19224 17956 19227
rect 18954 19224 18960 19236
rect 17944 19196 18960 19224
rect 17944 19193 17956 19196
rect 17898 19187 17956 19193
rect 18954 19184 18960 19196
rect 19012 19224 19018 19236
rect 19601 19227 19659 19233
rect 19601 19224 19613 19227
rect 19012 19196 19613 19224
rect 19012 19184 19018 19196
rect 19601 19193 19613 19196
rect 19647 19224 19659 19227
rect 20106 19227 20164 19233
rect 20106 19224 20118 19227
rect 19647 19196 20118 19224
rect 19647 19193 19659 19196
rect 19601 19187 19659 19193
rect 20106 19193 20118 19196
rect 20152 19224 20164 19227
rect 21070 19224 21076 19236
rect 20152 19196 21076 19224
rect 20152 19193 20164 19196
rect 20106 19187 20164 19193
rect 21070 19184 21076 19196
rect 21128 19224 21134 19236
rect 21533 19227 21591 19233
rect 21533 19224 21545 19227
rect 21128 19196 21545 19224
rect 21128 19184 21134 19196
rect 21533 19193 21545 19196
rect 21579 19193 21591 19227
rect 21533 19187 21591 19193
rect 22085 19227 22143 19233
rect 22085 19193 22097 19227
rect 22131 19224 22143 19227
rect 23370 19224 23376 19236
rect 22131 19196 23376 19224
rect 22131 19193 22143 19196
rect 22085 19187 22143 19193
rect 23370 19184 23376 19196
rect 23428 19184 23434 19236
rect 23465 19227 23523 19233
rect 23465 19193 23477 19227
rect 23511 19224 23523 19227
rect 23554 19224 23560 19236
rect 23511 19196 23560 19224
rect 23511 19193 23523 19196
rect 23465 19187 23523 19193
rect 10861 19159 10919 19165
rect 10861 19125 10873 19159
rect 10907 19156 10919 19159
rect 11137 19159 11195 19165
rect 11137 19156 11149 19159
rect 10907 19128 11149 19156
rect 10907 19125 10919 19128
rect 10861 19119 10919 19125
rect 11137 19125 11149 19128
rect 11183 19125 11195 19159
rect 11137 19119 11195 19125
rect 11962 19116 11968 19168
rect 12020 19156 12026 19168
rect 12057 19159 12115 19165
rect 12057 19156 12069 19159
rect 12020 19128 12069 19156
rect 12020 19116 12026 19128
rect 12057 19125 12069 19128
rect 12103 19125 12115 19159
rect 13618 19156 13624 19168
rect 13579 19128 13624 19156
rect 12057 19119 12115 19125
rect 13618 19116 13624 19128
rect 13676 19116 13682 19168
rect 21622 19116 21628 19168
rect 21680 19156 21686 19168
rect 21901 19159 21959 19165
rect 21901 19156 21913 19159
rect 21680 19128 21913 19156
rect 21680 19116 21686 19128
rect 21901 19125 21913 19128
rect 21947 19125 21959 19159
rect 21901 19119 21959 19125
rect 23005 19159 23063 19165
rect 23005 19125 23017 19159
rect 23051 19156 23063 19159
rect 23480 19156 23508 19187
rect 23554 19184 23560 19196
rect 23612 19184 23618 19236
rect 23051 19128 23508 19156
rect 23051 19125 23063 19128
rect 23005 19119 23063 19125
rect 24290 19116 24296 19168
rect 24348 19156 24354 19168
rect 24983 19159 25041 19165
rect 24983 19156 24995 19159
rect 24348 19128 24995 19156
rect 24348 19116 24354 19128
rect 24983 19125 24995 19128
rect 25029 19125 25041 19159
rect 24983 19119 25041 19125
rect 632 19066 26392 19088
rect 632 19014 9843 19066
rect 9895 19014 9907 19066
rect 9959 19014 9971 19066
rect 10023 19014 10035 19066
rect 10087 19014 19176 19066
rect 19228 19014 19240 19066
rect 19292 19014 19304 19066
rect 19356 19014 19368 19066
rect 19420 19014 26392 19066
rect 632 18992 26392 19014
rect 13253 18955 13311 18961
rect 13253 18921 13265 18955
rect 13299 18952 13311 18955
rect 13986 18952 13992 18964
rect 13299 18924 13992 18952
rect 13299 18921 13311 18924
rect 13253 18915 13311 18921
rect 13986 18912 13992 18924
rect 14044 18912 14050 18964
rect 17761 18955 17819 18961
rect 17761 18921 17773 18955
rect 17807 18952 17819 18955
rect 18494 18952 18500 18964
rect 17807 18924 18500 18952
rect 17807 18921 17819 18924
rect 17761 18915 17819 18921
rect 18494 18912 18500 18924
rect 18552 18912 18558 18964
rect 23370 18952 23376 18964
rect 23331 18924 23376 18952
rect 23370 18912 23376 18924
rect 23428 18912 23434 18964
rect 9202 18844 9208 18896
rect 9260 18884 9266 18896
rect 9846 18884 9852 18896
rect 9260 18856 9852 18884
rect 9260 18844 9266 18856
rect 9846 18844 9852 18856
rect 9904 18844 9910 18896
rect 9941 18887 9999 18893
rect 9941 18853 9953 18887
rect 9987 18884 9999 18887
rect 10214 18884 10220 18896
rect 9987 18856 10220 18884
rect 9987 18853 9999 18856
rect 9941 18847 9999 18853
rect 10214 18844 10220 18856
rect 10272 18844 10278 18896
rect 14906 18844 14912 18896
rect 14964 18884 14970 18896
rect 16565 18887 16623 18893
rect 14964 18856 15872 18884
rect 14964 18844 14970 18856
rect 15844 18828 15872 18856
rect 16565 18853 16577 18887
rect 16611 18884 16623 18887
rect 17574 18884 17580 18896
rect 16611 18856 17580 18884
rect 16611 18853 16623 18856
rect 16565 18847 16623 18853
rect 17574 18844 17580 18856
rect 17632 18844 17638 18896
rect 19509 18887 19567 18893
rect 19509 18853 19521 18887
rect 19555 18884 19567 18887
rect 19782 18884 19788 18896
rect 19555 18856 19788 18884
rect 19555 18853 19567 18856
rect 19509 18847 19567 18853
rect 19782 18844 19788 18856
rect 19840 18844 19846 18896
rect 21162 18884 21168 18896
rect 21123 18856 21168 18884
rect 21162 18844 21168 18856
rect 21220 18844 21226 18896
rect 23646 18884 23652 18896
rect 23607 18856 23652 18884
rect 23646 18844 23652 18856
rect 23704 18844 23710 18896
rect 24198 18884 24204 18896
rect 24159 18856 24204 18884
rect 24198 18844 24204 18856
rect 24256 18844 24262 18896
rect 15274 18816 15280 18828
rect 13912 18788 15280 18816
rect 10493 18751 10551 18757
rect 10493 18717 10505 18751
rect 10539 18748 10551 18751
rect 10674 18748 10680 18760
rect 10539 18720 10680 18748
rect 10539 18717 10551 18720
rect 10493 18711 10551 18717
rect 10674 18708 10680 18720
rect 10732 18708 10738 18760
rect 11318 18748 11324 18760
rect 11279 18720 11324 18748
rect 11318 18708 11324 18720
rect 11376 18708 11382 18760
rect 11962 18708 11968 18760
rect 12020 18748 12026 18760
rect 13710 18748 13716 18760
rect 12020 18720 13716 18748
rect 12020 18708 12026 18720
rect 13710 18708 13716 18720
rect 13768 18748 13774 18760
rect 13912 18757 13940 18788
rect 15274 18776 15280 18788
rect 15332 18776 15338 18828
rect 15826 18816 15832 18828
rect 15739 18788 15832 18816
rect 15826 18776 15832 18788
rect 15884 18776 15890 18828
rect 16289 18819 16347 18825
rect 16289 18785 16301 18819
rect 16335 18785 16347 18819
rect 18862 18816 18868 18828
rect 18823 18788 18868 18816
rect 16289 18779 16347 18785
rect 13897 18751 13955 18757
rect 13897 18748 13909 18751
rect 13768 18720 13909 18748
rect 13768 18708 13774 18720
rect 13897 18717 13909 18720
rect 13943 18717 13955 18751
rect 14630 18748 14636 18760
rect 14591 18720 14636 18748
rect 13897 18711 13955 18717
rect 14630 18708 14636 18720
rect 14688 18708 14694 18760
rect 16304 18748 16332 18779
rect 18862 18776 18868 18788
rect 18920 18776 18926 18828
rect 19046 18776 19052 18828
rect 19104 18816 19110 18828
rect 19233 18819 19291 18825
rect 19233 18816 19245 18819
rect 19104 18788 19245 18816
rect 19104 18776 19110 18788
rect 19233 18785 19245 18788
rect 19279 18785 19291 18819
rect 20702 18816 20708 18828
rect 20663 18788 20708 18816
rect 19233 18779 19291 18785
rect 20702 18776 20708 18788
rect 20760 18776 20766 18828
rect 20978 18816 20984 18828
rect 20939 18788 20984 18816
rect 20978 18776 20984 18788
rect 21036 18776 21042 18828
rect 16562 18748 16568 18760
rect 15660 18720 16568 18748
rect 9570 18612 9576 18624
rect 9531 18584 9576 18612
rect 9570 18572 9576 18584
rect 9628 18572 9634 18624
rect 10582 18572 10588 18624
rect 10640 18612 10646 18624
rect 10769 18615 10827 18621
rect 10769 18612 10781 18615
rect 10640 18584 10781 18612
rect 10640 18572 10646 18584
rect 10769 18581 10781 18584
rect 10815 18581 10827 18615
rect 10769 18575 10827 18581
rect 12054 18572 12060 18624
rect 12112 18612 12118 18624
rect 12333 18615 12391 18621
rect 12333 18612 12345 18615
rect 12112 18584 12345 18612
rect 12112 18572 12118 18584
rect 12333 18581 12345 18584
rect 12379 18581 12391 18615
rect 13618 18612 13624 18624
rect 13579 18584 13624 18612
rect 12333 18575 12391 18581
rect 13618 18572 13624 18584
rect 13676 18572 13682 18624
rect 15550 18572 15556 18624
rect 15608 18612 15614 18624
rect 15660 18621 15688 18720
rect 16562 18708 16568 18720
rect 16620 18708 16626 18760
rect 23554 18748 23560 18760
rect 23515 18720 23560 18748
rect 23554 18708 23560 18720
rect 23612 18708 23618 18760
rect 15645 18615 15703 18621
rect 15645 18612 15657 18615
rect 15608 18584 15657 18612
rect 15608 18572 15614 18584
rect 15645 18581 15657 18584
rect 15691 18581 15703 18615
rect 15645 18575 15703 18581
rect 21346 18572 21352 18624
rect 21404 18612 21410 18624
rect 21441 18615 21499 18621
rect 21441 18612 21453 18615
rect 21404 18584 21453 18612
rect 21404 18572 21410 18584
rect 21441 18581 21453 18584
rect 21487 18581 21499 18615
rect 21441 18575 21499 18581
rect 632 18522 26392 18544
rect 632 18470 5176 18522
rect 5228 18470 5240 18522
rect 5292 18470 5304 18522
rect 5356 18470 5368 18522
rect 5420 18470 14510 18522
rect 14562 18470 14574 18522
rect 14626 18470 14638 18522
rect 14690 18470 14702 18522
rect 14754 18470 23843 18522
rect 23895 18470 23907 18522
rect 23959 18470 23971 18522
rect 24023 18470 24035 18522
rect 24087 18470 26392 18522
rect 632 18448 26392 18470
rect 9846 18368 9852 18420
rect 9904 18408 9910 18420
rect 11321 18411 11379 18417
rect 11321 18408 11333 18411
rect 9904 18380 11333 18408
rect 9904 18368 9910 18380
rect 11321 18377 11333 18380
rect 11367 18377 11379 18411
rect 11321 18371 11379 18377
rect 13618 18368 13624 18420
rect 13676 18417 13682 18420
rect 13676 18411 13725 18417
rect 13676 18377 13679 18411
rect 13713 18377 13725 18411
rect 13986 18408 13992 18420
rect 13947 18380 13992 18408
rect 13676 18371 13725 18377
rect 13676 18368 13682 18371
rect 13986 18368 13992 18380
rect 14044 18368 14050 18420
rect 15826 18408 15832 18420
rect 15787 18380 15832 18408
rect 15826 18368 15832 18380
rect 15884 18408 15890 18420
rect 16102 18408 16108 18420
rect 15884 18380 16108 18408
rect 15884 18368 15890 18380
rect 16102 18368 16108 18380
rect 16160 18368 16166 18420
rect 16562 18408 16568 18420
rect 16523 18380 16568 18408
rect 16562 18368 16568 18380
rect 16620 18368 16626 18420
rect 18954 18368 18960 18420
rect 19012 18408 19018 18420
rect 19049 18411 19107 18417
rect 19049 18408 19061 18411
rect 19012 18380 19061 18408
rect 19012 18368 19018 18380
rect 19049 18377 19061 18380
rect 19095 18377 19107 18411
rect 20150 18408 20156 18420
rect 20111 18380 20156 18408
rect 19049 18371 19107 18377
rect 20150 18368 20156 18380
rect 20208 18368 20214 18420
rect 21070 18368 21076 18420
rect 21128 18408 21134 18420
rect 21165 18411 21223 18417
rect 21165 18408 21177 18411
rect 21128 18380 21177 18408
rect 21128 18368 21134 18380
rect 21165 18377 21177 18380
rect 21211 18408 21223 18411
rect 21622 18408 21628 18420
rect 21211 18380 21628 18408
rect 21211 18377 21223 18380
rect 21165 18371 21223 18377
rect 21622 18368 21628 18380
rect 21680 18368 21686 18420
rect 22266 18408 22272 18420
rect 22227 18380 22272 18408
rect 22266 18368 22272 18380
rect 22324 18368 22330 18420
rect 22637 18411 22695 18417
rect 22637 18377 22649 18411
rect 22683 18408 22695 18411
rect 23554 18408 23560 18420
rect 22683 18380 23560 18408
rect 22683 18377 22695 18380
rect 22637 18371 22695 18377
rect 23554 18368 23560 18380
rect 23612 18368 23618 18420
rect 10582 18340 10588 18352
rect 10416 18312 10588 18340
rect 10416 18281 10444 18312
rect 10582 18300 10588 18312
rect 10640 18300 10646 18352
rect 12606 18340 12612 18352
rect 12567 18312 12612 18340
rect 12606 18300 12612 18312
rect 12664 18300 12670 18352
rect 13805 18343 13863 18349
rect 13805 18309 13817 18343
rect 13851 18340 13863 18343
rect 13851 18312 14032 18340
rect 13851 18309 13863 18312
rect 13805 18303 13863 18309
rect 14004 18284 14032 18312
rect 10401 18275 10459 18281
rect 10401 18241 10413 18275
rect 10447 18241 10459 18275
rect 10674 18272 10680 18284
rect 10635 18244 10680 18272
rect 10401 18235 10459 18241
rect 10674 18232 10680 18244
rect 10732 18272 10738 18284
rect 12054 18272 12060 18284
rect 10732 18244 12060 18272
rect 10732 18232 10738 18244
rect 12054 18232 12060 18244
rect 12112 18232 12118 18284
rect 13434 18232 13440 18284
rect 13492 18272 13498 18284
rect 13897 18275 13955 18281
rect 13897 18272 13909 18275
rect 13492 18244 13909 18272
rect 13492 18232 13498 18244
rect 13897 18241 13909 18244
rect 13943 18241 13955 18275
rect 13897 18235 13955 18241
rect 13986 18232 13992 18284
rect 14044 18232 14050 18284
rect 19233 18275 19291 18281
rect 19233 18241 19245 18275
rect 19279 18272 19291 18275
rect 19506 18272 19512 18284
rect 19279 18244 19512 18272
rect 19279 18241 19291 18244
rect 19233 18235 19291 18241
rect 19506 18232 19512 18244
rect 19564 18232 19570 18284
rect 23572 18272 23600 18368
rect 24201 18275 24259 18281
rect 24201 18272 24213 18275
rect 23572 18244 24213 18272
rect 24201 18241 24213 18244
rect 24247 18272 24259 18275
rect 24382 18272 24388 18284
rect 24247 18244 24388 18272
rect 24247 18241 24259 18244
rect 24201 18235 24259 18241
rect 24382 18232 24388 18244
rect 24440 18232 24446 18284
rect 8653 18207 8711 18213
rect 8653 18173 8665 18207
rect 8699 18204 8711 18207
rect 9389 18207 9447 18213
rect 9389 18204 9401 18207
rect 8699 18176 9401 18204
rect 8699 18173 8711 18176
rect 8653 18167 8711 18173
rect 9389 18173 9401 18176
rect 9435 18204 9447 18207
rect 9849 18207 9907 18213
rect 9849 18204 9861 18207
rect 9435 18176 9861 18204
rect 9435 18173 9447 18176
rect 9389 18167 9447 18173
rect 9849 18173 9861 18176
rect 9895 18204 9907 18207
rect 10214 18204 10220 18216
rect 9895 18176 10220 18204
rect 9895 18173 9907 18176
rect 9849 18167 9907 18173
rect 10214 18164 10220 18176
rect 10272 18164 10278 18216
rect 18218 18204 18224 18216
rect 18131 18176 18224 18204
rect 18218 18164 18224 18176
rect 18276 18204 18282 18216
rect 18681 18207 18739 18213
rect 18681 18204 18693 18207
rect 18276 18176 18693 18204
rect 18276 18164 18282 18176
rect 18681 18173 18693 18176
rect 18727 18173 18739 18207
rect 21346 18204 21352 18216
rect 21307 18176 21352 18204
rect 18681 18167 18739 18173
rect 21346 18164 21352 18176
rect 21404 18164 21410 18216
rect 9481 18139 9539 18145
rect 9481 18105 9493 18139
rect 9527 18136 9539 18139
rect 10125 18139 10183 18145
rect 10125 18136 10137 18139
rect 9527 18108 10137 18136
rect 9527 18105 9539 18108
rect 9481 18099 9539 18105
rect 10125 18105 10137 18108
rect 10171 18105 10183 18139
rect 10125 18099 10183 18105
rect 10493 18139 10551 18145
rect 10493 18105 10505 18139
rect 10539 18105 10551 18139
rect 11778 18136 11784 18148
rect 11691 18108 11784 18136
rect 10493 18099 10551 18105
rect 10140 18068 10168 18099
rect 10508 18068 10536 18099
rect 11778 18096 11784 18108
rect 11836 18136 11842 18148
rect 12149 18139 12207 18145
rect 12149 18136 12161 18139
rect 11836 18108 12161 18136
rect 11836 18096 11842 18108
rect 12149 18105 12161 18108
rect 12195 18105 12207 18139
rect 12149 18099 12207 18105
rect 13069 18139 13127 18145
rect 13069 18105 13081 18139
rect 13115 18136 13127 18139
rect 13529 18139 13587 18145
rect 13529 18136 13541 18139
rect 13115 18108 13541 18136
rect 13115 18105 13127 18108
rect 13069 18099 13127 18105
rect 13529 18105 13541 18108
rect 13575 18136 13587 18139
rect 13710 18136 13716 18148
rect 13575 18108 13716 18136
rect 13575 18105 13587 18108
rect 13529 18099 13587 18105
rect 13710 18096 13716 18108
rect 13768 18096 13774 18148
rect 18954 18096 18960 18148
rect 19012 18136 19018 18148
rect 19554 18139 19612 18145
rect 19554 18136 19566 18139
rect 19012 18108 19566 18136
rect 19012 18096 19018 18108
rect 19554 18105 19566 18108
rect 19600 18105 19612 18139
rect 19554 18099 19612 18105
rect 21622 18096 21628 18148
rect 21680 18145 21686 18148
rect 21680 18139 21728 18145
rect 21680 18105 21682 18139
rect 21716 18105 21728 18139
rect 21680 18099 21728 18105
rect 23005 18139 23063 18145
rect 23005 18105 23017 18139
rect 23051 18136 23063 18139
rect 23922 18136 23928 18148
rect 23051 18108 23928 18136
rect 23051 18105 23063 18108
rect 23005 18099 23063 18105
rect 21680 18096 21686 18099
rect 23922 18096 23928 18108
rect 23980 18096 23986 18148
rect 24017 18139 24075 18145
rect 24017 18105 24029 18139
rect 24063 18105 24075 18139
rect 24017 18099 24075 18105
rect 13434 18068 13440 18080
rect 10140 18040 10536 18068
rect 13395 18040 13440 18068
rect 13434 18028 13440 18040
rect 13492 18028 13498 18080
rect 14538 18068 14544 18080
rect 14499 18040 14544 18068
rect 14538 18028 14544 18040
rect 14596 18028 14602 18080
rect 15001 18071 15059 18077
rect 15001 18037 15013 18071
rect 15047 18068 15059 18071
rect 15182 18068 15188 18080
rect 15047 18040 15188 18068
rect 15047 18037 15059 18040
rect 15001 18031 15059 18037
rect 15182 18028 15188 18040
rect 15240 18068 15246 18080
rect 15277 18071 15335 18077
rect 15277 18068 15289 18071
rect 15240 18040 15289 18068
rect 15240 18028 15246 18040
rect 15277 18037 15289 18040
rect 15323 18037 15335 18071
rect 16194 18068 16200 18080
rect 16155 18040 16200 18068
rect 15277 18031 15335 18037
rect 16194 18028 16200 18040
rect 16252 18028 16258 18080
rect 18129 18071 18187 18077
rect 18129 18037 18141 18071
rect 18175 18068 18187 18071
rect 18405 18071 18463 18077
rect 18405 18068 18417 18071
rect 18175 18040 18417 18068
rect 18175 18037 18187 18040
rect 18129 18031 18187 18037
rect 18405 18037 18417 18040
rect 18451 18068 18463 18071
rect 18862 18068 18868 18080
rect 18451 18040 18868 18068
rect 18451 18037 18463 18040
rect 18405 18031 18463 18037
rect 18862 18028 18868 18040
rect 18920 18028 18926 18080
rect 19046 18028 19052 18080
rect 19104 18068 19110 18080
rect 20429 18071 20487 18077
rect 20429 18068 20441 18071
rect 19104 18040 20441 18068
rect 19104 18028 19110 18040
rect 20429 18037 20441 18040
rect 20475 18037 20487 18071
rect 20429 18031 20487 18037
rect 20702 18028 20708 18080
rect 20760 18068 20766 18080
rect 20797 18071 20855 18077
rect 20797 18068 20809 18071
rect 20760 18040 20809 18068
rect 20760 18028 20766 18040
rect 20797 18037 20809 18040
rect 20843 18037 20855 18071
rect 23646 18068 23652 18080
rect 23607 18040 23652 18068
rect 20797 18031 20855 18037
rect 23646 18028 23652 18040
rect 23704 18068 23710 18080
rect 24032 18068 24060 18099
rect 23704 18040 24060 18068
rect 23704 18028 23710 18040
rect 632 17978 26392 18000
rect 632 17926 9843 17978
rect 9895 17926 9907 17978
rect 9959 17926 9971 17978
rect 10023 17926 10035 17978
rect 10087 17926 19176 17978
rect 19228 17926 19240 17978
rect 19292 17926 19304 17978
rect 19356 17926 19368 17978
rect 19420 17926 26392 17978
rect 632 17904 26392 17926
rect 10214 17824 10220 17876
rect 10272 17864 10278 17876
rect 10401 17867 10459 17873
rect 10401 17864 10413 17867
rect 10272 17836 10413 17864
rect 10272 17824 10278 17836
rect 10401 17833 10413 17836
rect 10447 17833 10459 17867
rect 13802 17864 13808 17876
rect 13763 17836 13808 17864
rect 10401 17827 10459 17833
rect 13802 17824 13808 17836
rect 13860 17824 13866 17876
rect 13986 17824 13992 17876
rect 14044 17864 14050 17876
rect 14538 17864 14544 17876
rect 14044 17836 14544 17864
rect 14044 17824 14050 17836
rect 14538 17824 14544 17836
rect 14596 17824 14602 17876
rect 16102 17824 16108 17876
rect 16160 17864 16166 17876
rect 16565 17867 16623 17873
rect 16565 17864 16577 17867
rect 16160 17836 16577 17864
rect 16160 17824 16166 17836
rect 16565 17833 16577 17836
rect 16611 17833 16623 17867
rect 23554 17864 23560 17876
rect 23515 17836 23560 17864
rect 16565 17827 16623 17833
rect 23554 17824 23560 17836
rect 23612 17824 23618 17876
rect 9662 17756 9668 17808
rect 9720 17796 9726 17808
rect 9802 17799 9860 17805
rect 9802 17796 9814 17799
rect 9720 17768 9814 17796
rect 9720 17756 9726 17768
rect 9802 17765 9814 17768
rect 9848 17765 9860 17799
rect 9802 17759 9860 17765
rect 11594 17756 11600 17808
rect 11652 17796 11658 17808
rect 11689 17799 11747 17805
rect 11689 17796 11701 17799
rect 11652 17768 11701 17796
rect 11652 17756 11658 17768
rect 11689 17765 11701 17768
rect 11735 17765 11747 17799
rect 11689 17759 11747 17765
rect 12241 17799 12299 17805
rect 12241 17765 12253 17799
rect 12287 17796 12299 17799
rect 12606 17796 12612 17808
rect 12287 17768 12612 17796
rect 12287 17765 12299 17768
rect 12241 17759 12299 17765
rect 12606 17756 12612 17768
rect 12664 17756 12670 17808
rect 13069 17799 13127 17805
rect 13069 17765 13081 17799
rect 13115 17796 13127 17799
rect 13618 17796 13624 17808
rect 13115 17768 13624 17796
rect 13115 17765 13127 17768
rect 13069 17759 13127 17765
rect 9478 17660 9484 17672
rect 9439 17632 9484 17660
rect 9478 17620 9484 17632
rect 9536 17620 9542 17672
rect 11318 17620 11324 17672
rect 11376 17660 11382 17672
rect 11597 17663 11655 17669
rect 11597 17660 11609 17663
rect 11376 17632 11609 17660
rect 11376 17620 11382 17632
rect 11597 17629 11609 17632
rect 11643 17629 11655 17663
rect 11597 17623 11655 17629
rect 10674 17524 10680 17536
rect 10635 17496 10680 17524
rect 10674 17484 10680 17496
rect 10732 17484 10738 17536
rect 12698 17524 12704 17536
rect 12659 17496 12704 17524
rect 12698 17484 12704 17496
rect 12756 17484 12762 17536
rect 12974 17484 12980 17536
rect 13032 17524 13038 17536
rect 13084 17524 13112 17759
rect 13618 17756 13624 17768
rect 13676 17796 13682 17808
rect 15550 17796 15556 17808
rect 13676 17768 15044 17796
rect 15511 17768 15556 17796
rect 13676 17756 13682 17768
rect 15016 17740 15044 17768
rect 15550 17756 15556 17768
rect 15608 17756 15614 17808
rect 18862 17756 18868 17808
rect 18920 17796 18926 17808
rect 19417 17799 19475 17805
rect 18920 17768 19276 17796
rect 18920 17756 18926 17768
rect 13161 17731 13219 17737
rect 13161 17697 13173 17731
rect 13207 17728 13219 17731
rect 13710 17728 13716 17740
rect 13207 17700 13716 17728
rect 13207 17697 13219 17700
rect 13161 17691 13219 17697
rect 13710 17688 13716 17700
rect 13768 17728 13774 17740
rect 14998 17737 15004 17740
rect 14817 17731 14875 17737
rect 13768 17700 14308 17728
rect 13768 17688 13774 17700
rect 13250 17620 13256 17672
rect 13308 17660 13314 17672
rect 13434 17660 13440 17672
rect 13308 17632 13440 17660
rect 13308 17620 13314 17632
rect 13434 17620 13440 17632
rect 13492 17660 13498 17672
rect 13529 17663 13587 17669
rect 13529 17660 13541 17663
rect 13492 17632 13541 17660
rect 13492 17620 13498 17632
rect 13529 17629 13541 17632
rect 13575 17629 13587 17663
rect 13529 17623 13587 17629
rect 13299 17527 13357 17533
rect 13299 17524 13311 17527
rect 13032 17496 13311 17524
rect 13032 17484 13038 17496
rect 13299 17493 13311 17496
rect 13345 17493 13357 17527
rect 13299 17487 13357 17493
rect 13434 17484 13440 17536
rect 13492 17524 13498 17536
rect 14170 17524 14176 17536
rect 13492 17496 14176 17524
rect 13492 17484 13498 17496
rect 14170 17484 14176 17496
rect 14228 17484 14234 17536
rect 14280 17533 14308 17700
rect 14817 17697 14829 17731
rect 14863 17697 14875 17731
rect 14817 17691 14875 17697
rect 14964 17731 15004 17737
rect 14964 17697 14976 17731
rect 15056 17728 15062 17740
rect 16378 17728 16384 17740
rect 15056 17700 15149 17728
rect 16339 17700 16384 17728
rect 14964 17691 15004 17697
rect 14832 17660 14860 17691
rect 14998 17688 15004 17691
rect 15056 17688 15062 17700
rect 16378 17688 16384 17700
rect 16436 17688 16442 17740
rect 18678 17728 18684 17740
rect 18639 17700 18684 17728
rect 18678 17688 18684 17700
rect 18736 17688 18742 17740
rect 19138 17728 19144 17740
rect 19099 17700 19144 17728
rect 19138 17688 19144 17700
rect 19196 17688 19202 17740
rect 19248 17728 19276 17768
rect 19417 17765 19429 17799
rect 19463 17796 19475 17799
rect 19506 17796 19512 17808
rect 19463 17768 19512 17796
rect 19463 17765 19475 17768
rect 19417 17759 19475 17765
rect 19506 17756 19512 17768
rect 19564 17796 19570 17808
rect 19693 17799 19751 17805
rect 19693 17796 19705 17799
rect 19564 17768 19705 17796
rect 19564 17756 19570 17768
rect 19693 17765 19705 17768
rect 19739 17765 19751 17799
rect 19693 17759 19751 17765
rect 21165 17799 21223 17805
rect 21165 17765 21177 17799
rect 21211 17796 21223 17799
rect 21530 17796 21536 17808
rect 21211 17768 21536 17796
rect 21211 17765 21223 17768
rect 21165 17759 21223 17765
rect 21530 17756 21536 17768
rect 21588 17756 21594 17808
rect 21622 17756 21628 17808
rect 21680 17796 21686 17808
rect 22314 17799 22372 17805
rect 22314 17796 22326 17799
rect 21680 17768 22326 17796
rect 21680 17756 21686 17768
rect 22314 17765 22326 17768
rect 22360 17765 22372 17799
rect 23925 17799 23983 17805
rect 23925 17796 23937 17799
rect 22314 17759 22372 17765
rect 22928 17768 23937 17796
rect 20705 17731 20763 17737
rect 20705 17728 20717 17731
rect 19248 17700 20717 17728
rect 20705 17697 20717 17700
rect 20751 17728 20763 17731
rect 20794 17728 20800 17740
rect 20751 17700 20800 17728
rect 20751 17697 20763 17700
rect 20705 17691 20763 17697
rect 20794 17688 20800 17700
rect 20852 17688 20858 17740
rect 20978 17688 20984 17740
rect 21036 17728 21042 17740
rect 22928 17737 22956 17768
rect 23925 17765 23937 17768
rect 23971 17796 23983 17799
rect 24198 17796 24204 17808
rect 23971 17768 24204 17796
rect 23971 17765 23983 17768
rect 23925 17759 23983 17765
rect 24198 17756 24204 17768
rect 24256 17756 24262 17808
rect 22913 17731 22971 17737
rect 21036 17700 21129 17728
rect 21036 17688 21042 17700
rect 22913 17697 22925 17731
rect 22959 17697 22971 17731
rect 22913 17691 22971 17697
rect 15182 17660 15188 17672
rect 14832 17632 14952 17660
rect 15143 17632 15188 17660
rect 14924 17604 14952 17632
rect 15182 17620 15188 17632
rect 15240 17620 15246 17672
rect 14906 17552 14912 17604
rect 14964 17592 14970 17604
rect 15921 17595 15979 17601
rect 15921 17592 15933 17595
rect 14964 17564 15933 17592
rect 14964 17552 14970 17564
rect 15921 17561 15933 17564
rect 15967 17561 15979 17595
rect 20996 17592 21024 17688
rect 21993 17663 22051 17669
rect 21993 17629 22005 17663
rect 22039 17660 22051 17663
rect 22358 17660 22364 17672
rect 22039 17632 22364 17660
rect 22039 17629 22051 17632
rect 21993 17623 22051 17629
rect 22358 17620 22364 17632
rect 22416 17620 22422 17672
rect 23833 17663 23891 17669
rect 23833 17629 23845 17663
rect 23879 17660 23891 17663
rect 24290 17660 24296 17672
rect 23879 17632 24296 17660
rect 23879 17629 23891 17632
rect 23833 17623 23891 17629
rect 24290 17620 24296 17632
rect 24348 17620 24354 17672
rect 21530 17592 21536 17604
rect 15921 17555 15979 17561
rect 20168 17564 21536 17592
rect 20168 17536 20196 17564
rect 21530 17552 21536 17564
rect 21588 17552 21594 17604
rect 24382 17592 24388 17604
rect 24343 17564 24388 17592
rect 24382 17552 24388 17564
rect 24440 17552 24446 17604
rect 14265 17527 14323 17533
rect 14265 17493 14277 17527
rect 14311 17524 14323 17527
rect 14354 17524 14360 17536
rect 14311 17496 14360 17524
rect 14311 17493 14323 17496
rect 14265 17487 14323 17493
rect 14354 17484 14360 17496
rect 14412 17484 14418 17536
rect 15093 17527 15151 17533
rect 15093 17493 15105 17527
rect 15139 17524 15151 17527
rect 15366 17524 15372 17536
rect 15139 17496 15372 17524
rect 15139 17493 15151 17496
rect 15093 17487 15151 17493
rect 15366 17484 15372 17496
rect 15424 17484 15430 17536
rect 16838 17524 16844 17536
rect 16799 17496 16844 17524
rect 16838 17484 16844 17496
rect 16896 17484 16902 17536
rect 17669 17527 17727 17533
rect 17669 17493 17681 17527
rect 17715 17524 17727 17527
rect 17850 17524 17856 17536
rect 17715 17496 17856 17524
rect 17715 17493 17727 17496
rect 17669 17487 17727 17493
rect 17850 17484 17856 17496
rect 17908 17484 17914 17536
rect 20150 17524 20156 17536
rect 20111 17496 20156 17524
rect 20150 17484 20156 17496
rect 20208 17484 20214 17536
rect 21438 17524 21444 17536
rect 21399 17496 21444 17524
rect 21438 17484 21444 17496
rect 21496 17484 21502 17536
rect 632 17434 26392 17456
rect 632 17382 5176 17434
rect 5228 17382 5240 17434
rect 5292 17382 5304 17434
rect 5356 17382 5368 17434
rect 5420 17382 14510 17434
rect 14562 17382 14574 17434
rect 14626 17382 14638 17434
rect 14690 17382 14702 17434
rect 14754 17382 23843 17434
rect 23895 17382 23907 17434
rect 23959 17382 23971 17434
rect 24023 17382 24035 17434
rect 24087 17382 26392 17434
rect 632 17360 26392 17382
rect 9662 17320 9668 17332
rect 9623 17292 9668 17320
rect 9662 17280 9668 17292
rect 9720 17320 9726 17332
rect 9849 17323 9907 17329
rect 9849 17320 9861 17323
rect 9720 17292 9861 17320
rect 9720 17280 9726 17292
rect 9849 17289 9861 17292
rect 9895 17320 9907 17323
rect 9941 17323 9999 17329
rect 9941 17320 9953 17323
rect 9895 17292 9953 17320
rect 9895 17289 9907 17292
rect 9849 17283 9907 17289
rect 9941 17289 9953 17292
rect 9987 17289 9999 17323
rect 11594 17320 11600 17332
rect 11555 17292 11600 17320
rect 9941 17283 9999 17289
rect 11594 17280 11600 17292
rect 11652 17280 11658 17332
rect 12974 17329 12980 17332
rect 12958 17323 12980 17329
rect 12958 17289 12970 17323
rect 12958 17283 12980 17289
rect 12974 17280 12980 17283
rect 13032 17280 13038 17332
rect 13342 17280 13348 17332
rect 13400 17320 13406 17332
rect 13437 17323 13495 17329
rect 13437 17320 13449 17323
rect 13400 17292 13449 17320
rect 13400 17280 13406 17292
rect 13437 17289 13449 17292
rect 13483 17289 13495 17323
rect 13437 17283 13495 17289
rect 14262 17280 14268 17332
rect 14320 17320 14326 17332
rect 15001 17323 15059 17329
rect 14320 17292 14768 17320
rect 14320 17280 14326 17292
rect 12514 17212 12520 17264
rect 12572 17252 12578 17264
rect 13069 17255 13127 17261
rect 13069 17252 13081 17255
rect 12572 17224 13081 17252
rect 12572 17212 12578 17224
rect 13069 17221 13081 17224
rect 13115 17252 13127 17255
rect 13986 17252 13992 17264
rect 13115 17224 13992 17252
rect 13115 17221 13127 17224
rect 13069 17215 13127 17221
rect 13986 17212 13992 17224
rect 14044 17252 14050 17264
rect 14630 17252 14636 17264
rect 14044 17224 14636 17252
rect 14044 17212 14050 17224
rect 14630 17212 14636 17224
rect 14688 17212 14694 17264
rect 14740 17252 14768 17292
rect 15001 17289 15013 17323
rect 15047 17320 15059 17323
rect 15918 17320 15924 17332
rect 15047 17292 15924 17320
rect 15047 17289 15059 17292
rect 15001 17283 15059 17289
rect 15918 17280 15924 17292
rect 15976 17280 15982 17332
rect 16565 17323 16623 17329
rect 16565 17289 16577 17323
rect 16611 17320 16623 17323
rect 18681 17323 18739 17329
rect 18681 17320 18693 17323
rect 16611 17292 18693 17320
rect 16611 17289 16623 17292
rect 16565 17283 16623 17289
rect 18681 17289 18693 17292
rect 18727 17320 18739 17323
rect 19138 17320 19144 17332
rect 18727 17292 19144 17320
rect 18727 17289 18739 17292
rect 18681 17283 18739 17289
rect 19138 17280 19144 17292
rect 19196 17280 19202 17332
rect 21530 17280 21536 17332
rect 21588 17320 21594 17332
rect 21625 17323 21683 17329
rect 21625 17320 21637 17323
rect 21588 17292 21637 17320
rect 21588 17280 21594 17292
rect 21625 17289 21637 17292
rect 21671 17289 21683 17323
rect 23646 17320 23652 17332
rect 23607 17292 23652 17320
rect 21625 17283 21683 17289
rect 23646 17280 23652 17292
rect 23704 17280 23710 17332
rect 24474 17280 24480 17332
rect 24532 17320 24538 17332
rect 25075 17323 25133 17329
rect 25075 17320 25087 17323
rect 24532 17292 25087 17320
rect 24532 17280 24538 17292
rect 25075 17289 25087 17292
rect 25121 17289 25133 17323
rect 25486 17320 25492 17332
rect 25447 17292 25492 17320
rect 25075 17283 25133 17289
rect 25486 17280 25492 17292
rect 25544 17280 25550 17332
rect 15366 17252 15372 17264
rect 14740 17224 15372 17252
rect 15366 17212 15372 17224
rect 15424 17212 15430 17264
rect 16194 17252 16200 17264
rect 16155 17224 16200 17252
rect 16194 17212 16200 17224
rect 16252 17212 16258 17264
rect 16378 17212 16384 17264
rect 16436 17252 16442 17264
rect 17025 17255 17083 17261
rect 17025 17252 17037 17255
rect 16436 17224 17037 17252
rect 16436 17212 16442 17224
rect 17025 17221 17037 17224
rect 17071 17252 17083 17255
rect 17206 17252 17212 17264
rect 17071 17224 17212 17252
rect 17071 17221 17083 17224
rect 17025 17215 17083 17221
rect 17206 17212 17212 17224
rect 17264 17252 17270 17264
rect 18218 17252 18224 17264
rect 17264 17224 18224 17252
rect 17264 17212 17270 17224
rect 18218 17212 18224 17224
rect 18276 17212 18282 17264
rect 9297 17187 9355 17193
rect 9297 17153 9309 17187
rect 9343 17184 9355 17187
rect 9478 17184 9484 17196
rect 9343 17156 9484 17184
rect 9343 17153 9355 17156
rect 9297 17147 9355 17153
rect 9478 17144 9484 17156
rect 9536 17144 9542 17196
rect 10398 17184 10404 17196
rect 9772 17156 10404 17184
rect 8837 17119 8895 17125
rect 8837 17085 8849 17119
rect 8883 17116 8895 17119
rect 9018 17116 9024 17128
rect 8883 17088 9024 17116
rect 8883 17085 8895 17088
rect 8837 17079 8895 17085
rect 9018 17076 9024 17088
rect 9076 17076 9082 17128
rect 9113 17119 9171 17125
rect 9113 17085 9125 17119
rect 9159 17116 9171 17119
rect 9772 17116 9800 17156
rect 10398 17144 10404 17156
rect 10456 17144 10462 17196
rect 12701 17187 12759 17193
rect 12701 17153 12713 17187
rect 12747 17184 12759 17187
rect 13161 17187 13219 17193
rect 13161 17184 13173 17187
rect 12747 17156 13173 17184
rect 12747 17153 12759 17156
rect 12701 17147 12759 17153
rect 13161 17153 13173 17156
rect 13207 17184 13219 17187
rect 13250 17184 13256 17196
rect 13207 17156 13256 17184
rect 13207 17153 13219 17156
rect 13161 17147 13219 17153
rect 13250 17144 13256 17156
rect 13308 17144 13314 17196
rect 14725 17187 14783 17193
rect 14725 17153 14737 17187
rect 14771 17184 14783 17187
rect 15182 17184 15188 17196
rect 14771 17156 15188 17184
rect 14771 17153 14783 17156
rect 14725 17147 14783 17153
rect 15182 17144 15188 17156
rect 15240 17184 15246 17196
rect 16289 17187 16347 17193
rect 16289 17184 16301 17187
rect 15240 17156 16301 17184
rect 15240 17144 15246 17156
rect 16289 17153 16301 17156
rect 16335 17184 16347 17187
rect 16838 17184 16844 17196
rect 16335 17156 16844 17184
rect 16335 17153 16347 17156
rect 16289 17147 16347 17153
rect 16838 17144 16844 17156
rect 16896 17144 16902 17196
rect 17669 17187 17727 17193
rect 17669 17153 17681 17187
rect 17715 17184 17727 17187
rect 17850 17184 17856 17196
rect 17715 17156 17856 17184
rect 17715 17153 17727 17156
rect 17669 17147 17727 17153
rect 17850 17144 17856 17156
rect 17908 17144 17914 17196
rect 17942 17144 17948 17196
rect 18000 17184 18006 17196
rect 21346 17184 21352 17196
rect 18000 17156 18045 17184
rect 21307 17156 21352 17184
rect 18000 17144 18006 17156
rect 21346 17144 21352 17156
rect 21404 17144 21410 17196
rect 9159 17088 9800 17116
rect 10125 17119 10183 17125
rect 9159 17085 9171 17088
rect 9113 17079 9171 17085
rect 10125 17085 10137 17119
rect 10171 17116 10183 17119
rect 10674 17116 10680 17128
rect 10171 17088 10680 17116
rect 10171 17085 10183 17088
rect 10125 17079 10183 17085
rect 8469 17051 8527 17057
rect 8469 17017 8481 17051
rect 8515 17048 8527 17051
rect 9128 17048 9156 17079
rect 10674 17076 10680 17088
rect 10732 17076 10738 17128
rect 11045 17119 11103 17125
rect 11045 17085 11057 17119
rect 11091 17116 11103 17119
rect 11778 17116 11784 17128
rect 11091 17088 11784 17116
rect 11091 17085 11103 17088
rect 11045 17079 11103 17085
rect 11778 17076 11784 17088
rect 11836 17076 11842 17128
rect 12333 17119 12391 17125
rect 12333 17085 12345 17119
rect 12379 17116 12391 17119
rect 13434 17116 13440 17128
rect 12379 17088 13440 17116
rect 12379 17085 12391 17088
rect 12333 17079 12391 17085
rect 13434 17076 13440 17088
rect 13492 17076 13498 17128
rect 14504 17119 14562 17125
rect 14504 17116 14516 17119
rect 14188 17088 14516 17116
rect 8515 17020 9156 17048
rect 9849 17051 9907 17057
rect 8515 17017 8527 17020
rect 8469 17011 8527 17017
rect 9849 17017 9861 17051
rect 9895 17048 9907 17051
rect 10446 17051 10504 17057
rect 10446 17048 10458 17051
rect 9895 17020 10458 17048
rect 9895 17017 9907 17020
rect 9849 17011 9907 17017
rect 10446 17017 10458 17020
rect 10492 17017 10504 17051
rect 10446 17011 10504 17017
rect 12698 17008 12704 17060
rect 12756 17048 12762 17060
rect 12793 17051 12851 17057
rect 12793 17048 12805 17051
rect 12756 17020 12805 17048
rect 12756 17008 12762 17020
rect 12793 17017 12805 17020
rect 12839 17048 12851 17051
rect 13158 17048 13164 17060
rect 12839 17020 13164 17048
rect 12839 17017 12851 17020
rect 12793 17011 12851 17017
rect 13158 17008 13164 17020
rect 13216 17008 13222 17060
rect 14188 16992 14216 17088
rect 14504 17085 14516 17088
rect 14550 17116 14562 17119
rect 15737 17119 15795 17125
rect 15737 17116 15749 17119
rect 14550 17088 15749 17116
rect 14550 17085 14562 17088
rect 14504 17079 14562 17085
rect 15737 17085 15749 17088
rect 15783 17116 15795 17119
rect 16068 17119 16126 17125
rect 16068 17116 16080 17119
rect 15783 17088 16080 17116
rect 15783 17085 15795 17088
rect 15737 17079 15795 17085
rect 16068 17085 16080 17088
rect 16114 17085 16126 17119
rect 16068 17079 16126 17085
rect 19141 17119 19199 17125
rect 19141 17085 19153 17119
rect 19187 17085 19199 17119
rect 19141 17079 19199 17085
rect 20153 17119 20211 17125
rect 20153 17085 20165 17119
rect 20199 17116 20211 17119
rect 20521 17119 20579 17125
rect 20521 17116 20533 17119
rect 20199 17088 20533 17116
rect 20199 17085 20211 17088
rect 20153 17079 20211 17085
rect 20521 17085 20533 17088
rect 20567 17116 20579 17119
rect 20794 17116 20800 17128
rect 20567 17088 20800 17116
rect 20567 17085 20579 17088
rect 20521 17079 20579 17085
rect 14354 17048 14360 17060
rect 14315 17020 14360 17048
rect 14354 17008 14360 17020
rect 14412 17008 14418 17060
rect 15642 17008 15648 17060
rect 15700 17048 15706 17060
rect 15921 17051 15979 17057
rect 15921 17048 15933 17051
rect 15700 17020 15933 17048
rect 15700 17008 15706 17020
rect 15921 17017 15933 17020
rect 15967 17017 15979 17051
rect 15921 17011 15979 17017
rect 17761 17051 17819 17057
rect 17761 17017 17773 17051
rect 17807 17017 17819 17051
rect 17761 17011 17819 17017
rect 13250 16940 13256 16992
rect 13308 16980 13314 16992
rect 13805 16983 13863 16989
rect 13805 16980 13817 16983
rect 13308 16952 13817 16980
rect 13308 16940 13314 16952
rect 13805 16949 13817 16952
rect 13851 16949 13863 16983
rect 14170 16980 14176 16992
rect 14131 16952 14176 16980
rect 13805 16943 13863 16949
rect 14170 16940 14176 16952
rect 14228 16940 14234 16992
rect 17298 16980 17304 16992
rect 17259 16952 17304 16980
rect 17298 16940 17304 16952
rect 17356 16980 17362 16992
rect 17776 16980 17804 17011
rect 18034 17008 18040 17060
rect 18092 17048 18098 17060
rect 19156 17048 19184 17079
rect 20794 17076 20800 17088
rect 20852 17076 20858 17128
rect 20886 17076 20892 17128
rect 20944 17116 20950 17128
rect 21073 17119 21131 17125
rect 21073 17116 21085 17119
rect 20944 17088 21085 17116
rect 20944 17076 20950 17088
rect 21073 17085 21085 17088
rect 21119 17116 21131 17119
rect 21438 17116 21444 17128
rect 21119 17088 21444 17116
rect 21119 17085 21131 17088
rect 21073 17079 21131 17085
rect 21438 17076 21444 17088
rect 21496 17076 21502 17128
rect 21622 17076 21628 17128
rect 21680 17116 21686 17128
rect 21993 17119 22051 17125
rect 21993 17116 22005 17119
rect 21680 17088 22005 17116
rect 21680 17076 21686 17088
rect 21993 17085 22005 17088
rect 22039 17085 22051 17119
rect 21993 17079 22051 17085
rect 23005 17119 23063 17125
rect 23005 17085 23017 17119
rect 23051 17116 23063 17119
rect 24017 17119 24075 17125
rect 24017 17116 24029 17119
rect 23051 17088 24029 17116
rect 23051 17085 23063 17088
rect 23005 17079 23063 17085
rect 24017 17085 24029 17088
rect 24063 17116 24075 17119
rect 24198 17116 24204 17128
rect 24063 17088 24204 17116
rect 24063 17085 24075 17088
rect 24017 17079 24075 17085
rect 24198 17076 24204 17088
rect 24256 17116 24262 17128
rect 24385 17119 24443 17125
rect 24385 17116 24397 17119
rect 24256 17088 24397 17116
rect 24256 17076 24262 17088
rect 24385 17085 24397 17088
rect 24431 17085 24443 17119
rect 24385 17079 24443 17085
rect 25004 17119 25062 17125
rect 25004 17085 25016 17119
rect 25050 17116 25062 17119
rect 25486 17116 25492 17128
rect 25050 17088 25492 17116
rect 25050 17085 25062 17088
rect 25004 17079 25062 17085
rect 25486 17076 25492 17088
rect 25544 17076 25550 17128
rect 19601 17051 19659 17057
rect 19601 17048 19613 17051
rect 18092 17020 19613 17048
rect 18092 17008 18098 17020
rect 19601 17017 19613 17020
rect 19647 17017 19659 17051
rect 19601 17011 19659 17017
rect 17356 16952 17804 16980
rect 17356 16940 17362 16952
rect 18678 16940 18684 16992
rect 18736 16980 18742 16992
rect 19325 16983 19383 16989
rect 19325 16980 19337 16983
rect 18736 16952 19337 16980
rect 18736 16940 18742 16952
rect 19325 16949 19337 16952
rect 19371 16980 19383 16983
rect 20702 16980 20708 16992
rect 19371 16952 20708 16980
rect 19371 16949 19383 16952
rect 19325 16943 19383 16949
rect 20702 16940 20708 16952
rect 20760 16940 20766 16992
rect 22358 16980 22364 16992
rect 22319 16952 22364 16980
rect 22358 16940 22364 16952
rect 22416 16940 22422 16992
rect 632 16890 26392 16912
rect 632 16838 9843 16890
rect 9895 16838 9907 16890
rect 9959 16838 9971 16890
rect 10023 16838 10035 16890
rect 10087 16838 19176 16890
rect 19228 16838 19240 16890
rect 19292 16838 19304 16890
rect 19356 16838 19368 16890
rect 19420 16838 26392 16890
rect 632 16816 26392 16838
rect 8653 16779 8711 16785
rect 8653 16745 8665 16779
rect 8699 16776 8711 16779
rect 9018 16776 9024 16788
rect 8699 16748 9024 16776
rect 8699 16745 8711 16748
rect 8653 16739 8711 16745
rect 9018 16736 9024 16748
rect 9076 16736 9082 16788
rect 9478 16776 9484 16788
rect 9439 16748 9484 16776
rect 9478 16736 9484 16748
rect 9536 16736 9542 16788
rect 11318 16776 11324 16788
rect 11279 16748 11324 16776
rect 11318 16736 11324 16748
rect 11376 16736 11382 16788
rect 11594 16736 11600 16788
rect 11652 16776 11658 16788
rect 11781 16779 11839 16785
rect 11781 16776 11793 16779
rect 11652 16748 11793 16776
rect 11652 16736 11658 16748
rect 11781 16745 11793 16748
rect 11827 16745 11839 16779
rect 11781 16739 11839 16745
rect 12885 16779 12943 16785
rect 12885 16745 12897 16779
rect 12931 16776 12943 16779
rect 12974 16776 12980 16788
rect 12931 16748 12980 16776
rect 12931 16745 12943 16748
rect 12885 16739 12943 16745
rect 12974 16736 12980 16748
rect 13032 16736 13038 16788
rect 13802 16776 13808 16788
rect 13763 16748 13808 16776
rect 13802 16736 13808 16748
rect 13860 16736 13866 16788
rect 14998 16776 15004 16788
rect 14959 16748 15004 16776
rect 14998 16736 15004 16748
rect 15056 16776 15062 16788
rect 15277 16779 15335 16785
rect 15277 16776 15289 16779
rect 15056 16748 15289 16776
rect 15056 16736 15062 16748
rect 15277 16745 15289 16748
rect 15323 16745 15335 16779
rect 18678 16776 18684 16788
rect 18639 16748 18684 16776
rect 15277 16739 15335 16745
rect 18678 16736 18684 16748
rect 18736 16736 18742 16788
rect 24109 16779 24167 16785
rect 24109 16745 24121 16779
rect 24155 16776 24167 16779
rect 24290 16776 24296 16788
rect 24155 16748 24296 16776
rect 24155 16745 24167 16748
rect 24109 16739 24167 16745
rect 24290 16736 24296 16748
rect 24348 16736 24354 16788
rect 10674 16708 10680 16720
rect 10635 16680 10680 16708
rect 10674 16668 10680 16680
rect 10732 16668 10738 16720
rect 12606 16668 12612 16720
rect 12664 16708 12670 16720
rect 14170 16708 14176 16720
rect 12664 16680 14176 16708
rect 12664 16668 12670 16680
rect 14170 16668 14176 16680
rect 14228 16708 14234 16720
rect 14228 16680 14860 16708
rect 14228 16668 14234 16680
rect 10214 16640 10220 16652
rect 10175 16612 10220 16640
rect 10214 16600 10220 16612
rect 10272 16600 10278 16652
rect 10398 16640 10404 16652
rect 10359 16612 10404 16640
rect 10398 16600 10404 16612
rect 10456 16600 10462 16652
rect 11778 16640 11784 16652
rect 11739 16612 11784 16640
rect 11778 16600 11784 16612
rect 11836 16600 11842 16652
rect 13158 16640 13164 16652
rect 13119 16612 13164 16640
rect 13158 16600 13164 16612
rect 13216 16600 13222 16652
rect 14832 16649 14860 16680
rect 14906 16668 14912 16720
rect 14964 16708 14970 16720
rect 15642 16708 15648 16720
rect 14964 16680 15648 16708
rect 14964 16668 14970 16680
rect 15642 16668 15648 16680
rect 15700 16668 15706 16720
rect 16010 16708 16016 16720
rect 15971 16680 16016 16708
rect 16010 16668 16016 16680
rect 16068 16668 16074 16720
rect 16105 16711 16163 16717
rect 16105 16677 16117 16711
rect 16151 16708 16163 16711
rect 16194 16708 16200 16720
rect 16151 16680 16200 16708
rect 16151 16677 16163 16680
rect 16105 16671 16163 16677
rect 16194 16668 16200 16680
rect 16252 16668 16258 16720
rect 17942 16708 17948 16720
rect 17408 16680 17948 16708
rect 14817 16643 14875 16649
rect 14817 16609 14829 16643
rect 14863 16640 14875 16643
rect 14998 16640 15004 16652
rect 14863 16612 15004 16640
rect 14863 16609 14875 16612
rect 14817 16603 14875 16609
rect 14998 16600 15004 16612
rect 15056 16600 15062 16652
rect 13250 16532 13256 16584
rect 13308 16572 13314 16584
rect 13529 16575 13587 16581
rect 13529 16572 13541 16575
rect 13308 16544 13541 16572
rect 13308 16532 13314 16544
rect 13529 16541 13541 16544
rect 13575 16541 13587 16575
rect 13529 16535 13587 16541
rect 16657 16575 16715 16581
rect 16657 16541 16669 16575
rect 16703 16572 16715 16575
rect 17408 16572 17436 16680
rect 17942 16668 17948 16680
rect 18000 16708 18006 16720
rect 18770 16708 18776 16720
rect 18000 16680 18776 16708
rect 18000 16668 18006 16680
rect 18770 16668 18776 16680
rect 18828 16668 18834 16720
rect 21349 16711 21407 16717
rect 21349 16677 21361 16711
rect 21395 16708 21407 16711
rect 22358 16708 22364 16720
rect 21395 16680 22364 16708
rect 21395 16677 21407 16680
rect 21349 16671 21407 16677
rect 22358 16668 22364 16680
rect 22416 16668 22422 16720
rect 23327 16711 23385 16717
rect 23327 16677 23339 16711
rect 23373 16708 23385 16711
rect 24382 16708 24388 16720
rect 23373 16680 24388 16708
rect 23373 16677 23385 16680
rect 23327 16671 23385 16677
rect 24382 16668 24388 16680
rect 24440 16668 24446 16720
rect 17574 16640 17580 16652
rect 17535 16612 17580 16640
rect 17574 16600 17580 16612
rect 17632 16640 17638 16652
rect 18034 16640 18040 16652
rect 17632 16612 18040 16640
rect 17632 16600 17638 16612
rect 18034 16600 18040 16612
rect 18092 16600 18098 16652
rect 18218 16640 18224 16652
rect 18179 16612 18224 16640
rect 18218 16600 18224 16612
rect 18276 16600 18282 16652
rect 19046 16640 19052 16652
rect 19007 16612 19052 16640
rect 19046 16600 19052 16612
rect 19104 16600 19110 16652
rect 20702 16640 20708 16652
rect 20663 16612 20708 16640
rect 20702 16600 20708 16612
rect 20760 16600 20766 16652
rect 20886 16600 20892 16652
rect 20944 16640 20950 16652
rect 21073 16643 21131 16649
rect 21073 16640 21085 16643
rect 20944 16612 21085 16640
rect 20944 16600 20950 16612
rect 21073 16609 21085 16612
rect 21119 16609 21131 16643
rect 21073 16603 21131 16609
rect 23186 16600 23192 16652
rect 23244 16649 23250 16652
rect 23244 16643 23282 16649
rect 23270 16640 23282 16643
rect 23649 16643 23707 16649
rect 23649 16640 23661 16643
rect 23270 16612 23661 16640
rect 23270 16609 23282 16612
rect 23244 16603 23282 16609
rect 23649 16609 23661 16612
rect 23695 16609 23707 16643
rect 23649 16603 23707 16609
rect 23244 16600 23250 16603
rect 23738 16600 23744 16652
rect 23796 16640 23802 16652
rect 24290 16649 24296 16652
rect 24268 16643 24296 16649
rect 24268 16640 24280 16643
rect 23796 16612 24280 16640
rect 23796 16600 23802 16612
rect 24268 16609 24280 16612
rect 24268 16603 24296 16609
rect 24290 16600 24296 16603
rect 24348 16600 24354 16652
rect 16703 16544 17436 16572
rect 16703 16541 16715 16544
rect 16657 16535 16715 16541
rect 13437 16507 13495 16513
rect 13437 16473 13449 16507
rect 13483 16504 13495 16507
rect 14262 16504 14268 16516
rect 13483 16476 14268 16504
rect 13483 16473 13495 16476
rect 13437 16467 13495 16473
rect 14262 16464 14268 16476
rect 14320 16464 14326 16516
rect 12974 16396 12980 16448
rect 13032 16436 13038 16448
rect 13299 16439 13357 16445
rect 13299 16436 13311 16439
rect 13032 16408 13311 16436
rect 13032 16396 13038 16408
rect 13299 16405 13311 16408
rect 13345 16405 13357 16439
rect 14354 16436 14360 16448
rect 14315 16408 14360 16436
rect 13299 16399 13357 16405
rect 14354 16396 14360 16408
rect 14412 16396 14418 16448
rect 23002 16396 23008 16448
rect 23060 16436 23066 16448
rect 24339 16439 24397 16445
rect 24339 16436 24351 16439
rect 23060 16408 24351 16436
rect 23060 16396 23066 16408
rect 24339 16405 24351 16408
rect 24385 16405 24397 16439
rect 24339 16399 24397 16405
rect 632 16346 26392 16368
rect 632 16294 5176 16346
rect 5228 16294 5240 16346
rect 5292 16294 5304 16346
rect 5356 16294 5368 16346
rect 5420 16294 14510 16346
rect 14562 16294 14574 16346
rect 14626 16294 14638 16346
rect 14690 16294 14702 16346
rect 14754 16294 23843 16346
rect 23895 16294 23907 16346
rect 23959 16294 23971 16346
rect 24023 16294 24035 16346
rect 24087 16294 26392 16346
rect 632 16272 26392 16294
rect 9202 16192 9208 16244
rect 9260 16232 9266 16244
rect 9665 16235 9723 16241
rect 9665 16232 9677 16235
rect 9260 16204 9677 16232
rect 9260 16192 9266 16204
rect 9665 16201 9677 16204
rect 9711 16201 9723 16235
rect 9665 16195 9723 16201
rect 10214 16192 10220 16244
rect 10272 16232 10278 16244
rect 10309 16235 10367 16241
rect 10309 16232 10321 16235
rect 10272 16204 10321 16232
rect 10272 16192 10278 16204
rect 10309 16201 10321 16204
rect 10355 16201 10367 16235
rect 10766 16232 10772 16244
rect 10727 16204 10772 16232
rect 10309 16195 10367 16201
rect 10766 16192 10772 16204
rect 10824 16192 10830 16244
rect 11597 16235 11655 16241
rect 11597 16201 11609 16235
rect 11643 16232 11655 16235
rect 11778 16232 11784 16244
rect 11643 16204 11784 16232
rect 11643 16201 11655 16204
rect 11597 16195 11655 16201
rect 11778 16192 11784 16204
rect 11836 16192 11842 16244
rect 12885 16235 12943 16241
rect 12885 16201 12897 16235
rect 12931 16232 12943 16235
rect 12974 16232 12980 16244
rect 12931 16204 12980 16232
rect 12931 16201 12943 16204
rect 12885 16195 12943 16201
rect 12974 16192 12980 16204
rect 13032 16232 13038 16244
rect 14078 16232 14084 16244
rect 13032 16204 14084 16232
rect 13032 16192 13038 16204
rect 14078 16192 14084 16204
rect 14136 16232 14142 16244
rect 14219 16235 14277 16241
rect 14219 16232 14231 16235
rect 14136 16204 14231 16232
rect 14136 16192 14142 16204
rect 14219 16201 14231 16204
rect 14265 16201 14277 16235
rect 14219 16195 14277 16201
rect 14725 16235 14783 16241
rect 14725 16201 14737 16235
rect 14771 16232 14783 16235
rect 14814 16232 14820 16244
rect 14771 16204 14820 16232
rect 14771 16201 14783 16204
rect 14725 16195 14783 16201
rect 14814 16192 14820 16204
rect 14872 16192 14878 16244
rect 14998 16192 15004 16244
rect 15056 16232 15062 16244
rect 15093 16235 15151 16241
rect 15093 16232 15105 16235
rect 15056 16204 15105 16232
rect 15056 16192 15062 16204
rect 15093 16201 15105 16204
rect 15139 16201 15151 16235
rect 18862 16232 18868 16244
rect 18823 16204 18868 16232
rect 15093 16195 15151 16201
rect 18862 16192 18868 16204
rect 18920 16232 18926 16244
rect 24290 16232 24296 16244
rect 18920 16204 19552 16232
rect 24251 16204 24296 16232
rect 18920 16192 18926 16204
rect 14357 16167 14415 16173
rect 14357 16164 14369 16167
rect 14280 16136 14369 16164
rect 14280 16108 14308 16136
rect 14357 16133 14369 16136
rect 14403 16133 14415 16167
rect 14357 16127 14415 16133
rect 13434 16056 13440 16108
rect 13492 16096 13498 16108
rect 13621 16099 13679 16105
rect 13621 16096 13633 16099
rect 13492 16068 13633 16096
rect 13492 16056 13498 16068
rect 13621 16065 13633 16068
rect 13667 16096 13679 16099
rect 13989 16099 14047 16105
rect 13989 16096 14001 16099
rect 13667 16068 14001 16096
rect 13667 16065 13679 16068
rect 13621 16059 13679 16065
rect 13989 16065 14001 16068
rect 14035 16096 14047 16099
rect 14262 16096 14268 16108
rect 14035 16068 14268 16096
rect 14035 16065 14047 16068
rect 13989 16059 14047 16065
rect 14262 16056 14268 16068
rect 14320 16056 14326 16108
rect 14449 16099 14507 16105
rect 14449 16065 14461 16099
rect 14495 16096 14507 16099
rect 15182 16096 15188 16108
rect 14495 16068 15188 16096
rect 14495 16065 14507 16068
rect 14449 16059 14507 16065
rect 15182 16056 15188 16068
rect 15240 16056 15246 16108
rect 16657 16099 16715 16105
rect 16657 16065 16669 16099
rect 16703 16096 16715 16099
rect 17298 16096 17304 16108
rect 16703 16068 17304 16096
rect 16703 16065 16715 16068
rect 16657 16059 16715 16065
rect 17298 16056 17304 16068
rect 17356 16056 17362 16108
rect 19524 16105 19552 16204
rect 24290 16192 24296 16204
rect 24348 16192 24354 16244
rect 24934 16232 24940 16244
rect 24895 16204 24940 16232
rect 24934 16192 24940 16204
rect 24992 16192 24998 16244
rect 19509 16099 19567 16105
rect 19509 16065 19521 16099
rect 19555 16065 19567 16099
rect 20150 16096 20156 16108
rect 20111 16068 20156 16096
rect 19509 16059 19567 16065
rect 20150 16056 20156 16068
rect 20208 16056 20214 16108
rect 22637 16099 22695 16105
rect 22637 16065 22649 16099
rect 22683 16096 22695 16099
rect 23281 16099 23339 16105
rect 23281 16096 23293 16099
rect 22683 16068 23293 16096
rect 22683 16065 22695 16068
rect 22637 16059 22695 16065
rect 23281 16065 23293 16068
rect 23327 16096 23339 16099
rect 25026 16096 25032 16108
rect 23327 16068 25032 16096
rect 23327 16065 23339 16068
rect 23281 16059 23339 16065
rect 25026 16056 25032 16068
rect 25084 16056 25090 16108
rect 9481 16031 9539 16037
rect 9481 15997 9493 16031
rect 9527 16028 9539 16031
rect 9527 16000 10076 16028
rect 9527 15997 9539 16000
rect 9481 15991 9539 15997
rect 10048 15901 10076 16000
rect 16194 15988 16200 16040
rect 16252 16028 16258 16040
rect 16565 16031 16623 16037
rect 16565 16028 16577 16031
rect 16252 16000 16577 16028
rect 16252 15988 16258 16000
rect 16565 15997 16577 16000
rect 16611 16028 16623 16031
rect 16933 16031 16991 16037
rect 16933 16028 16945 16031
rect 16611 16000 16945 16028
rect 16611 15997 16623 16000
rect 16565 15991 16623 15997
rect 16933 15997 16945 16000
rect 16979 15997 16991 16031
rect 16933 15991 16991 15997
rect 17942 15988 17948 16040
rect 18000 16028 18006 16040
rect 18497 16031 18555 16037
rect 18497 16028 18509 16031
rect 18000 16000 18509 16028
rect 18000 15988 18006 16000
rect 18497 15997 18509 16000
rect 18543 16028 18555 16031
rect 18543 16000 19368 16028
rect 18543 15997 18555 16000
rect 18497 15991 18555 15997
rect 14081 15963 14139 15969
rect 14081 15929 14093 15963
rect 14127 15960 14139 15963
rect 14354 15960 14360 15972
rect 14127 15932 14360 15960
rect 14127 15929 14139 15932
rect 14081 15923 14139 15929
rect 14354 15920 14360 15932
rect 14412 15920 14418 15972
rect 18586 15960 18592 15972
rect 18547 15932 18592 15960
rect 18586 15920 18592 15932
rect 18644 15920 18650 15972
rect 10033 15895 10091 15901
rect 10033 15861 10045 15895
rect 10079 15892 10091 15895
rect 10214 15892 10220 15904
rect 10079 15864 10220 15892
rect 10079 15861 10091 15864
rect 10033 15855 10091 15861
rect 10214 15852 10220 15864
rect 10272 15852 10278 15904
rect 12514 15892 12520 15904
rect 12475 15864 12520 15892
rect 12514 15852 12520 15864
rect 12572 15852 12578 15904
rect 13250 15892 13256 15904
rect 13211 15864 13256 15892
rect 13250 15852 13256 15864
rect 13308 15852 13314 15904
rect 15182 15852 15188 15904
rect 15240 15892 15246 15904
rect 15461 15895 15519 15901
rect 15461 15892 15473 15895
rect 15240 15864 15473 15892
rect 15240 15852 15246 15864
rect 15461 15861 15473 15864
rect 15507 15861 15519 15895
rect 17298 15892 17304 15904
rect 17259 15864 17304 15892
rect 15461 15855 15519 15861
rect 17298 15852 17304 15864
rect 17356 15852 17362 15904
rect 19340 15901 19368 16000
rect 24382 15988 24388 16040
rect 24440 16028 24446 16040
rect 24753 16031 24811 16037
rect 24753 16028 24765 16031
rect 24440 16000 24765 16028
rect 24440 15988 24446 16000
rect 24753 15997 24765 16000
rect 24799 16028 24811 16031
rect 25305 16031 25363 16037
rect 25305 16028 25317 16031
rect 24799 16000 25317 16028
rect 24799 15997 24811 16000
rect 24753 15991 24811 15997
rect 25305 15997 25317 16000
rect 25351 15997 25363 16031
rect 25305 15991 25363 15997
rect 19601 15963 19659 15969
rect 19601 15929 19613 15963
rect 19647 15929 19659 15963
rect 20702 15960 20708 15972
rect 20615 15932 20708 15960
rect 19601 15923 19659 15929
rect 19325 15895 19383 15901
rect 19325 15861 19337 15895
rect 19371 15892 19383 15895
rect 19616 15892 19644 15923
rect 20702 15920 20708 15932
rect 20760 15960 20766 15972
rect 21438 15960 21444 15972
rect 20760 15932 21444 15960
rect 20760 15920 20766 15932
rect 21438 15920 21444 15932
rect 21496 15920 21502 15972
rect 23370 15920 23376 15972
rect 23428 15960 23434 15972
rect 23922 15960 23928 15972
rect 23428 15932 23473 15960
rect 23883 15932 23928 15960
rect 23428 15920 23434 15932
rect 23922 15920 23928 15932
rect 23980 15920 23986 15972
rect 19371 15864 19644 15892
rect 19371 15861 19383 15864
rect 19325 15855 19383 15861
rect 20886 15852 20892 15904
rect 20944 15892 20950 15904
rect 20981 15895 21039 15901
rect 20981 15892 20993 15895
rect 20944 15864 20993 15892
rect 20944 15852 20950 15864
rect 20981 15861 20993 15864
rect 21027 15861 21039 15895
rect 20981 15855 21039 15861
rect 23005 15895 23063 15901
rect 23005 15861 23017 15895
rect 23051 15892 23063 15895
rect 23388 15892 23416 15920
rect 23051 15864 23416 15892
rect 23051 15861 23063 15864
rect 23005 15855 23063 15861
rect 632 15802 26392 15824
rect 632 15750 9843 15802
rect 9895 15750 9907 15802
rect 9959 15750 9971 15802
rect 10023 15750 10035 15802
rect 10087 15750 19176 15802
rect 19228 15750 19240 15802
rect 19292 15750 19304 15802
rect 19356 15750 19368 15802
rect 19420 15750 26392 15802
rect 632 15728 26392 15750
rect 14078 15688 14084 15700
rect 14039 15660 14084 15688
rect 14078 15648 14084 15660
rect 14136 15648 14142 15700
rect 15829 15691 15887 15697
rect 15829 15657 15841 15691
rect 15875 15688 15887 15691
rect 16194 15688 16200 15700
rect 15875 15660 16200 15688
rect 15875 15657 15887 15660
rect 15829 15651 15887 15657
rect 16194 15648 16200 15660
rect 16252 15648 16258 15700
rect 17577 15691 17635 15697
rect 17577 15657 17589 15691
rect 17623 15688 17635 15691
rect 17942 15688 17948 15700
rect 17623 15660 17948 15688
rect 17623 15657 17635 15660
rect 17577 15651 17635 15657
rect 17942 15648 17948 15660
rect 18000 15648 18006 15700
rect 18218 15688 18224 15700
rect 18179 15660 18224 15688
rect 18218 15648 18224 15660
rect 18276 15648 18282 15700
rect 23370 15648 23376 15700
rect 23428 15688 23434 15700
rect 23557 15691 23615 15697
rect 23557 15688 23569 15691
rect 23428 15660 23569 15688
rect 23428 15648 23434 15660
rect 23557 15657 23569 15660
rect 23603 15657 23615 15691
rect 23557 15651 23615 15657
rect 15271 15623 15329 15629
rect 15271 15589 15283 15623
rect 15317 15620 15329 15623
rect 15734 15620 15740 15632
rect 15317 15592 15740 15620
rect 15317 15589 15329 15592
rect 15271 15583 15329 15589
rect 15734 15580 15740 15592
rect 15792 15620 15798 15632
rect 15792 15592 16056 15620
rect 15792 15580 15798 15592
rect 16028 15552 16056 15592
rect 16102 15580 16108 15632
rect 16160 15620 16166 15632
rect 16473 15623 16531 15629
rect 16473 15620 16485 15623
rect 16160 15592 16485 15620
rect 16160 15580 16166 15592
rect 16473 15589 16485 15592
rect 16519 15589 16531 15623
rect 16978 15623 17036 15629
rect 16978 15620 16990 15623
rect 16473 15583 16531 15589
rect 16764 15592 16990 15620
rect 16764 15564 16792 15592
rect 16978 15589 16990 15592
rect 17024 15589 17036 15623
rect 18586 15620 18592 15632
rect 18547 15592 18592 15620
rect 16978 15583 17036 15589
rect 18586 15580 18592 15592
rect 18644 15580 18650 15632
rect 19141 15623 19199 15629
rect 19141 15589 19153 15623
rect 19187 15620 19199 15623
rect 20150 15620 20156 15632
rect 19187 15592 20156 15620
rect 19187 15589 19199 15592
rect 19141 15583 19199 15589
rect 20150 15580 20156 15592
rect 20208 15580 20214 15632
rect 21898 15620 21904 15632
rect 21859 15592 21904 15620
rect 21898 15580 21904 15592
rect 21956 15580 21962 15632
rect 22453 15623 22511 15629
rect 22453 15589 22465 15623
rect 22499 15620 22511 15623
rect 23186 15620 23192 15632
rect 22499 15592 23192 15620
rect 22499 15589 22511 15592
rect 22453 15583 22511 15589
rect 23186 15580 23192 15592
rect 23244 15620 23250 15632
rect 23922 15620 23928 15632
rect 23244 15592 23928 15620
rect 23244 15580 23250 15592
rect 23922 15580 23928 15592
rect 23980 15580 23986 15632
rect 16746 15552 16752 15564
rect 16028 15524 16752 15552
rect 16746 15512 16752 15524
rect 16804 15512 16810 15564
rect 23370 15552 23376 15564
rect 23331 15524 23376 15552
rect 23370 15512 23376 15524
rect 23428 15512 23434 15564
rect 24842 15512 24848 15564
rect 24900 15561 24906 15564
rect 24900 15555 24938 15561
rect 24926 15521 24938 15555
rect 24900 15515 24938 15521
rect 24900 15512 24906 15515
rect 14906 15484 14912 15496
rect 14867 15456 14912 15484
rect 14906 15444 14912 15456
rect 14964 15444 14970 15496
rect 16654 15484 16660 15496
rect 16615 15456 16660 15484
rect 16654 15444 16660 15456
rect 16712 15444 16718 15496
rect 18497 15487 18555 15493
rect 18497 15453 18509 15487
rect 18543 15484 18555 15487
rect 18770 15484 18776 15496
rect 18543 15456 18776 15484
rect 18543 15453 18555 15456
rect 18497 15447 18555 15453
rect 18770 15444 18776 15456
rect 18828 15444 18834 15496
rect 20429 15487 20487 15493
rect 20429 15453 20441 15487
rect 20475 15484 20487 15487
rect 20518 15484 20524 15496
rect 20475 15456 20524 15484
rect 20475 15453 20487 15456
rect 20429 15447 20487 15453
rect 20518 15444 20524 15456
rect 20576 15444 20582 15496
rect 21806 15484 21812 15496
rect 21767 15456 21812 15484
rect 21806 15444 21812 15456
rect 21864 15444 21870 15496
rect 13158 15308 13164 15360
rect 13216 15348 13222 15360
rect 13253 15351 13311 15357
rect 13253 15348 13265 15351
rect 13216 15320 13265 15348
rect 13216 15308 13222 15320
rect 13253 15317 13265 15320
rect 13299 15348 13311 15351
rect 13342 15348 13348 15360
rect 13299 15320 13348 15348
rect 13299 15317 13311 15320
rect 13253 15311 13311 15317
rect 13342 15308 13348 15320
rect 13400 15308 13406 15360
rect 14354 15308 14360 15360
rect 14412 15348 14418 15360
rect 14449 15351 14507 15357
rect 14449 15348 14461 15351
rect 14412 15320 14461 15348
rect 14412 15308 14418 15320
rect 14449 15317 14461 15320
rect 14495 15317 14507 15351
rect 14449 15311 14507 15317
rect 18954 15308 18960 15360
rect 19012 15348 19018 15360
rect 19417 15351 19475 15357
rect 19417 15348 19429 15351
rect 19012 15320 19429 15348
rect 19012 15308 19018 15320
rect 19417 15317 19429 15320
rect 19463 15317 19475 15351
rect 20978 15348 20984 15360
rect 20939 15320 20984 15348
rect 19417 15311 19475 15317
rect 20978 15308 20984 15320
rect 21036 15308 21042 15360
rect 24290 15308 24296 15360
rect 24348 15348 24354 15360
rect 24983 15351 25041 15357
rect 24983 15348 24995 15351
rect 24348 15320 24995 15348
rect 24348 15308 24354 15320
rect 24983 15317 24995 15320
rect 25029 15317 25041 15351
rect 24983 15311 25041 15317
rect 632 15258 26392 15280
rect 632 15206 5176 15258
rect 5228 15206 5240 15258
rect 5292 15206 5304 15258
rect 5356 15206 5368 15258
rect 5420 15206 14510 15258
rect 14562 15206 14574 15258
rect 14626 15206 14638 15258
rect 14690 15206 14702 15258
rect 14754 15206 23843 15258
rect 23895 15206 23907 15258
rect 23959 15206 23971 15258
rect 24023 15206 24035 15258
rect 24087 15206 26392 15258
rect 632 15184 26392 15206
rect 15734 15144 15740 15156
rect 15695 15116 15740 15144
rect 15734 15104 15740 15116
rect 15792 15104 15798 15156
rect 16746 15144 16752 15156
rect 16707 15116 16752 15144
rect 16746 15104 16752 15116
rect 16804 15104 16810 15156
rect 17206 15144 17212 15156
rect 17167 15116 17212 15144
rect 17206 15104 17212 15116
rect 17264 15104 17270 15156
rect 18586 15144 18592 15156
rect 18547 15116 18592 15144
rect 18586 15104 18592 15116
rect 18644 15104 18650 15156
rect 19046 15144 19052 15156
rect 19007 15116 19052 15144
rect 19046 15104 19052 15116
rect 19104 15104 19110 15156
rect 21898 15144 21904 15156
rect 21811 15116 21904 15144
rect 21898 15104 21904 15116
rect 21956 15144 21962 15156
rect 22269 15147 22327 15153
rect 22269 15144 22281 15147
rect 21956 15116 22281 15144
rect 21956 15104 21962 15116
rect 22269 15113 22281 15116
rect 22315 15144 22327 15147
rect 23370 15144 23376 15156
rect 22315 15116 23376 15144
rect 22315 15113 22327 15116
rect 22269 15107 22327 15113
rect 23370 15104 23376 15116
rect 23428 15104 23434 15156
rect 24017 15147 24075 15153
rect 24017 15113 24029 15147
rect 24063 15144 24075 15147
rect 24290 15144 24296 15156
rect 24063 15116 24296 15144
rect 24063 15113 24075 15116
rect 24017 15107 24075 15113
rect 21806 15036 21812 15088
rect 21864 15076 21870 15088
rect 22545 15079 22603 15085
rect 22545 15076 22557 15079
rect 21864 15048 22557 15076
rect 21864 15036 21870 15048
rect 22545 15045 22557 15048
rect 22591 15045 22603 15079
rect 22545 15039 22603 15045
rect 17666 15008 17672 15020
rect 17627 14980 17672 15008
rect 17666 14968 17672 14980
rect 17724 14968 17730 15020
rect 14265 14943 14323 14949
rect 14265 14909 14277 14943
rect 14311 14940 14323 14943
rect 14354 14940 14360 14952
rect 14311 14912 14360 14940
rect 14311 14909 14323 14912
rect 14265 14903 14323 14909
rect 14354 14900 14360 14912
rect 14412 14940 14418 14952
rect 14630 14940 14636 14952
rect 14412 14912 14636 14940
rect 14412 14900 14418 14912
rect 14630 14900 14636 14912
rect 14688 14900 14694 14952
rect 14817 14943 14875 14949
rect 14817 14909 14829 14943
rect 14863 14940 14875 14943
rect 14998 14940 15004 14952
rect 14863 14912 15004 14940
rect 14863 14909 14875 14912
rect 14817 14903 14875 14909
rect 14832 14872 14860 14903
rect 14998 14900 15004 14912
rect 15056 14900 15062 14952
rect 15182 14940 15188 14952
rect 15095 14912 15188 14940
rect 15182 14900 15188 14912
rect 15240 14940 15246 14952
rect 16289 14943 16347 14949
rect 15240 14912 16240 14940
rect 15240 14900 15246 14912
rect 13912 14844 14860 14872
rect 13912 14816 13940 14844
rect 14906 14832 14912 14884
rect 14964 14872 14970 14884
rect 16105 14875 16163 14881
rect 16105 14872 16117 14875
rect 14964 14844 16117 14872
rect 14964 14832 14970 14844
rect 16105 14841 16117 14844
rect 16151 14841 16163 14875
rect 16105 14835 16163 14841
rect 13894 14804 13900 14816
rect 13855 14776 13900 14804
rect 13894 14764 13900 14776
rect 13952 14764 13958 14816
rect 15458 14804 15464 14816
rect 15419 14776 15464 14804
rect 15458 14764 15464 14776
rect 15516 14764 15522 14816
rect 16212 14804 16240 14912
rect 16289 14909 16301 14943
rect 16335 14940 16347 14943
rect 17206 14940 17212 14952
rect 16335 14912 17212 14940
rect 16335 14909 16347 14912
rect 16289 14903 16347 14909
rect 17206 14900 17212 14912
rect 17264 14900 17270 14952
rect 20978 14940 20984 14952
rect 20939 14912 20984 14940
rect 20978 14900 20984 14912
rect 21036 14940 21042 14952
rect 22082 14940 22088 14952
rect 21036 14912 22088 14940
rect 21036 14900 21042 14912
rect 22082 14900 22088 14912
rect 22140 14900 22146 14952
rect 24124 14949 24152 15116
rect 24290 15104 24296 15116
rect 24348 15104 24354 15156
rect 24109 14943 24167 14949
rect 24109 14909 24121 14943
rect 24155 14909 24167 14943
rect 24109 14903 24167 14909
rect 17758 14832 17764 14884
rect 17816 14872 17822 14884
rect 18313 14875 18371 14881
rect 17816 14844 17861 14872
rect 17816 14832 17822 14844
rect 18313 14841 18325 14875
rect 18359 14872 18371 14875
rect 18954 14872 18960 14884
rect 18359 14844 18960 14872
rect 18359 14841 18371 14844
rect 18313 14835 18371 14841
rect 18954 14832 18960 14844
rect 19012 14872 19018 14884
rect 19233 14875 19291 14881
rect 19233 14872 19245 14875
rect 19012 14844 19245 14872
rect 19012 14832 19018 14844
rect 19233 14841 19245 14844
rect 19279 14841 19291 14875
rect 19233 14835 19291 14841
rect 19325 14875 19383 14881
rect 19325 14841 19337 14875
rect 19371 14841 19383 14875
rect 19325 14835 19383 14841
rect 19877 14875 19935 14881
rect 19877 14841 19889 14875
rect 19923 14872 19935 14875
rect 20702 14872 20708 14884
rect 19923 14844 20708 14872
rect 19923 14841 19935 14844
rect 19877 14835 19935 14841
rect 16473 14807 16531 14813
rect 16473 14804 16485 14807
rect 16212 14776 16485 14804
rect 16473 14773 16485 14776
rect 16519 14773 16531 14807
rect 16473 14767 16531 14773
rect 19046 14764 19052 14816
rect 19104 14804 19110 14816
rect 19340 14804 19368 14835
rect 20702 14832 20708 14844
rect 20760 14832 20766 14884
rect 20889 14875 20947 14881
rect 20889 14841 20901 14875
rect 20935 14872 20947 14875
rect 21343 14875 21401 14881
rect 21343 14872 21355 14875
rect 20935 14844 21355 14872
rect 20935 14841 20947 14844
rect 20889 14835 20947 14841
rect 21343 14841 21355 14844
rect 21389 14872 21401 14875
rect 21530 14872 21536 14884
rect 21389 14844 21536 14872
rect 21389 14841 21401 14844
rect 21343 14835 21401 14841
rect 21530 14832 21536 14844
rect 21588 14832 21594 14884
rect 19104 14776 19368 14804
rect 19104 14764 19110 14776
rect 24198 14764 24204 14816
rect 24256 14804 24262 14816
rect 24293 14807 24351 14813
rect 24293 14804 24305 14807
rect 24256 14776 24305 14804
rect 24256 14764 24262 14776
rect 24293 14773 24305 14776
rect 24339 14773 24351 14807
rect 24842 14804 24848 14816
rect 24803 14776 24848 14804
rect 24293 14767 24351 14773
rect 24842 14764 24848 14776
rect 24900 14764 24906 14816
rect 632 14714 26392 14736
rect 632 14662 9843 14714
rect 9895 14662 9907 14714
rect 9959 14662 9971 14714
rect 10023 14662 10035 14714
rect 10087 14662 19176 14714
rect 19228 14662 19240 14714
rect 19292 14662 19304 14714
rect 19356 14662 19368 14714
rect 19420 14662 26392 14714
rect 632 14640 26392 14662
rect 13894 14560 13900 14612
rect 13952 14600 13958 14612
rect 13989 14603 14047 14609
rect 13989 14600 14001 14603
rect 13952 14572 14001 14600
rect 13952 14560 13958 14572
rect 13989 14569 14001 14572
rect 14035 14569 14047 14603
rect 14906 14600 14912 14612
rect 14867 14572 14912 14600
rect 13989 14563 14047 14569
rect 14906 14560 14912 14572
rect 14964 14560 14970 14612
rect 15458 14560 15464 14612
rect 15516 14600 15522 14612
rect 16654 14600 16660 14612
rect 15516 14572 16660 14600
rect 15516 14560 15522 14572
rect 16654 14560 16660 14572
rect 16712 14560 16718 14612
rect 17669 14603 17727 14609
rect 17669 14569 17681 14603
rect 17715 14600 17727 14603
rect 17758 14600 17764 14612
rect 17715 14572 17764 14600
rect 17715 14569 17727 14572
rect 17669 14563 17727 14569
rect 17758 14560 17764 14572
rect 17816 14560 17822 14612
rect 22082 14600 22088 14612
rect 22043 14572 22088 14600
rect 22082 14560 22088 14572
rect 22140 14560 22146 14612
rect 23186 14600 23192 14612
rect 23147 14572 23192 14600
rect 23186 14560 23192 14572
rect 23244 14560 23250 14612
rect 14449 14535 14507 14541
rect 14449 14501 14461 14535
rect 14495 14532 14507 14535
rect 15182 14532 15188 14544
rect 14495 14504 15188 14532
rect 14495 14501 14507 14504
rect 14449 14495 14507 14501
rect 15182 14492 15188 14504
rect 15240 14492 15246 14544
rect 16746 14492 16752 14544
rect 16804 14532 16810 14544
rect 17942 14532 17948 14544
rect 16804 14504 17948 14532
rect 16804 14492 16810 14504
rect 17942 14492 17948 14504
rect 18000 14532 18006 14544
rect 18082 14535 18140 14541
rect 18082 14532 18094 14535
rect 18000 14504 18094 14532
rect 18000 14492 18006 14504
rect 18082 14501 18094 14504
rect 18128 14501 18140 14535
rect 20610 14532 20616 14544
rect 20571 14504 20616 14532
rect 18082 14495 18140 14501
rect 20610 14492 20616 14504
rect 20668 14492 20674 14544
rect 14630 14424 14636 14476
rect 14688 14464 14694 14476
rect 14909 14467 14967 14473
rect 14909 14464 14921 14467
rect 14688 14436 14921 14464
rect 14688 14424 14694 14436
rect 14909 14433 14921 14436
rect 14955 14433 14967 14467
rect 14909 14427 14967 14433
rect 14924 14396 14952 14427
rect 14998 14424 15004 14476
rect 15056 14464 15062 14476
rect 15277 14467 15335 14473
rect 15277 14464 15289 14467
rect 15056 14436 15289 14464
rect 15056 14424 15062 14436
rect 15277 14433 15289 14436
rect 15323 14433 15335 14467
rect 15642 14464 15648 14476
rect 15603 14436 15648 14464
rect 15277 14427 15335 14433
rect 15642 14424 15648 14436
rect 15700 14424 15706 14476
rect 21438 14424 21444 14476
rect 21496 14464 21502 14476
rect 21993 14467 22051 14473
rect 21993 14464 22005 14467
rect 21496 14436 22005 14464
rect 21496 14424 21502 14436
rect 21993 14433 22005 14436
rect 22039 14464 22051 14467
rect 22358 14464 22364 14476
rect 22039 14436 22364 14464
rect 22039 14433 22051 14436
rect 21993 14427 22051 14433
rect 22358 14424 22364 14436
rect 22416 14424 22422 14476
rect 22453 14467 22511 14473
rect 22453 14433 22465 14467
rect 22499 14433 22511 14467
rect 24198 14464 24204 14476
rect 24159 14436 24204 14464
rect 22453 14427 22511 14433
rect 15734 14396 15740 14408
rect 14924 14368 15740 14396
rect 15734 14356 15740 14368
rect 15792 14356 15798 14408
rect 17761 14399 17819 14405
rect 17761 14365 17773 14399
rect 17807 14396 17819 14399
rect 18126 14396 18132 14408
rect 17807 14368 18132 14396
rect 17807 14365 17819 14368
rect 17761 14359 17819 14365
rect 18126 14356 18132 14368
rect 18184 14356 18190 14408
rect 20518 14396 20524 14408
rect 20479 14368 20524 14396
rect 20518 14356 20524 14368
rect 20576 14356 20582 14408
rect 20702 14356 20708 14408
rect 20760 14396 20766 14408
rect 20797 14399 20855 14405
rect 20797 14396 20809 14399
rect 20760 14368 20809 14396
rect 20760 14356 20766 14368
rect 20797 14365 20809 14368
rect 20843 14365 20855 14399
rect 20797 14359 20855 14365
rect 21806 14356 21812 14408
rect 21864 14396 21870 14408
rect 22468 14396 22496 14427
rect 24198 14424 24204 14436
rect 24256 14424 24262 14476
rect 23554 14396 23560 14408
rect 21864 14368 22496 14396
rect 23515 14368 23560 14396
rect 21864 14356 21870 14368
rect 23554 14356 23560 14368
rect 23612 14356 23618 14408
rect 18681 14263 18739 14269
rect 18681 14229 18693 14263
rect 18727 14260 18739 14263
rect 19138 14260 19144 14272
rect 18727 14232 19144 14260
rect 18727 14229 18739 14232
rect 18681 14223 18739 14229
rect 19138 14220 19144 14232
rect 19196 14220 19202 14272
rect 21346 14220 21352 14272
rect 21404 14260 21410 14272
rect 21441 14263 21499 14269
rect 21441 14260 21453 14263
rect 21404 14232 21453 14260
rect 21404 14220 21410 14232
rect 21441 14229 21453 14232
rect 21487 14229 21499 14263
rect 21441 14223 21499 14229
rect 632 14170 26392 14192
rect 632 14118 5176 14170
rect 5228 14118 5240 14170
rect 5292 14118 5304 14170
rect 5356 14118 5368 14170
rect 5420 14118 14510 14170
rect 14562 14118 14574 14170
rect 14626 14118 14638 14170
rect 14690 14118 14702 14170
rect 14754 14118 23843 14170
rect 23895 14118 23907 14170
rect 23959 14118 23971 14170
rect 24023 14118 24035 14170
rect 24087 14118 26392 14170
rect 632 14096 26392 14118
rect 13161 14059 13219 14065
rect 13161 14025 13173 14059
rect 13207 14056 13219 14059
rect 14354 14056 14360 14068
rect 13207 14028 14360 14056
rect 13207 14025 13219 14028
rect 13161 14019 13219 14025
rect 14354 14016 14360 14028
rect 14412 14016 14418 14068
rect 15734 14056 15740 14068
rect 15695 14028 15740 14056
rect 15734 14016 15740 14028
rect 15792 14016 15798 14068
rect 17853 14059 17911 14065
rect 17853 14025 17865 14059
rect 17899 14056 17911 14059
rect 17942 14056 17948 14068
rect 17899 14028 17948 14056
rect 17899 14025 17911 14028
rect 17853 14019 17911 14025
rect 17942 14016 17948 14028
rect 18000 14016 18006 14068
rect 20518 14016 20524 14068
rect 20576 14056 20582 14068
rect 20797 14059 20855 14065
rect 20797 14056 20809 14059
rect 20576 14028 20809 14056
rect 20576 14016 20582 14028
rect 20797 14025 20809 14028
rect 20843 14025 20855 14059
rect 20797 14019 20855 14025
rect 22269 14059 22327 14065
rect 22269 14025 22281 14059
rect 22315 14056 22327 14059
rect 23005 14059 23063 14065
rect 23005 14056 23017 14059
rect 22315 14028 23017 14056
rect 22315 14025 22327 14028
rect 22269 14019 22327 14025
rect 23005 14025 23017 14028
rect 23051 14056 23063 14059
rect 23370 14056 23376 14068
rect 23051 14028 23376 14056
rect 23051 14025 23063 14028
rect 23005 14019 23063 14025
rect 23370 14016 23376 14028
rect 23428 14056 23434 14068
rect 24198 14056 24204 14068
rect 23428 14028 24204 14056
rect 23428 14016 23434 14028
rect 24198 14016 24204 14028
rect 24256 14016 24262 14068
rect 13342 13948 13348 14000
rect 13400 13988 13406 14000
rect 14173 13991 14231 13997
rect 14173 13988 14185 13991
rect 13400 13960 14185 13988
rect 13400 13948 13406 13960
rect 12977 13855 13035 13861
rect 12977 13821 12989 13855
rect 13023 13852 13035 13855
rect 13158 13852 13164 13864
rect 13023 13824 13164 13852
rect 13023 13821 13035 13824
rect 12977 13815 13035 13821
rect 13158 13812 13164 13824
rect 13216 13852 13222 13864
rect 13437 13855 13495 13861
rect 13437 13852 13449 13855
rect 13216 13824 13449 13852
rect 13216 13812 13222 13824
rect 13437 13821 13449 13824
rect 13483 13821 13495 13855
rect 13437 13815 13495 13821
rect 12330 13744 12336 13796
rect 12388 13784 12394 13796
rect 13544 13784 13572 13960
rect 14173 13957 14185 13960
rect 14219 13988 14231 13991
rect 14262 13988 14268 14000
rect 14219 13960 14268 13988
rect 14219 13957 14231 13960
rect 14173 13951 14231 13957
rect 14262 13948 14268 13960
rect 14320 13948 14326 14000
rect 22358 13948 22364 14000
rect 22416 13988 22422 14000
rect 22545 13991 22603 13997
rect 22545 13988 22557 13991
rect 22416 13960 22557 13988
rect 22416 13948 22422 13960
rect 22545 13957 22557 13960
rect 22591 13957 22603 13991
rect 22545 13951 22603 13957
rect 23186 13948 23192 14000
rect 23244 13948 23250 14000
rect 19785 13923 19843 13929
rect 14096 13892 15228 13920
rect 14096 13864 14124 13892
rect 13897 13855 13955 13861
rect 13897 13821 13909 13855
rect 13943 13852 13955 13855
rect 14078 13852 14084 13864
rect 13943 13824 14084 13852
rect 13943 13821 13955 13824
rect 13897 13815 13955 13821
rect 14078 13812 14084 13824
rect 14136 13812 14142 13864
rect 14262 13812 14268 13864
rect 14320 13852 14326 13864
rect 14357 13855 14415 13861
rect 14357 13852 14369 13855
rect 14320 13824 14369 13852
rect 14320 13812 14326 13824
rect 14357 13821 14369 13824
rect 14403 13852 14415 13855
rect 14722 13852 14728 13864
rect 14403 13824 14728 13852
rect 14403 13821 14415 13824
rect 14357 13815 14415 13821
rect 14722 13812 14728 13824
rect 14780 13812 14786 13864
rect 14998 13852 15004 13864
rect 14959 13824 15004 13852
rect 14998 13812 15004 13824
rect 15056 13812 15062 13864
rect 15200 13861 15228 13892
rect 19785 13889 19797 13923
rect 19831 13920 19843 13923
rect 20429 13923 20487 13929
rect 20429 13920 20441 13923
rect 19831 13892 20441 13920
rect 19831 13889 19843 13892
rect 19785 13883 19843 13889
rect 20429 13889 20441 13892
rect 20475 13920 20487 13923
rect 20610 13920 20616 13932
rect 20475 13892 20616 13920
rect 20475 13889 20487 13892
rect 20429 13883 20487 13889
rect 20610 13880 20616 13892
rect 20668 13880 20674 13932
rect 21257 13923 21315 13929
rect 21257 13889 21269 13923
rect 21303 13920 21315 13923
rect 23204 13920 23232 13948
rect 23281 13923 23339 13929
rect 23281 13920 23293 13923
rect 21303 13892 21484 13920
rect 23204 13892 23293 13920
rect 21303 13889 21315 13892
rect 21257 13883 21315 13889
rect 15185 13855 15243 13861
rect 15185 13821 15197 13855
rect 15231 13852 15243 13855
rect 15642 13852 15648 13864
rect 15231 13824 15648 13852
rect 15231 13821 15243 13824
rect 15185 13815 15243 13821
rect 15642 13812 15648 13824
rect 15700 13852 15706 13864
rect 16105 13855 16163 13861
rect 16105 13852 16117 13855
rect 15700 13824 16117 13852
rect 15700 13812 15706 13824
rect 16105 13821 16117 13824
rect 16151 13821 16163 13855
rect 16473 13855 16531 13861
rect 16473 13852 16485 13855
rect 16105 13815 16163 13821
rect 16212 13824 16485 13852
rect 12388 13756 13572 13784
rect 15016 13784 15044 13812
rect 16212 13784 16240 13824
rect 16473 13821 16485 13824
rect 16519 13821 16531 13855
rect 18126 13852 18132 13864
rect 18087 13824 18132 13852
rect 16473 13815 16531 13821
rect 18126 13812 18132 13824
rect 18184 13812 18190 13864
rect 18957 13855 19015 13861
rect 18957 13821 18969 13855
rect 19003 13852 19015 13855
rect 19138 13852 19144 13864
rect 19003 13824 19144 13852
rect 19003 13821 19015 13824
rect 18957 13815 19015 13821
rect 19138 13812 19144 13824
rect 19196 13812 19202 13864
rect 21346 13852 21352 13864
rect 21307 13824 21352 13852
rect 21346 13812 21352 13824
rect 21404 13812 21410 13864
rect 15016 13756 16240 13784
rect 21456 13784 21484 13892
rect 23281 13889 23293 13892
rect 23327 13889 23339 13923
rect 23281 13883 23339 13889
rect 21530 13784 21536 13796
rect 21456 13756 21536 13784
rect 12388 13744 12394 13756
rect 21530 13744 21536 13756
rect 21588 13784 21594 13796
rect 21670 13787 21728 13793
rect 21670 13784 21682 13787
rect 21588 13756 21682 13784
rect 21588 13744 21594 13756
rect 21670 13753 21682 13756
rect 21716 13753 21728 13787
rect 21670 13747 21728 13753
rect 23370 13744 23376 13796
rect 23428 13784 23434 13796
rect 23922 13784 23928 13796
rect 23428 13756 23473 13784
rect 23883 13756 23928 13784
rect 23428 13744 23434 13756
rect 23922 13744 23928 13756
rect 23980 13744 23986 13796
rect 15458 13716 15464 13728
rect 15419 13688 15464 13716
rect 15458 13676 15464 13688
rect 15516 13676 15522 13728
rect 23462 13676 23468 13728
rect 23520 13716 23526 13728
rect 24753 13719 24811 13725
rect 24753 13716 24765 13719
rect 23520 13688 24765 13716
rect 23520 13676 23526 13688
rect 24753 13685 24765 13688
rect 24799 13685 24811 13719
rect 24753 13679 24811 13685
rect 632 13626 26392 13648
rect 632 13574 9843 13626
rect 9895 13574 9907 13626
rect 9959 13574 9971 13626
rect 10023 13574 10035 13626
rect 10087 13574 19176 13626
rect 19228 13574 19240 13626
rect 19292 13574 19304 13626
rect 19356 13574 19368 13626
rect 19420 13574 26392 13626
rect 632 13552 26392 13574
rect 12330 13512 12336 13524
rect 12291 13484 12336 13512
rect 12330 13472 12336 13484
rect 12388 13472 12394 13524
rect 15458 13472 15464 13524
rect 15516 13512 15522 13524
rect 16197 13515 16255 13521
rect 16197 13512 16209 13515
rect 15516 13484 16209 13512
rect 15516 13472 15522 13484
rect 16197 13481 16209 13484
rect 16243 13481 16255 13515
rect 16197 13475 16255 13481
rect 22315 13515 22373 13521
rect 22315 13481 22327 13515
rect 22361 13512 22373 13515
rect 24934 13512 24940 13524
rect 22361 13484 24796 13512
rect 24895 13484 24940 13512
rect 22361 13481 22373 13484
rect 22315 13475 22373 13481
rect 13894 13444 13900 13456
rect 13855 13416 13900 13444
rect 13894 13404 13900 13416
rect 13952 13404 13958 13456
rect 15918 13444 15924 13456
rect 15879 13416 15924 13444
rect 15918 13404 15924 13416
rect 15976 13404 15982 13456
rect 17853 13447 17911 13453
rect 17853 13413 17865 13447
rect 17899 13444 17911 13447
rect 18770 13444 18776 13456
rect 17899 13416 18776 13444
rect 17899 13413 17911 13416
rect 17853 13407 17911 13413
rect 18770 13404 18776 13416
rect 18828 13444 18834 13456
rect 18865 13447 18923 13453
rect 18865 13444 18877 13447
rect 18828 13416 18877 13444
rect 18828 13404 18834 13416
rect 18865 13413 18877 13416
rect 18911 13413 18923 13447
rect 21346 13444 21352 13456
rect 21307 13416 21352 13444
rect 18865 13407 18923 13413
rect 21346 13404 21352 13416
rect 21404 13404 21410 13456
rect 23373 13447 23431 13453
rect 23373 13413 23385 13447
rect 23419 13444 23431 13447
rect 23554 13444 23560 13456
rect 23419 13416 23560 13444
rect 23419 13413 23431 13416
rect 23373 13407 23431 13413
rect 23554 13404 23560 13416
rect 23612 13404 23618 13456
rect 23922 13444 23928 13456
rect 23883 13416 23928 13444
rect 23922 13404 23928 13416
rect 23980 13444 23986 13456
rect 24198 13444 24204 13456
rect 23980 13416 24204 13444
rect 23980 13404 23986 13416
rect 24198 13404 24204 13416
rect 24256 13404 24262 13456
rect 24768 13388 24796 13484
rect 24934 13472 24940 13484
rect 24992 13472 24998 13524
rect 12146 13376 12152 13388
rect 12107 13348 12152 13376
rect 12146 13336 12152 13348
rect 12204 13336 12210 13388
rect 13158 13376 13164 13388
rect 13119 13348 13164 13376
rect 13158 13336 13164 13348
rect 13216 13336 13222 13388
rect 14722 13336 14728 13388
rect 14780 13376 14786 13388
rect 14817 13379 14875 13385
rect 14817 13376 14829 13379
rect 14780 13348 14829 13376
rect 14780 13336 14786 13348
rect 14817 13345 14829 13348
rect 14863 13345 14875 13379
rect 14817 13339 14875 13345
rect 15182 13336 15188 13388
rect 15240 13376 15246 13388
rect 15645 13379 15703 13385
rect 15645 13376 15657 13379
rect 15240 13348 15657 13376
rect 15240 13336 15246 13348
rect 15645 13345 15657 13348
rect 15691 13376 15703 13379
rect 15734 13376 15740 13388
rect 15691 13348 15740 13376
rect 15691 13345 15703 13348
rect 15645 13339 15703 13345
rect 15734 13336 15740 13348
rect 15792 13336 15798 13388
rect 17758 13376 17764 13388
rect 17719 13348 17764 13376
rect 17758 13336 17764 13348
rect 17816 13336 17822 13388
rect 20794 13376 20800 13388
rect 20755 13348 20800 13376
rect 20794 13336 20800 13348
rect 20852 13336 20858 13388
rect 21070 13376 21076 13388
rect 21031 13348 21076 13376
rect 21070 13336 21076 13348
rect 21128 13376 21134 13388
rect 21806 13376 21812 13388
rect 21128 13348 21812 13376
rect 21128 13336 21134 13348
rect 21806 13336 21812 13348
rect 21864 13376 21870 13388
rect 21993 13379 22051 13385
rect 21993 13376 22005 13379
rect 21864 13348 22005 13376
rect 21864 13336 21870 13348
rect 21993 13345 22005 13348
rect 22039 13345 22051 13379
rect 21993 13339 22051 13345
rect 22174 13336 22180 13388
rect 22232 13385 22238 13388
rect 22232 13379 22270 13385
rect 22258 13345 22270 13379
rect 24750 13376 24756 13388
rect 24663 13348 24756 13376
rect 22232 13339 22270 13345
rect 22232 13336 22238 13339
rect 24750 13336 24756 13348
rect 24808 13336 24814 13388
rect 13526 13308 13532 13320
rect 13487 13280 13532 13308
rect 13526 13268 13532 13280
rect 13584 13268 13590 13320
rect 14998 13268 15004 13320
rect 15056 13308 15062 13320
rect 15553 13311 15611 13317
rect 15553 13308 15565 13311
rect 15056 13280 15565 13308
rect 15056 13268 15062 13280
rect 15553 13277 15565 13280
rect 15599 13277 15611 13311
rect 18773 13311 18831 13317
rect 18773 13308 18785 13311
rect 15553 13271 15611 13277
rect 18696 13280 18785 13308
rect 18696 13252 18724 13280
rect 18773 13277 18785 13280
rect 18819 13277 18831 13311
rect 18773 13271 18831 13277
rect 18954 13268 18960 13320
rect 19012 13308 19018 13320
rect 19049 13311 19107 13317
rect 19049 13308 19061 13311
rect 19012 13280 19061 13308
rect 19012 13268 19018 13280
rect 19049 13277 19061 13280
rect 19095 13277 19107 13311
rect 19049 13271 19107 13277
rect 23281 13311 23339 13317
rect 23281 13277 23293 13311
rect 23327 13308 23339 13311
rect 23462 13308 23468 13320
rect 23327 13280 23468 13308
rect 23327 13277 23339 13280
rect 23281 13271 23339 13277
rect 23462 13268 23468 13280
rect 23520 13268 23526 13320
rect 13069 13243 13127 13249
rect 13069 13209 13081 13243
rect 13115 13240 13127 13243
rect 13326 13243 13384 13249
rect 13326 13240 13338 13243
rect 13115 13212 13338 13240
rect 13115 13209 13127 13212
rect 13069 13203 13127 13209
rect 13326 13209 13338 13212
rect 13372 13240 13384 13243
rect 13372 13212 14308 13240
rect 13372 13209 13384 13212
rect 13326 13203 13384 13209
rect 14280 13184 14308 13212
rect 18678 13200 18684 13252
rect 18736 13200 18742 13252
rect 13434 13172 13440 13184
rect 13395 13144 13440 13172
rect 13434 13132 13440 13144
rect 13492 13132 13498 13184
rect 13802 13132 13808 13184
rect 13860 13172 13866 13184
rect 14173 13175 14231 13181
rect 14173 13172 14185 13175
rect 13860 13144 14185 13172
rect 13860 13132 13866 13144
rect 14173 13141 14185 13144
rect 14219 13141 14231 13175
rect 14173 13135 14231 13141
rect 14262 13132 14268 13184
rect 14320 13172 14326 13184
rect 14541 13175 14599 13181
rect 14541 13172 14553 13175
rect 14320 13144 14553 13172
rect 14320 13132 14326 13144
rect 14541 13141 14553 13144
rect 14587 13141 14599 13175
rect 14541 13135 14599 13141
rect 632 13082 26392 13104
rect 632 13030 5176 13082
rect 5228 13030 5240 13082
rect 5292 13030 5304 13082
rect 5356 13030 5368 13082
rect 5420 13030 14510 13082
rect 14562 13030 14574 13082
rect 14626 13030 14638 13082
rect 14690 13030 14702 13082
rect 14754 13030 23843 13082
rect 23895 13030 23907 13082
rect 23959 13030 23971 13082
rect 24023 13030 24035 13082
rect 24087 13030 26392 13082
rect 632 13008 26392 13030
rect 12885 12971 12943 12977
rect 12885 12937 12897 12971
rect 12931 12968 12943 12971
rect 13066 12968 13072 12980
rect 12931 12940 13072 12968
rect 12931 12937 12943 12940
rect 12885 12931 12943 12937
rect 13066 12928 13072 12940
rect 13124 12968 13130 12980
rect 13434 12968 13440 12980
rect 13124 12940 13440 12968
rect 13124 12928 13130 12940
rect 13434 12928 13440 12940
rect 13492 12928 13498 12980
rect 13894 12977 13900 12980
rect 13878 12971 13900 12977
rect 13878 12968 13890 12971
rect 13807 12940 13890 12968
rect 13878 12937 13890 12940
rect 13952 12968 13958 12980
rect 14262 12968 14268 12980
rect 13952 12940 14268 12968
rect 13878 12931 13900 12937
rect 13894 12928 13900 12931
rect 13952 12928 13958 12940
rect 14262 12928 14268 12940
rect 14320 12928 14326 12980
rect 14354 12928 14360 12980
rect 14412 12968 14418 12980
rect 14814 12968 14820 12980
rect 14412 12940 14457 12968
rect 14775 12940 14820 12968
rect 14412 12928 14418 12940
rect 14814 12928 14820 12940
rect 14872 12928 14878 12980
rect 15550 12968 15556 12980
rect 15511 12940 15556 12968
rect 15550 12928 15556 12940
rect 15608 12928 15614 12980
rect 16565 12971 16623 12977
rect 16565 12937 16577 12971
rect 16611 12968 16623 12971
rect 17025 12971 17083 12977
rect 17025 12968 17037 12971
rect 16611 12940 17037 12968
rect 16611 12937 16623 12940
rect 16565 12931 16623 12937
rect 17025 12937 17037 12940
rect 17071 12968 17083 12971
rect 17758 12968 17764 12980
rect 17071 12940 17764 12968
rect 17071 12937 17083 12940
rect 17025 12931 17083 12937
rect 17758 12928 17764 12940
rect 17816 12928 17822 12980
rect 18770 12968 18776 12980
rect 18731 12940 18776 12968
rect 18770 12928 18776 12940
rect 18828 12928 18834 12980
rect 21806 12968 21812 12980
rect 21767 12940 21812 12968
rect 21806 12928 21812 12940
rect 21864 12928 21870 12980
rect 23465 12971 23523 12977
rect 23465 12937 23477 12971
rect 23511 12968 23523 12971
rect 23554 12968 23560 12980
rect 23511 12940 23560 12968
rect 23511 12937 23523 12940
rect 23465 12931 23523 12937
rect 23554 12928 23560 12940
rect 23612 12928 23618 12980
rect 24198 12968 24204 12980
rect 24159 12940 24204 12968
rect 24198 12928 24204 12940
rect 24256 12928 24262 12980
rect 24750 12968 24756 12980
rect 24711 12940 24756 12968
rect 24750 12928 24756 12940
rect 24808 12928 24814 12980
rect 13452 12900 13480 12928
rect 13989 12903 14047 12909
rect 13989 12900 14001 12903
rect 13452 12872 14001 12900
rect 13989 12869 14001 12872
rect 14035 12900 14047 12903
rect 14170 12900 14176 12912
rect 14035 12872 14176 12900
rect 14035 12869 14047 12872
rect 13989 12863 14047 12869
rect 14170 12860 14176 12872
rect 14228 12860 14234 12912
rect 21438 12900 21444 12912
rect 20812 12872 21444 12900
rect 14081 12835 14139 12841
rect 14081 12801 14093 12835
rect 14127 12801 14139 12835
rect 14081 12795 14139 12801
rect 12146 12724 12152 12776
rect 12204 12764 12210 12776
rect 12241 12767 12299 12773
rect 12241 12764 12253 12767
rect 12204 12736 12253 12764
rect 12204 12724 12210 12736
rect 12241 12733 12253 12736
rect 12287 12764 12299 12767
rect 13713 12767 13771 12773
rect 13713 12764 13725 12767
rect 12287 12736 13725 12764
rect 12287 12733 12299 12736
rect 12241 12727 12299 12733
rect 13713 12733 13725 12736
rect 13759 12764 13771 12767
rect 13802 12764 13808 12776
rect 13759 12736 13808 12764
rect 13759 12733 13771 12736
rect 13713 12727 13771 12733
rect 13802 12724 13808 12736
rect 13860 12724 13866 12776
rect 13250 12628 13256 12640
rect 13211 12600 13256 12628
rect 13250 12588 13256 12600
rect 13308 12628 13314 12640
rect 13526 12628 13532 12640
rect 13308 12600 13532 12628
rect 13308 12588 13314 12600
rect 13526 12588 13532 12600
rect 13584 12628 13590 12640
rect 14096 12628 14124 12795
rect 15458 12792 15464 12844
rect 15516 12832 15522 12844
rect 15645 12835 15703 12841
rect 15645 12832 15657 12835
rect 15516 12804 15657 12832
rect 15516 12792 15522 12804
rect 15645 12801 15657 12804
rect 15691 12801 15703 12835
rect 15645 12795 15703 12801
rect 19325 12835 19383 12841
rect 19325 12801 19337 12835
rect 19371 12832 19383 12835
rect 19506 12832 19512 12844
rect 19371 12804 19512 12832
rect 19371 12801 19383 12804
rect 19325 12795 19383 12801
rect 19506 12792 19512 12804
rect 19564 12792 19570 12844
rect 17393 12767 17451 12773
rect 17393 12733 17405 12767
rect 17439 12764 17451 12767
rect 17482 12764 17488 12776
rect 17439 12736 17488 12764
rect 17439 12733 17451 12736
rect 17393 12727 17451 12733
rect 17482 12724 17488 12736
rect 17540 12764 17546 12776
rect 17669 12767 17727 12773
rect 17669 12764 17681 12767
rect 17540 12736 17681 12764
rect 17540 12724 17546 12736
rect 17669 12733 17681 12736
rect 17715 12733 17727 12767
rect 17669 12727 17727 12733
rect 20518 12724 20524 12776
rect 20576 12764 20582 12776
rect 20812 12773 20840 12872
rect 21438 12860 21444 12872
rect 21496 12860 21502 12912
rect 21346 12832 21352 12844
rect 21307 12804 21352 12832
rect 21346 12792 21352 12804
rect 21404 12792 21410 12844
rect 23005 12835 23063 12841
rect 23005 12801 23017 12835
rect 23051 12832 23063 12835
rect 23462 12832 23468 12844
rect 23051 12804 23468 12832
rect 23051 12801 23063 12804
rect 23005 12795 23063 12801
rect 23462 12792 23468 12804
rect 23520 12792 23526 12844
rect 20797 12767 20855 12773
rect 20797 12764 20809 12767
rect 20576 12736 20809 12764
rect 20576 12724 20582 12736
rect 20797 12733 20809 12736
rect 20843 12733 20855 12767
rect 20797 12727 20855 12733
rect 21162 12724 21168 12776
rect 21220 12764 21226 12776
rect 21257 12767 21315 12773
rect 21257 12764 21269 12767
rect 21220 12736 21269 12764
rect 21220 12724 21226 12736
rect 21257 12733 21269 12736
rect 21303 12733 21315 12767
rect 21257 12727 21315 12733
rect 23716 12767 23774 12773
rect 23716 12733 23728 12767
rect 23762 12764 23774 12767
rect 24198 12764 24204 12776
rect 23762 12736 24204 12764
rect 23762 12733 23774 12736
rect 23716 12727 23774 12733
rect 24198 12724 24204 12736
rect 24256 12724 24262 12776
rect 15550 12656 15556 12708
rect 15608 12696 15614 12708
rect 15966 12699 16024 12705
rect 15966 12696 15978 12699
rect 15608 12668 15978 12696
rect 15608 12656 15614 12668
rect 15966 12665 15978 12668
rect 16012 12696 16024 12699
rect 16102 12696 16108 12708
rect 16012 12668 16108 12696
rect 16012 12665 16024 12668
rect 15966 12659 16024 12665
rect 16102 12656 16108 12668
rect 16160 12656 16166 12708
rect 18310 12696 18316 12708
rect 18271 12668 18316 12696
rect 18310 12656 18316 12668
rect 18368 12656 18374 12708
rect 19417 12699 19475 12705
rect 19417 12665 19429 12699
rect 19463 12665 19475 12699
rect 19966 12696 19972 12708
rect 19927 12668 19972 12696
rect 19417 12659 19475 12665
rect 13584 12600 14124 12628
rect 13584 12588 13590 12600
rect 18954 12588 18960 12640
rect 19012 12628 19018 12640
rect 19049 12631 19107 12637
rect 19049 12628 19061 12631
rect 19012 12600 19061 12628
rect 19012 12588 19018 12600
rect 19049 12597 19061 12600
rect 19095 12628 19107 12631
rect 19432 12628 19460 12659
rect 19966 12656 19972 12668
rect 20024 12696 20030 12708
rect 22174 12696 22180 12708
rect 20024 12668 22180 12696
rect 20024 12656 20030 12668
rect 22174 12656 22180 12668
rect 22232 12656 22238 12708
rect 19095 12600 19460 12628
rect 20337 12631 20395 12637
rect 19095 12597 19107 12600
rect 19049 12591 19107 12597
rect 20337 12597 20349 12631
rect 20383 12628 20395 12631
rect 20518 12628 20524 12640
rect 20383 12600 20524 12628
rect 20383 12597 20395 12600
rect 20337 12591 20395 12597
rect 20518 12588 20524 12600
rect 20576 12588 20582 12640
rect 20705 12631 20763 12637
rect 20705 12597 20717 12631
rect 20751 12628 20763 12631
rect 20794 12628 20800 12640
rect 20751 12600 20800 12628
rect 20751 12597 20763 12600
rect 20705 12591 20763 12597
rect 20794 12588 20800 12600
rect 20852 12588 20858 12640
rect 23370 12588 23376 12640
rect 23428 12628 23434 12640
rect 23787 12631 23845 12637
rect 23787 12628 23799 12631
rect 23428 12600 23799 12628
rect 23428 12588 23434 12600
rect 23787 12597 23799 12600
rect 23833 12597 23845 12631
rect 23787 12591 23845 12597
rect 632 12538 26392 12560
rect 632 12486 9843 12538
rect 9895 12486 9907 12538
rect 9959 12486 9971 12538
rect 10023 12486 10035 12538
rect 10087 12486 19176 12538
rect 19228 12486 19240 12538
rect 19292 12486 19304 12538
rect 19356 12486 19368 12538
rect 19420 12486 26392 12538
rect 632 12464 26392 12486
rect 12885 12427 12943 12433
rect 12885 12393 12897 12427
rect 12931 12424 12943 12427
rect 13250 12424 13256 12436
rect 12931 12396 13256 12424
rect 12931 12393 12943 12396
rect 12885 12387 12943 12393
rect 13250 12384 13256 12396
rect 13308 12384 13314 12436
rect 14170 12424 14176 12436
rect 14131 12396 14176 12424
rect 14170 12384 14176 12396
rect 14228 12384 14234 12436
rect 14906 12384 14912 12436
rect 14964 12424 14970 12436
rect 15001 12427 15059 12433
rect 15001 12424 15013 12427
rect 14964 12396 15013 12424
rect 14964 12384 14970 12396
rect 15001 12393 15013 12396
rect 15047 12424 15059 12427
rect 16197 12427 16255 12433
rect 16197 12424 16209 12427
rect 15047 12396 16209 12424
rect 15047 12393 15059 12396
rect 15001 12387 15059 12393
rect 16197 12393 16209 12396
rect 16243 12393 16255 12427
rect 16197 12387 16255 12393
rect 15734 12316 15740 12368
rect 15792 12356 15798 12368
rect 15829 12359 15887 12365
rect 15829 12356 15841 12359
rect 15792 12328 15841 12356
rect 15792 12316 15798 12328
rect 15829 12325 15841 12328
rect 15875 12325 15887 12359
rect 17482 12356 17488 12368
rect 17443 12328 17488 12356
rect 15829 12319 15887 12325
rect 17482 12316 17488 12328
rect 17540 12316 17546 12368
rect 19141 12359 19199 12365
rect 19141 12325 19153 12359
rect 19187 12356 19199 12359
rect 19506 12356 19512 12368
rect 19187 12328 19512 12356
rect 19187 12325 19199 12328
rect 19141 12319 19199 12325
rect 19506 12316 19512 12328
rect 19564 12356 19570 12368
rect 19601 12359 19659 12365
rect 19601 12356 19613 12359
rect 19564 12328 19613 12356
rect 19564 12316 19570 12328
rect 19601 12325 19613 12328
rect 19647 12325 19659 12359
rect 19601 12319 19659 12325
rect 12698 12288 12704 12300
rect 12659 12260 12704 12288
rect 12698 12248 12704 12260
rect 12756 12248 12762 12300
rect 13710 12288 13716 12300
rect 13671 12260 13716 12288
rect 13710 12248 13716 12260
rect 13768 12248 13774 12300
rect 14170 12248 14176 12300
rect 14228 12288 14234 12300
rect 14814 12288 14820 12300
rect 14228 12260 14820 12288
rect 14228 12248 14234 12260
rect 14814 12248 14820 12260
rect 14872 12248 14878 12300
rect 20794 12288 20800 12300
rect 20755 12260 20800 12288
rect 20794 12248 20800 12260
rect 20852 12248 20858 12300
rect 20981 12291 21039 12297
rect 20981 12257 20993 12291
rect 21027 12288 21039 12291
rect 21162 12288 21168 12300
rect 21027 12260 21168 12288
rect 21027 12257 21039 12260
rect 20981 12251 21039 12257
rect 13621 12223 13679 12229
rect 13621 12189 13633 12223
rect 13667 12220 13679 12223
rect 13986 12220 13992 12232
rect 13667 12192 13992 12220
rect 13667 12189 13679 12192
rect 13621 12183 13679 12189
rect 13986 12180 13992 12192
rect 14044 12180 14050 12232
rect 17390 12220 17396 12232
rect 17351 12192 17396 12220
rect 17390 12180 17396 12192
rect 17448 12180 17454 12232
rect 18037 12223 18095 12229
rect 18037 12189 18049 12223
rect 18083 12220 18095 12223
rect 18494 12220 18500 12232
rect 18083 12192 18500 12220
rect 18083 12189 18095 12192
rect 18037 12183 18095 12189
rect 18494 12180 18500 12192
rect 18552 12180 18558 12232
rect 20610 12180 20616 12232
rect 20668 12220 20674 12232
rect 20996 12220 21024 12251
rect 21162 12248 21168 12260
rect 21220 12288 21226 12300
rect 21533 12291 21591 12297
rect 21533 12288 21545 12291
rect 21220 12260 21545 12288
rect 21220 12248 21226 12260
rect 21533 12257 21545 12260
rect 21579 12257 21591 12291
rect 22910 12288 22916 12300
rect 22871 12260 22916 12288
rect 21533 12251 21591 12257
rect 22910 12248 22916 12260
rect 22968 12248 22974 12300
rect 21254 12220 21260 12232
rect 20668 12192 21024 12220
rect 21215 12192 21260 12220
rect 20668 12180 20674 12192
rect 21254 12180 21260 12192
rect 21312 12180 21318 12232
rect 23462 12220 23468 12232
rect 23423 12192 23468 12220
rect 23462 12180 23468 12192
rect 23520 12180 23526 12232
rect 13158 12112 13164 12164
rect 13216 12152 13222 12164
rect 13253 12155 13311 12161
rect 13253 12152 13265 12155
rect 13216 12124 13265 12152
rect 13216 12112 13222 12124
rect 13253 12121 13265 12124
rect 13299 12152 13311 12155
rect 13299 12124 15412 12152
rect 13299 12121 13311 12124
rect 13253 12115 13311 12121
rect 15384 12096 15412 12124
rect 13897 12087 13955 12093
rect 13897 12053 13909 12087
rect 13943 12084 13955 12087
rect 14078 12084 14084 12096
rect 13943 12056 14084 12084
rect 13943 12053 13955 12056
rect 13897 12047 13955 12053
rect 14078 12044 14084 12056
rect 14136 12044 14142 12096
rect 14354 12044 14360 12096
rect 14412 12084 14418 12096
rect 14541 12087 14599 12093
rect 14541 12084 14553 12087
rect 14412 12056 14553 12084
rect 14412 12044 14418 12056
rect 14541 12053 14553 12056
rect 14587 12053 14599 12087
rect 14541 12047 14599 12053
rect 15366 12044 15372 12096
rect 15424 12084 15430 12096
rect 15461 12087 15519 12093
rect 15461 12084 15473 12087
rect 15424 12056 15473 12084
rect 15424 12044 15430 12056
rect 15461 12053 15473 12056
rect 15507 12053 15519 12087
rect 18770 12084 18776 12096
rect 18731 12056 18776 12084
rect 15461 12047 15519 12053
rect 18770 12044 18776 12056
rect 18828 12044 18834 12096
rect 632 11994 26392 12016
rect 632 11942 5176 11994
rect 5228 11942 5240 11994
rect 5292 11942 5304 11994
rect 5356 11942 5368 11994
rect 5420 11942 14510 11994
rect 14562 11942 14574 11994
rect 14626 11942 14638 11994
rect 14690 11942 14702 11994
rect 14754 11942 23843 11994
rect 23895 11942 23907 11994
rect 23959 11942 23971 11994
rect 24023 11942 24035 11994
rect 24087 11942 26392 11994
rect 632 11920 26392 11942
rect 13066 11880 13072 11892
rect 13027 11852 13072 11880
rect 13066 11840 13072 11852
rect 13124 11840 13130 11892
rect 14814 11840 14820 11892
rect 14872 11880 14878 11892
rect 16473 11883 16531 11889
rect 16473 11880 16485 11883
rect 14872 11852 16485 11880
rect 14872 11840 14878 11852
rect 16473 11849 16485 11852
rect 16519 11849 16531 11883
rect 16473 11843 16531 11849
rect 17025 11883 17083 11889
rect 17025 11849 17037 11883
rect 17071 11880 17083 11883
rect 17482 11880 17488 11892
rect 17071 11852 17488 11880
rect 17071 11849 17083 11852
rect 17025 11843 17083 11849
rect 17482 11840 17488 11852
rect 17540 11840 17546 11892
rect 20613 11883 20671 11889
rect 20613 11849 20625 11883
rect 20659 11880 20671 11883
rect 20794 11880 20800 11892
rect 20659 11852 20800 11880
rect 20659 11849 20671 11852
rect 20613 11843 20671 11849
rect 20794 11840 20800 11852
rect 20852 11840 20858 11892
rect 21257 11883 21315 11889
rect 21257 11849 21269 11883
rect 21303 11880 21315 11883
rect 21530 11880 21536 11892
rect 21303 11852 21536 11880
rect 21303 11849 21315 11852
rect 21257 11843 21315 11849
rect 21530 11840 21536 11852
rect 21588 11840 21594 11892
rect 22269 11883 22327 11889
rect 22269 11849 22281 11883
rect 22315 11880 22327 11883
rect 22637 11883 22695 11889
rect 22637 11880 22649 11883
rect 22315 11852 22649 11880
rect 22315 11849 22327 11852
rect 22269 11843 22327 11849
rect 22637 11849 22649 11852
rect 22683 11880 22695 11883
rect 22910 11880 22916 11892
rect 22683 11852 22916 11880
rect 22683 11849 22695 11852
rect 22637 11843 22695 11849
rect 22910 11840 22916 11852
rect 22968 11840 22974 11892
rect 12514 11772 12520 11824
rect 12572 11812 12578 11824
rect 14173 11815 14231 11821
rect 14173 11812 14185 11815
rect 12572 11784 14185 11812
rect 12572 11772 12578 11784
rect 14173 11781 14185 11784
rect 14219 11812 14231 11815
rect 14354 11812 14360 11824
rect 14219 11784 14360 11812
rect 14219 11781 14231 11784
rect 14173 11775 14231 11781
rect 14354 11772 14360 11784
rect 14412 11812 14418 11824
rect 14909 11815 14967 11821
rect 14909 11812 14921 11815
rect 14412 11784 14921 11812
rect 14412 11772 14418 11784
rect 14909 11781 14921 11784
rect 14955 11812 14967 11815
rect 15737 11815 15795 11821
rect 15737 11812 15749 11815
rect 14955 11784 15749 11812
rect 14955 11781 14967 11784
rect 14909 11775 14967 11781
rect 15737 11781 15749 11784
rect 15783 11781 15795 11815
rect 15737 11775 15795 11781
rect 16102 11772 16108 11824
rect 16160 11812 16166 11824
rect 16746 11812 16752 11824
rect 16160 11784 16752 11812
rect 16160 11772 16166 11784
rect 16746 11772 16752 11784
rect 16804 11812 16810 11824
rect 17301 11815 17359 11821
rect 17301 11812 17313 11815
rect 16804 11784 17313 11812
rect 16804 11772 16810 11784
rect 17301 11781 17313 11784
rect 17347 11781 17359 11815
rect 19966 11812 19972 11824
rect 19927 11784 19972 11812
rect 17301 11775 17359 11781
rect 12698 11704 12704 11756
rect 12756 11744 12762 11756
rect 12793 11747 12851 11753
rect 12793 11744 12805 11747
rect 12756 11716 12805 11744
rect 12756 11704 12762 11716
rect 12793 11713 12805 11716
rect 12839 11744 12851 11747
rect 14262 11744 14268 11756
rect 12839 11716 14268 11744
rect 12839 11713 12851 11716
rect 12793 11707 12851 11713
rect 14262 11704 14268 11716
rect 14320 11704 14326 11756
rect 15829 11747 15887 11753
rect 15829 11744 15841 11747
rect 15292 11716 15841 11744
rect 12885 11679 12943 11685
rect 12885 11645 12897 11679
rect 12931 11676 12943 11679
rect 12931 11648 13480 11676
rect 12931 11645 12943 11648
rect 12885 11639 12943 11645
rect 13452 11617 13480 11648
rect 13986 11636 13992 11688
rect 14044 11685 14050 11688
rect 14044 11679 14102 11685
rect 14044 11645 14056 11679
rect 14090 11645 14102 11679
rect 14044 11639 14102 11645
rect 14044 11636 14050 11639
rect 13437 11611 13495 11617
rect 13437 11577 13449 11611
rect 13483 11608 13495 11611
rect 13618 11608 13624 11620
rect 13483 11580 13624 11608
rect 13483 11577 13495 11580
rect 13437 11571 13495 11577
rect 13618 11568 13624 11580
rect 13676 11568 13682 11620
rect 13802 11568 13808 11620
rect 13860 11608 13866 11620
rect 13897 11611 13955 11617
rect 13897 11608 13909 11611
rect 13860 11580 13909 11608
rect 13860 11568 13866 11580
rect 13897 11577 13909 11580
rect 13943 11577 13955 11611
rect 13897 11571 13955 11577
rect 13710 11540 13716 11552
rect 13671 11512 13716 11540
rect 13710 11500 13716 11512
rect 13768 11500 13774 11552
rect 14354 11500 14360 11552
rect 14412 11540 14418 11552
rect 14541 11543 14599 11549
rect 14541 11540 14553 11543
rect 14412 11512 14553 11540
rect 14412 11500 14418 11512
rect 14541 11509 14553 11512
rect 14587 11509 14599 11543
rect 14541 11503 14599 11509
rect 15182 11500 15188 11552
rect 15240 11540 15246 11552
rect 15292 11549 15320 11716
rect 15829 11713 15841 11716
rect 15875 11713 15887 11747
rect 15829 11707 15887 11713
rect 15642 11685 15648 11688
rect 15608 11679 15648 11685
rect 15608 11645 15620 11679
rect 15608 11639 15648 11645
rect 15642 11636 15648 11639
rect 15700 11636 15706 11688
rect 15366 11568 15372 11620
rect 15424 11608 15430 11620
rect 15461 11611 15519 11617
rect 15461 11608 15473 11611
rect 15424 11580 15473 11608
rect 15424 11568 15430 11580
rect 15461 11577 15473 11580
rect 15507 11577 15519 11611
rect 16194 11608 16200 11620
rect 16155 11580 16200 11608
rect 15461 11571 15519 11577
rect 16194 11568 16200 11580
rect 16252 11568 16258 11620
rect 17316 11608 17344 11775
rect 19966 11772 19972 11784
rect 20024 11772 20030 11824
rect 18494 11704 18500 11756
rect 18552 11744 18558 11756
rect 19417 11747 19475 11753
rect 19417 11744 19429 11747
rect 18552 11716 19429 11744
rect 18552 11704 18558 11716
rect 19417 11713 19429 11716
rect 19463 11713 19475 11747
rect 21346 11744 21352 11756
rect 21307 11716 21352 11744
rect 19417 11707 19475 11713
rect 21346 11704 21352 11716
rect 21404 11704 21410 11756
rect 17574 11676 17580 11688
rect 17535 11648 17580 11676
rect 17574 11636 17580 11648
rect 17632 11636 17638 11688
rect 17898 11611 17956 11617
rect 17898 11608 17910 11611
rect 17316 11580 17910 11608
rect 17898 11577 17910 11580
rect 17944 11577 17956 11611
rect 17898 11571 17956 11577
rect 19509 11611 19567 11617
rect 19509 11577 19521 11611
rect 19555 11577 19567 11611
rect 19509 11571 19567 11577
rect 15277 11543 15335 11549
rect 15277 11540 15289 11543
rect 15240 11512 15289 11540
rect 15240 11500 15246 11512
rect 15277 11509 15289 11512
rect 15323 11509 15335 11543
rect 15277 11503 15335 11509
rect 18497 11543 18555 11549
rect 18497 11509 18509 11543
rect 18543 11540 18555 11543
rect 18586 11540 18592 11552
rect 18543 11512 18592 11540
rect 18543 11509 18555 11512
rect 18497 11503 18555 11509
rect 18586 11500 18592 11512
rect 18644 11540 18650 11552
rect 19141 11543 19199 11549
rect 19141 11540 19153 11543
rect 18644 11512 19153 11540
rect 18644 11500 18650 11512
rect 19141 11509 19153 11512
rect 19187 11540 19199 11543
rect 19524 11540 19552 11571
rect 21530 11568 21536 11620
rect 21588 11608 21594 11620
rect 21670 11611 21728 11617
rect 21670 11608 21682 11611
rect 21588 11580 21682 11608
rect 21588 11568 21594 11580
rect 21670 11577 21682 11580
rect 21716 11577 21728 11611
rect 23278 11608 23284 11620
rect 23239 11580 23284 11608
rect 21670 11571 21728 11577
rect 23278 11568 23284 11580
rect 23336 11568 23342 11620
rect 23373 11611 23431 11617
rect 23373 11577 23385 11611
rect 23419 11577 23431 11611
rect 23373 11571 23431 11577
rect 23925 11611 23983 11617
rect 23925 11577 23937 11611
rect 23971 11608 23983 11611
rect 24198 11608 24204 11620
rect 23971 11580 24204 11608
rect 23971 11577 23983 11580
rect 23925 11571 23983 11577
rect 19187 11512 19552 11540
rect 19187 11509 19199 11512
rect 19141 11503 19199 11509
rect 22910 11500 22916 11552
rect 22968 11540 22974 11552
rect 23388 11540 23416 11571
rect 24198 11568 24204 11580
rect 24256 11568 24262 11620
rect 22968 11512 23416 11540
rect 22968 11500 22974 11512
rect 632 11450 26392 11472
rect 632 11398 9843 11450
rect 9895 11398 9907 11450
rect 9959 11398 9971 11450
rect 10023 11398 10035 11450
rect 10087 11398 19176 11450
rect 19228 11398 19240 11450
rect 19292 11398 19304 11450
rect 19356 11398 19368 11450
rect 19420 11398 26392 11450
rect 632 11376 26392 11398
rect 12514 11296 12520 11348
rect 12572 11336 12578 11348
rect 12701 11339 12759 11345
rect 12701 11336 12713 11339
rect 12572 11308 12713 11336
rect 12572 11296 12578 11308
rect 12701 11305 12713 11308
rect 12747 11305 12759 11339
rect 12701 11299 12759 11305
rect 13713 11339 13771 11345
rect 13713 11305 13725 11339
rect 13759 11336 13771 11339
rect 13759 11308 14032 11336
rect 13759 11305 13771 11308
rect 13713 11299 13771 11305
rect 14004 11280 14032 11308
rect 14078 11296 14084 11348
rect 14136 11336 14142 11348
rect 14814 11336 14820 11348
rect 14136 11308 14820 11336
rect 14136 11296 14142 11308
rect 14814 11296 14820 11308
rect 14872 11296 14878 11348
rect 17301 11339 17359 11345
rect 17301 11305 17313 11339
rect 17347 11336 17359 11339
rect 17482 11336 17488 11348
rect 17347 11308 17488 11336
rect 17347 11305 17359 11308
rect 17301 11299 17359 11305
rect 17482 11296 17488 11308
rect 17540 11296 17546 11348
rect 21346 11336 21352 11348
rect 21307 11308 21352 11336
rect 21346 11296 21352 11308
rect 21404 11296 21410 11348
rect 23278 11336 23284 11348
rect 23239 11308 23284 11336
rect 23278 11296 23284 11308
rect 23336 11296 23342 11348
rect 13986 11228 13992 11280
rect 14044 11268 14050 11280
rect 15642 11268 15648 11280
rect 14044 11240 15648 11268
rect 14044 11228 14050 11240
rect 15642 11228 15648 11240
rect 15700 11268 15706 11280
rect 16746 11277 16752 11280
rect 15829 11271 15887 11277
rect 15829 11268 15841 11271
rect 15700 11240 15841 11268
rect 15700 11228 15706 11240
rect 15829 11237 15841 11240
rect 15875 11237 15887 11271
rect 16743 11268 16752 11277
rect 16707 11240 16752 11268
rect 15829 11231 15887 11237
rect 16743 11231 16752 11240
rect 16746 11228 16752 11231
rect 16804 11228 16810 11280
rect 17390 11228 17396 11280
rect 17448 11268 17454 11280
rect 17945 11271 18003 11277
rect 17945 11268 17957 11271
rect 17448 11240 17957 11268
rect 17448 11228 17454 11240
rect 17945 11237 17957 11240
rect 17991 11237 18003 11271
rect 18310 11268 18316 11280
rect 18271 11240 18316 11268
rect 17945 11231 18003 11237
rect 18310 11228 18316 11240
rect 18368 11228 18374 11280
rect 20610 11268 20616 11280
rect 20571 11240 20616 11268
rect 20610 11228 20616 11240
rect 20668 11228 20674 11280
rect 21530 11228 21536 11280
rect 21588 11268 21594 11280
rect 21806 11268 21812 11280
rect 21588 11240 21812 11268
rect 21588 11228 21594 11240
rect 21806 11228 21812 11240
rect 21864 11268 21870 11280
rect 22130 11271 22188 11277
rect 22130 11268 22142 11271
rect 21864 11240 22142 11268
rect 21864 11228 21870 11240
rect 22130 11237 22142 11240
rect 22176 11237 22188 11271
rect 22130 11231 22188 11237
rect 23462 11228 23468 11280
rect 23520 11268 23526 11280
rect 23741 11271 23799 11277
rect 23741 11268 23753 11271
rect 23520 11240 23753 11268
rect 23520 11228 23526 11240
rect 23741 11237 23753 11240
rect 23787 11268 23799 11271
rect 24382 11268 24388 11280
rect 23787 11240 24388 11268
rect 23787 11237 23799 11240
rect 23741 11231 23799 11237
rect 24382 11228 24388 11240
rect 24440 11228 24446 11280
rect 12514 11200 12520 11212
rect 12475 11172 12520 11200
rect 12514 11160 12520 11172
rect 12572 11160 12578 11212
rect 13529 11203 13587 11209
rect 13529 11169 13541 11203
rect 13575 11200 13587 11203
rect 14078 11200 14084 11212
rect 13575 11172 14084 11200
rect 13575 11169 13587 11172
rect 13529 11163 13587 11169
rect 14078 11160 14084 11172
rect 14136 11160 14142 11212
rect 14814 11200 14820 11212
rect 14775 11172 14820 11200
rect 14814 11160 14820 11172
rect 14872 11160 14878 11212
rect 15274 11200 15280 11212
rect 15235 11172 15280 11200
rect 15274 11160 15280 11172
rect 15332 11160 15338 11212
rect 21254 11160 21260 11212
rect 21312 11200 21318 11212
rect 22542 11200 22548 11212
rect 21312 11172 22548 11200
rect 21312 11160 21318 11172
rect 13802 11092 13808 11144
rect 13860 11132 13866 11144
rect 14357 11135 14415 11141
rect 14357 11132 14369 11135
rect 13860 11104 14369 11132
rect 13860 11092 13866 11104
rect 14357 11101 14369 11104
rect 14403 11101 14415 11135
rect 14357 11095 14415 11101
rect 15553 11135 15611 11141
rect 15553 11101 15565 11135
rect 15599 11132 15611 11135
rect 16378 11132 16384 11144
rect 15599 11104 16384 11132
rect 15599 11101 15611 11104
rect 15553 11095 15611 11101
rect 16378 11092 16384 11104
rect 16436 11092 16442 11144
rect 17942 11092 17948 11144
rect 18000 11132 18006 11144
rect 18221 11135 18279 11141
rect 18221 11132 18233 11135
rect 18000 11104 18233 11132
rect 18000 11092 18006 11104
rect 18221 11101 18233 11104
rect 18267 11101 18279 11135
rect 18494 11132 18500 11144
rect 18455 11104 18500 11132
rect 18221 11095 18279 11101
rect 18494 11092 18500 11104
rect 18552 11132 18558 11144
rect 21824 11141 21852 11172
rect 22542 11160 22548 11172
rect 22600 11160 22606 11212
rect 19325 11135 19383 11141
rect 19325 11132 19337 11135
rect 18552 11104 19337 11132
rect 18552 11092 18558 11104
rect 19325 11101 19337 11104
rect 19371 11101 19383 11135
rect 19325 11095 19383 11101
rect 21809 11135 21867 11141
rect 21809 11101 21821 11135
rect 21855 11101 21867 11135
rect 21809 11095 21867 11101
rect 23462 11092 23468 11144
rect 23520 11132 23526 11144
rect 23649 11135 23707 11141
rect 23649 11132 23661 11135
rect 23520 11104 23661 11132
rect 23520 11092 23526 11104
rect 23649 11101 23661 11104
rect 23695 11132 23707 11135
rect 23695 11104 24336 11132
rect 23695 11101 23707 11104
rect 23649 11095 23707 11101
rect 13526 11024 13532 11076
rect 13584 11064 13590 11076
rect 13989 11067 14047 11073
rect 13989 11064 14001 11067
rect 13584 11036 14001 11064
rect 13584 11024 13590 11036
rect 13989 11033 14001 11036
rect 14035 11064 14047 11067
rect 14262 11064 14268 11076
rect 14035 11036 14268 11064
rect 14035 11033 14047 11036
rect 13989 11027 14047 11033
rect 14262 11024 14268 11036
rect 14320 11064 14326 11076
rect 15182 11064 15188 11076
rect 14320 11036 15188 11064
rect 14320 11024 14326 11036
rect 15182 11024 15188 11036
rect 15240 11024 15246 11076
rect 17574 11064 17580 11076
rect 17408 11036 17580 11064
rect 16562 10956 16568 11008
rect 16620 10996 16626 11008
rect 17408 10996 17436 11036
rect 17574 11024 17580 11036
rect 17632 11024 17638 11076
rect 22729 11067 22787 11073
rect 22729 11033 22741 11067
rect 22775 11064 22787 11067
rect 24198 11064 24204 11076
rect 22775 11036 22956 11064
rect 24159 11036 24204 11064
rect 22775 11033 22787 11036
rect 22729 11027 22787 11033
rect 16620 10968 17436 10996
rect 22928 10996 22956 11036
rect 24198 11024 24204 11036
rect 24256 11024 24262 11076
rect 23002 10996 23008 11008
rect 22928 10968 23008 10996
rect 16620 10956 16626 10968
rect 23002 10956 23008 10968
rect 23060 10956 23066 11008
rect 24308 10996 24336 11104
rect 24750 10996 24756 11008
rect 24308 10968 24756 10996
rect 24750 10956 24756 10968
rect 24808 10956 24814 11008
rect 632 10906 26392 10928
rect 632 10854 5176 10906
rect 5228 10854 5240 10906
rect 5292 10854 5304 10906
rect 5356 10854 5368 10906
rect 5420 10854 14510 10906
rect 14562 10854 14574 10906
rect 14626 10854 14638 10906
rect 14690 10854 14702 10906
rect 14754 10854 23843 10906
rect 23895 10854 23907 10906
rect 23959 10854 23971 10906
rect 24023 10854 24035 10906
rect 24087 10854 26392 10906
rect 632 10832 26392 10854
rect 12514 10792 12520 10804
rect 12475 10764 12520 10792
rect 12514 10752 12520 10764
rect 12572 10792 12578 10804
rect 13342 10792 13348 10804
rect 12572 10764 13348 10792
rect 12572 10752 12578 10764
rect 13342 10752 13348 10764
rect 13400 10752 13406 10804
rect 14078 10792 14084 10804
rect 14039 10764 14084 10792
rect 14078 10752 14084 10764
rect 14136 10752 14142 10804
rect 14817 10795 14875 10801
rect 14817 10761 14829 10795
rect 14863 10792 14875 10795
rect 14998 10792 15004 10804
rect 14863 10764 15004 10792
rect 14863 10761 14875 10764
rect 14817 10755 14875 10761
rect 14998 10752 15004 10764
rect 15056 10752 15062 10804
rect 15734 10792 15740 10804
rect 15695 10764 15740 10792
rect 15734 10752 15740 10764
rect 15792 10752 15798 10804
rect 16378 10752 16384 10804
rect 16436 10792 16442 10804
rect 17209 10795 17267 10801
rect 17209 10792 17221 10795
rect 16436 10764 17221 10792
rect 16436 10752 16442 10764
rect 17209 10761 17221 10764
rect 17255 10761 17267 10795
rect 17209 10755 17267 10761
rect 18221 10795 18279 10801
rect 18221 10761 18233 10795
rect 18267 10792 18279 10795
rect 18310 10792 18316 10804
rect 18267 10764 18316 10792
rect 18267 10761 18279 10764
rect 18221 10755 18279 10761
rect 18310 10752 18316 10764
rect 18368 10752 18374 10804
rect 18586 10792 18592 10804
rect 18547 10764 18592 10792
rect 18586 10752 18592 10764
rect 18644 10752 18650 10804
rect 18954 10792 18960 10804
rect 18915 10764 18960 10792
rect 18954 10752 18960 10764
rect 19012 10752 19018 10804
rect 22542 10792 22548 10804
rect 22503 10764 22548 10792
rect 22542 10752 22548 10764
rect 22600 10752 22606 10804
rect 24382 10792 24388 10804
rect 24343 10764 24388 10792
rect 24382 10752 24388 10764
rect 24440 10752 24446 10804
rect 24750 10792 24756 10804
rect 24711 10764 24756 10792
rect 24750 10752 24756 10764
rect 24808 10752 24814 10804
rect 25118 10792 25124 10804
rect 25079 10764 25124 10792
rect 25118 10752 25124 10764
rect 25176 10752 25182 10804
rect 16746 10684 16752 10736
rect 16804 10724 16810 10736
rect 16841 10727 16899 10733
rect 16841 10724 16853 10727
rect 16804 10696 16853 10724
rect 16804 10684 16810 10696
rect 16841 10693 16853 10696
rect 16887 10693 16899 10727
rect 16841 10687 16899 10693
rect 16562 10656 16568 10668
rect 16523 10628 16568 10656
rect 16562 10616 16568 10628
rect 16620 10616 16626 10668
rect 19690 10656 19696 10668
rect 19651 10628 19696 10656
rect 19690 10616 19696 10628
rect 19748 10616 19754 10668
rect 20153 10659 20211 10665
rect 20153 10625 20165 10659
rect 20199 10656 20211 10659
rect 20794 10656 20800 10668
rect 20199 10628 20800 10656
rect 20199 10625 20211 10628
rect 20153 10619 20211 10625
rect 13529 10591 13587 10597
rect 13529 10557 13541 10591
rect 13575 10557 13587 10591
rect 13529 10551 13587 10557
rect 12977 10455 13035 10461
rect 12977 10421 12989 10455
rect 13023 10452 13035 10455
rect 13544 10452 13572 10551
rect 13894 10548 13900 10600
rect 13952 10588 13958 10600
rect 14633 10591 14691 10597
rect 14633 10588 14645 10591
rect 13952 10560 14645 10588
rect 13952 10548 13958 10560
rect 14633 10557 14645 10560
rect 14679 10588 14691 10591
rect 15093 10591 15151 10597
rect 15093 10588 15105 10591
rect 14679 10560 15105 10588
rect 14679 10557 14691 10560
rect 14633 10551 14691 10557
rect 15093 10557 15105 10560
rect 15139 10588 15151 10591
rect 15182 10588 15188 10600
rect 15139 10560 15188 10588
rect 15139 10557 15151 10560
rect 15093 10551 15151 10557
rect 15182 10548 15188 10560
rect 15240 10548 15246 10600
rect 15734 10548 15740 10600
rect 15792 10588 15798 10600
rect 15829 10591 15887 10597
rect 15829 10588 15841 10591
rect 15792 10560 15841 10588
rect 15792 10548 15798 10560
rect 15829 10557 15841 10560
rect 15875 10557 15887 10591
rect 16286 10588 16292 10600
rect 16247 10560 16292 10588
rect 15829 10551 15887 10557
rect 16286 10548 16292 10560
rect 16344 10548 16350 10600
rect 18586 10548 18592 10600
rect 18644 10588 18650 10600
rect 18773 10591 18831 10597
rect 18773 10588 18785 10591
rect 18644 10560 18785 10588
rect 18644 10548 18650 10560
rect 18773 10557 18785 10560
rect 18819 10557 18831 10591
rect 18773 10551 18831 10557
rect 19708 10520 19736 10616
rect 20536 10597 20564 10628
rect 20794 10616 20800 10628
rect 20852 10616 20858 10668
rect 23465 10659 23523 10665
rect 23465 10625 23477 10659
rect 23511 10656 23523 10659
rect 24198 10656 24204 10668
rect 23511 10628 24204 10656
rect 23511 10625 23523 10628
rect 23465 10619 23523 10625
rect 24198 10616 24204 10628
rect 24256 10616 24262 10668
rect 20521 10591 20579 10597
rect 20521 10557 20533 10591
rect 20567 10557 20579 10591
rect 20521 10551 20579 10557
rect 20705 10591 20763 10597
rect 20705 10557 20717 10591
rect 20751 10557 20763 10591
rect 24934 10588 24940 10600
rect 24895 10560 24940 10588
rect 20705 10551 20763 10557
rect 20720 10520 20748 10551
rect 24934 10548 24940 10560
rect 24992 10588 24998 10600
rect 25489 10591 25547 10597
rect 25489 10588 25501 10591
rect 24992 10560 25501 10588
rect 24992 10548 24998 10560
rect 25489 10557 25501 10560
rect 25535 10557 25547 10591
rect 25489 10551 25547 10557
rect 20886 10520 20892 10532
rect 19708 10492 20892 10520
rect 20886 10480 20892 10492
rect 20944 10480 20950 10532
rect 20981 10523 21039 10529
rect 20981 10489 20993 10523
rect 21027 10520 21039 10523
rect 21530 10520 21536 10532
rect 21027 10492 21536 10520
rect 21027 10489 21039 10492
rect 20981 10483 21039 10489
rect 21530 10480 21536 10492
rect 21588 10480 21594 10532
rect 23557 10523 23615 10529
rect 23557 10489 23569 10523
rect 23603 10489 23615 10523
rect 23557 10483 23615 10489
rect 13618 10452 13624 10464
rect 13023 10424 13624 10452
rect 13023 10421 13035 10424
rect 12977 10415 13035 10421
rect 13618 10412 13624 10424
rect 13676 10412 13682 10464
rect 14541 10455 14599 10461
rect 14541 10421 14553 10455
rect 14587 10452 14599 10455
rect 14630 10452 14636 10464
rect 14587 10424 14636 10452
rect 14587 10421 14599 10424
rect 14541 10415 14599 10421
rect 14630 10412 14636 10424
rect 14688 10412 14694 10464
rect 17853 10455 17911 10461
rect 17853 10421 17865 10455
rect 17899 10452 17911 10455
rect 17942 10452 17948 10464
rect 17899 10424 17948 10452
rect 17899 10421 17911 10424
rect 17853 10415 17911 10421
rect 17942 10412 17948 10424
rect 18000 10412 18006 10464
rect 21806 10452 21812 10464
rect 21767 10424 21812 10452
rect 21806 10412 21812 10424
rect 21864 10412 21870 10464
rect 22082 10452 22088 10464
rect 22043 10424 22088 10452
rect 22082 10412 22088 10424
rect 22140 10412 22146 10464
rect 23002 10452 23008 10464
rect 22915 10424 23008 10452
rect 23002 10412 23008 10424
rect 23060 10452 23066 10464
rect 23278 10452 23284 10464
rect 23060 10424 23284 10452
rect 23060 10412 23066 10424
rect 23278 10412 23284 10424
rect 23336 10452 23342 10464
rect 23572 10452 23600 10483
rect 23922 10480 23928 10532
rect 23980 10520 23986 10532
rect 24109 10523 24167 10529
rect 24109 10520 24121 10523
rect 23980 10492 24121 10520
rect 23980 10480 23986 10492
rect 24109 10489 24121 10492
rect 24155 10489 24167 10523
rect 24109 10483 24167 10489
rect 23336 10424 23600 10452
rect 23336 10412 23342 10424
rect 632 10362 26392 10384
rect 632 10310 9843 10362
rect 9895 10310 9907 10362
rect 9959 10310 9971 10362
rect 10023 10310 10035 10362
rect 10087 10310 19176 10362
rect 19228 10310 19240 10362
rect 19292 10310 19304 10362
rect 19356 10310 19368 10362
rect 19420 10310 26392 10362
rect 632 10288 26392 10310
rect 14078 10208 14084 10260
rect 14136 10248 14142 10260
rect 14541 10251 14599 10257
rect 14541 10248 14553 10251
rect 14136 10220 14553 10248
rect 14136 10208 14142 10220
rect 14541 10217 14553 10220
rect 14587 10217 14599 10251
rect 16286 10248 16292 10260
rect 16247 10220 16292 10248
rect 14541 10211 14599 10217
rect 13894 10180 13900 10192
rect 13855 10152 13900 10180
rect 13894 10140 13900 10152
rect 13952 10140 13958 10192
rect 13526 10112 13532 10124
rect 13487 10084 13532 10112
rect 13526 10072 13532 10084
rect 13584 10072 13590 10124
rect 14556 10044 14584 10211
rect 16286 10208 16292 10220
rect 16344 10208 16350 10260
rect 20702 10248 20708 10260
rect 20663 10220 20708 10248
rect 20702 10208 20708 10220
rect 20760 10208 20766 10260
rect 22683 10251 22741 10257
rect 22683 10217 22695 10251
rect 22729 10248 22741 10251
rect 22910 10248 22916 10260
rect 22729 10220 22916 10248
rect 22729 10217 22741 10220
rect 22683 10211 22741 10217
rect 22910 10208 22916 10220
rect 22968 10208 22974 10260
rect 24198 10208 24204 10260
rect 24256 10248 24262 10260
rect 24569 10251 24627 10257
rect 24569 10248 24581 10251
rect 24256 10220 24581 10248
rect 24256 10208 24262 10220
rect 24569 10217 24581 10220
rect 24615 10217 24627 10251
rect 24569 10211 24627 10217
rect 23646 10140 23652 10192
rect 23704 10180 23710 10192
rect 23741 10183 23799 10189
rect 23741 10180 23753 10183
rect 23704 10152 23753 10180
rect 23704 10140 23710 10152
rect 23741 10149 23753 10152
rect 23787 10149 23799 10183
rect 23741 10143 23799 10149
rect 14814 10112 14820 10124
rect 14775 10084 14820 10112
rect 14814 10072 14820 10084
rect 14872 10072 14878 10124
rect 18862 10112 18868 10124
rect 18823 10084 18868 10112
rect 18862 10072 18868 10084
rect 18920 10072 18926 10124
rect 20518 10112 20524 10124
rect 20479 10084 20524 10112
rect 20518 10072 20524 10084
rect 20576 10072 20582 10124
rect 20886 10112 20892 10124
rect 20847 10084 20892 10112
rect 20886 10072 20892 10084
rect 20944 10072 20950 10124
rect 22634 10121 22640 10124
rect 22612 10115 22640 10121
rect 22612 10081 22624 10115
rect 22612 10075 22640 10081
rect 22634 10072 22640 10075
rect 22692 10072 22698 10124
rect 14964 10047 15022 10053
rect 14964 10044 14976 10047
rect 14556 10016 14976 10044
rect 14964 10013 14976 10016
rect 15010 10013 15022 10047
rect 15182 10044 15188 10056
rect 15143 10016 15188 10044
rect 14964 10007 15022 10013
rect 15182 10004 15188 10016
rect 15240 10004 15246 10056
rect 22910 10004 22916 10056
rect 22968 10044 22974 10056
rect 23649 10047 23707 10053
rect 23649 10044 23661 10047
rect 22968 10016 23661 10044
rect 22968 10004 22974 10016
rect 23649 10013 23661 10016
rect 23695 10013 23707 10047
rect 23922 10044 23928 10056
rect 23835 10016 23928 10044
rect 23649 10007 23707 10013
rect 23922 10004 23928 10016
rect 23980 10004 23986 10056
rect 14265 9979 14323 9985
rect 14265 9945 14277 9979
rect 14311 9976 14323 9979
rect 15274 9976 15280 9988
rect 14311 9948 15280 9976
rect 14311 9945 14323 9948
rect 14265 9939 14323 9945
rect 15274 9936 15280 9948
rect 15332 9976 15338 9988
rect 16286 9976 16292 9988
rect 15332 9948 16292 9976
rect 15332 9936 15338 9948
rect 16286 9936 16292 9948
rect 16344 9936 16350 9988
rect 22634 9936 22640 9988
rect 22692 9976 22698 9988
rect 23940 9976 23968 10004
rect 22692 9948 23968 9976
rect 22692 9936 22698 9948
rect 13342 9868 13348 9920
rect 13400 9908 13406 9920
rect 15093 9911 15151 9917
rect 15093 9908 15105 9911
rect 13400 9880 15105 9908
rect 13400 9868 13406 9880
rect 15093 9877 15105 9880
rect 15139 9908 15151 9911
rect 15550 9908 15556 9920
rect 15139 9880 15556 9908
rect 15139 9877 15151 9880
rect 15093 9871 15151 9877
rect 15550 9868 15556 9880
rect 15608 9908 15614 9920
rect 15826 9908 15832 9920
rect 15608 9880 15832 9908
rect 15608 9868 15614 9880
rect 15826 9868 15832 9880
rect 15884 9868 15890 9920
rect 18954 9908 18960 9920
rect 18915 9880 18960 9908
rect 18954 9868 18960 9880
rect 19012 9868 19018 9920
rect 23278 9908 23284 9920
rect 23239 9880 23284 9908
rect 23278 9868 23284 9880
rect 23336 9868 23342 9920
rect 632 9818 26392 9840
rect 632 9766 5176 9818
rect 5228 9766 5240 9818
rect 5292 9766 5304 9818
rect 5356 9766 5368 9818
rect 5420 9766 14510 9818
rect 14562 9766 14574 9818
rect 14626 9766 14638 9818
rect 14690 9766 14702 9818
rect 14754 9766 23843 9818
rect 23895 9766 23907 9818
rect 23959 9766 23971 9818
rect 24023 9766 24035 9818
rect 24087 9766 26392 9818
rect 632 9744 26392 9766
rect 12606 9704 12612 9716
rect 12567 9676 12612 9704
rect 12606 9664 12612 9676
rect 12664 9664 12670 9716
rect 15182 9664 15188 9716
rect 15240 9704 15246 9716
rect 15240 9676 15688 9704
rect 15240 9664 15246 9676
rect 15550 9636 15556 9648
rect 15511 9608 15556 9636
rect 15550 9596 15556 9608
rect 15608 9596 15614 9648
rect 14078 9568 14084 9580
rect 14039 9540 14084 9568
rect 14078 9528 14084 9540
rect 14136 9568 14142 9580
rect 15660 9577 15688 9676
rect 20886 9664 20892 9716
rect 20944 9704 20950 9716
rect 21257 9707 21315 9713
rect 21257 9704 21269 9707
rect 20944 9676 21269 9704
rect 20944 9664 20950 9676
rect 21257 9673 21269 9676
rect 21303 9673 21315 9707
rect 21257 9667 21315 9673
rect 22082 9664 22088 9716
rect 22140 9704 22146 9716
rect 22910 9704 22916 9716
rect 22140 9676 22916 9704
rect 22140 9664 22146 9676
rect 22910 9664 22916 9676
rect 22968 9664 22974 9716
rect 24198 9664 24204 9716
rect 24256 9704 24262 9716
rect 25762 9704 25768 9716
rect 24256 9676 25768 9704
rect 24256 9664 24262 9676
rect 25762 9664 25768 9676
rect 25820 9664 25826 9716
rect 15826 9596 15832 9648
rect 15884 9636 15890 9648
rect 16289 9639 16347 9645
rect 16289 9636 16301 9639
rect 15884 9608 16301 9636
rect 15884 9596 15890 9608
rect 16289 9605 16301 9608
rect 16335 9605 16347 9639
rect 16289 9599 16347 9605
rect 18405 9639 18463 9645
rect 18405 9605 18417 9639
rect 18451 9636 18463 9639
rect 18773 9639 18831 9645
rect 18773 9636 18785 9639
rect 18451 9608 18785 9636
rect 18451 9605 18463 9608
rect 18405 9599 18463 9605
rect 18773 9605 18785 9608
rect 18819 9636 18831 9639
rect 18862 9636 18868 9648
rect 18819 9608 18868 9636
rect 18819 9605 18831 9608
rect 18773 9599 18831 9605
rect 18862 9596 18868 9608
rect 18920 9596 18926 9648
rect 24382 9596 24388 9648
rect 24440 9636 24446 9648
rect 24937 9639 24995 9645
rect 24937 9636 24949 9639
rect 24440 9608 24949 9636
rect 24440 9596 24446 9608
rect 24937 9605 24949 9608
rect 24983 9605 24995 9639
rect 24937 9599 24995 9605
rect 15424 9571 15482 9577
rect 15424 9568 15436 9571
rect 14136 9540 15436 9568
rect 14136 9528 14142 9540
rect 15424 9537 15436 9540
rect 15470 9568 15482 9571
rect 15645 9571 15703 9577
rect 15470 9537 15504 9568
rect 15424 9531 15504 9537
rect 15645 9537 15657 9571
rect 15691 9537 15703 9571
rect 15645 9531 15703 9537
rect 12241 9503 12299 9509
rect 12241 9469 12253 9503
rect 12287 9500 12299 9503
rect 12517 9503 12575 9509
rect 12517 9500 12529 9503
rect 12287 9472 12529 9500
rect 12287 9469 12299 9472
rect 12241 9463 12299 9469
rect 12517 9469 12529 9472
rect 12563 9469 12575 9503
rect 13710 9500 13716 9512
rect 13671 9472 13716 9500
rect 12517 9463 12575 9469
rect 12330 9432 12336 9444
rect 12291 9404 12336 9432
rect 12330 9392 12336 9404
rect 12388 9392 12394 9444
rect 12532 9432 12560 9463
rect 13710 9460 13716 9472
rect 13768 9460 13774 9512
rect 14262 9500 14268 9512
rect 14223 9472 14268 9500
rect 14262 9460 14268 9472
rect 14320 9460 14326 9512
rect 14814 9500 14820 9512
rect 14727 9472 14820 9500
rect 14814 9460 14820 9472
rect 14872 9500 14878 9512
rect 15476 9500 15504 9531
rect 20518 9528 20524 9580
rect 20576 9568 20582 9580
rect 20889 9571 20947 9577
rect 20889 9568 20901 9571
rect 20576 9540 20901 9568
rect 20576 9528 20582 9540
rect 20889 9537 20901 9540
rect 20935 9537 20947 9571
rect 20889 9531 20947 9537
rect 23738 9528 23744 9580
rect 23796 9568 23802 9580
rect 23925 9571 23983 9577
rect 23925 9568 23937 9571
rect 23796 9540 23937 9568
rect 23796 9528 23802 9540
rect 23925 9537 23937 9540
rect 23971 9568 23983 9571
rect 24201 9571 24259 9577
rect 24201 9568 24213 9571
rect 23971 9540 24213 9568
rect 23971 9537 23983 9540
rect 23925 9531 23983 9537
rect 24201 9537 24213 9540
rect 24247 9537 24259 9571
rect 24201 9531 24259 9537
rect 16657 9503 16715 9509
rect 16657 9500 16669 9503
rect 14872 9472 15412 9500
rect 15476 9472 16669 9500
rect 14872 9460 14878 9472
rect 13621 9435 13679 9441
rect 13621 9432 13633 9435
rect 12532 9404 13633 9432
rect 13621 9401 13633 9404
rect 13667 9432 13679 9435
rect 14280 9432 14308 9460
rect 15384 9444 15412 9472
rect 16657 9469 16669 9472
rect 16703 9469 16715 9503
rect 16657 9463 16715 9469
rect 22082 9460 22088 9512
rect 22140 9509 22146 9512
rect 22140 9503 22178 9509
rect 22166 9500 22178 9503
rect 22545 9503 22603 9509
rect 22545 9500 22557 9503
rect 22166 9472 22557 9500
rect 22166 9469 22178 9472
rect 22140 9463 22178 9469
rect 22545 9469 22557 9472
rect 22591 9469 22603 9503
rect 23278 9500 23284 9512
rect 23239 9472 23284 9500
rect 22545 9463 22603 9469
rect 22140 9460 22146 9463
rect 23278 9460 23284 9472
rect 23336 9460 23342 9512
rect 24753 9503 24811 9509
rect 24753 9469 24765 9503
rect 24799 9469 24811 9503
rect 24753 9463 24811 9469
rect 13667 9404 14308 9432
rect 15277 9435 15335 9441
rect 13667 9401 13679 9404
rect 13621 9395 13679 9401
rect 15277 9401 15289 9435
rect 15323 9401 15335 9435
rect 15277 9395 15335 9401
rect 13253 9367 13311 9373
rect 13253 9333 13265 9367
rect 13299 9364 13311 9367
rect 13526 9364 13532 9376
rect 13299 9336 13532 9364
rect 13299 9333 13311 9336
rect 13253 9327 13311 9333
rect 13526 9324 13532 9336
rect 13584 9324 13590 9376
rect 15090 9364 15096 9376
rect 15051 9336 15096 9364
rect 15090 9324 15096 9336
rect 15148 9364 15154 9376
rect 15292 9364 15320 9395
rect 15366 9392 15372 9444
rect 15424 9392 15430 9444
rect 18037 9435 18095 9441
rect 18037 9401 18049 9435
rect 18083 9432 18095 9435
rect 18770 9432 18776 9444
rect 18083 9404 18776 9432
rect 18083 9401 18095 9404
rect 18037 9395 18095 9401
rect 18770 9392 18776 9404
rect 18828 9432 18834 9444
rect 18957 9435 19015 9441
rect 18957 9432 18969 9435
rect 18828 9404 18969 9432
rect 18828 9392 18834 9404
rect 18957 9401 18969 9404
rect 19003 9401 19015 9435
rect 18957 9395 19015 9401
rect 19049 9435 19107 9441
rect 19049 9401 19061 9435
rect 19095 9401 19107 9435
rect 19049 9395 19107 9401
rect 19601 9435 19659 9441
rect 19601 9401 19613 9435
rect 19647 9432 19659 9435
rect 19690 9432 19696 9444
rect 19647 9404 19696 9432
rect 19647 9401 19659 9404
rect 19601 9395 19659 9401
rect 15918 9364 15924 9376
rect 15148 9336 15320 9364
rect 15879 9336 15924 9364
rect 15148 9324 15154 9336
rect 15918 9324 15924 9336
rect 15976 9324 15982 9376
rect 18862 9324 18868 9376
rect 18920 9364 18926 9376
rect 19064 9364 19092 9395
rect 19690 9392 19696 9404
rect 19748 9392 19754 9444
rect 22223 9435 22281 9441
rect 22223 9401 22235 9435
rect 22269 9432 22281 9435
rect 24768 9432 24796 9463
rect 25305 9435 25363 9441
rect 25305 9432 25317 9435
rect 22269 9404 25317 9432
rect 22269 9401 22281 9404
rect 22223 9395 22281 9401
rect 25305 9401 25317 9404
rect 25351 9401 25363 9435
rect 25305 9395 25363 9401
rect 20426 9364 20432 9376
rect 18920 9336 19092 9364
rect 20387 9336 20432 9364
rect 18920 9324 18926 9336
rect 20426 9324 20432 9336
rect 20484 9324 20490 9376
rect 632 9274 26392 9296
rect 632 9222 9843 9274
rect 9895 9222 9907 9274
rect 9959 9222 9971 9274
rect 10023 9222 10035 9274
rect 10087 9222 19176 9274
rect 19228 9222 19240 9274
rect 19292 9222 19304 9274
rect 19356 9222 19368 9274
rect 19420 9222 26392 9274
rect 632 9200 26392 9222
rect 13805 9163 13863 9169
rect 13805 9129 13817 9163
rect 13851 9160 13863 9163
rect 14170 9160 14176 9172
rect 13851 9132 14176 9160
rect 13851 9129 13863 9132
rect 13805 9123 13863 9129
rect 14170 9120 14176 9132
rect 14228 9120 14234 9172
rect 14633 9163 14691 9169
rect 14633 9129 14645 9163
rect 14679 9160 14691 9163
rect 15182 9160 15188 9172
rect 14679 9132 15188 9160
rect 14679 9129 14691 9132
rect 14633 9123 14691 9129
rect 15182 9120 15188 9132
rect 15240 9160 15246 9172
rect 16013 9163 16071 9169
rect 16013 9160 16025 9163
rect 15240 9132 16025 9160
rect 15240 9120 15246 9132
rect 16013 9129 16025 9132
rect 16059 9129 16071 9163
rect 16013 9123 16071 9129
rect 19417 9163 19475 9169
rect 19417 9129 19429 9163
rect 19463 9160 19475 9163
rect 19506 9160 19512 9172
rect 19463 9132 19512 9160
rect 19463 9129 19475 9132
rect 19417 9123 19475 9129
rect 19506 9120 19512 9132
rect 19564 9160 19570 9172
rect 20426 9160 20432 9172
rect 19564 9132 20432 9160
rect 19564 9120 19570 9132
rect 20426 9120 20432 9132
rect 20484 9120 20490 9172
rect 21530 9120 21536 9172
rect 21588 9160 21594 9172
rect 21901 9163 21959 9169
rect 21901 9160 21913 9163
rect 21588 9132 21913 9160
rect 21588 9120 21594 9132
rect 21901 9129 21913 9132
rect 21947 9129 21959 9163
rect 22634 9160 22640 9172
rect 22595 9132 22640 9160
rect 21901 9123 21959 9129
rect 22634 9120 22640 9132
rect 22692 9120 22698 9172
rect 24658 9160 24664 9172
rect 24619 9132 24664 9160
rect 24658 9120 24664 9132
rect 24716 9120 24722 9172
rect 12330 9052 12336 9104
rect 12388 9092 12394 9104
rect 12425 9095 12483 9101
rect 12425 9092 12437 9095
rect 12388 9064 12437 9092
rect 12388 9052 12394 9064
rect 12425 9061 12437 9064
rect 12471 9092 12483 9095
rect 14354 9092 14360 9104
rect 12471 9064 14360 9092
rect 12471 9061 12483 9064
rect 12425 9055 12483 9061
rect 14354 9052 14360 9064
rect 14412 9052 14418 9104
rect 16746 9052 16752 9104
rect 16804 9092 16810 9104
rect 16886 9095 16944 9101
rect 16886 9092 16898 9095
rect 16804 9064 16898 9092
rect 16804 9052 16810 9064
rect 16886 9061 16898 9064
rect 16932 9061 16944 9095
rect 16886 9055 16944 9061
rect 17666 9052 17672 9104
rect 17724 9092 17730 9104
rect 18497 9095 18555 9101
rect 18497 9092 18509 9095
rect 17724 9064 18509 9092
rect 17724 9052 17730 9064
rect 18497 9061 18509 9064
rect 18543 9061 18555 9095
rect 18497 9055 18555 9061
rect 21067 9095 21125 9101
rect 21067 9061 21079 9095
rect 21113 9092 21125 9095
rect 21254 9092 21260 9104
rect 21113 9064 21260 9092
rect 21113 9061 21125 9064
rect 21067 9055 21125 9061
rect 21254 9052 21260 9064
rect 21312 9092 21318 9104
rect 21806 9092 21812 9104
rect 21312 9064 21812 9092
rect 21312 9052 21318 9064
rect 21806 9052 21812 9064
rect 21864 9052 21870 9104
rect 23094 9092 23100 9104
rect 23055 9064 23100 9092
rect 23094 9052 23100 9064
rect 23152 9052 23158 9104
rect 13161 9027 13219 9033
rect 13161 8993 13173 9027
rect 13207 9024 13219 9027
rect 13250 9024 13256 9036
rect 13207 8996 13256 9024
rect 13207 8993 13219 8996
rect 13161 8987 13219 8993
rect 13250 8984 13256 8996
rect 13308 9024 13314 9036
rect 13710 9024 13716 9036
rect 13308 8996 13716 9024
rect 13308 8984 13314 8996
rect 13710 8984 13716 8996
rect 13768 9024 13774 9036
rect 14173 9027 14231 9033
rect 14173 9024 14185 9027
rect 13768 8996 14185 9024
rect 13768 8984 13774 8996
rect 14173 8993 14185 8996
rect 14219 8993 14231 9027
rect 14173 8987 14231 8993
rect 14906 8984 14912 9036
rect 14964 9024 14970 9036
rect 15001 9027 15059 9033
rect 15001 9024 15013 9027
rect 14964 8996 15013 9024
rect 14964 8984 14970 8996
rect 15001 8993 15013 8996
rect 15047 8993 15059 9027
rect 15001 8987 15059 8993
rect 15458 8984 15464 9036
rect 15516 9024 15522 9036
rect 15553 9027 15611 9033
rect 15553 9024 15565 9027
rect 15516 8996 15565 9024
rect 15516 8984 15522 8996
rect 15553 8993 15565 8996
rect 15599 9024 15611 9027
rect 15918 9024 15924 9036
rect 15599 8996 15924 9024
rect 15599 8993 15611 8996
rect 15553 8987 15611 8993
rect 15918 8984 15924 8996
rect 15976 9024 15982 9036
rect 16378 9024 16384 9036
rect 15976 8996 16384 9024
rect 15976 8984 15982 8996
rect 16378 8984 16384 8996
rect 16436 8984 16442 9036
rect 20702 9024 20708 9036
rect 20663 8996 20708 9024
rect 20702 8984 20708 8996
rect 20760 8984 20766 9036
rect 24382 8984 24388 9036
rect 24440 9024 24446 9036
rect 24477 9027 24535 9033
rect 24477 9024 24489 9027
rect 24440 8996 24489 9024
rect 24440 8984 24446 8996
rect 24477 8993 24489 8996
rect 24523 8993 24535 9027
rect 24477 8987 24535 8993
rect 13526 8956 13532 8968
rect 13487 8928 13532 8956
rect 13526 8916 13532 8928
rect 13584 8916 13590 8968
rect 15737 8959 15795 8965
rect 15737 8925 15749 8959
rect 15783 8956 15795 8959
rect 16562 8956 16568 8968
rect 15783 8928 16568 8956
rect 15783 8925 15795 8928
rect 15737 8919 15795 8925
rect 16562 8916 16568 8928
rect 16620 8916 16626 8968
rect 18402 8956 18408 8968
rect 18363 8928 18408 8956
rect 18402 8916 18408 8928
rect 18460 8916 18466 8968
rect 18770 8956 18776 8968
rect 18731 8928 18776 8956
rect 18770 8916 18776 8928
rect 18828 8916 18834 8968
rect 23002 8956 23008 8968
rect 22963 8928 23008 8956
rect 23002 8916 23008 8928
rect 23060 8916 23066 8968
rect 12882 8848 12888 8900
rect 12940 8888 12946 8900
rect 13326 8891 13384 8897
rect 13326 8888 13338 8891
rect 12940 8860 13338 8888
rect 12940 8848 12946 8860
rect 13326 8857 13338 8860
rect 13372 8888 13384 8891
rect 14262 8888 14268 8900
rect 13372 8860 14268 8888
rect 13372 8857 13384 8860
rect 13326 8851 13384 8857
rect 14262 8848 14268 8860
rect 14320 8848 14326 8900
rect 23554 8888 23560 8900
rect 23515 8860 23560 8888
rect 23554 8848 23560 8860
rect 23612 8848 23618 8900
rect 13437 8823 13495 8829
rect 13437 8789 13449 8823
rect 13483 8820 13495 8823
rect 13618 8820 13624 8832
rect 13483 8792 13624 8820
rect 13483 8789 13495 8792
rect 13437 8783 13495 8789
rect 13618 8780 13624 8792
rect 13676 8780 13682 8832
rect 16378 8820 16384 8832
rect 16339 8792 16384 8820
rect 16378 8780 16384 8792
rect 16436 8780 16442 8832
rect 17485 8823 17543 8829
rect 17485 8789 17497 8823
rect 17531 8820 17543 8823
rect 17666 8820 17672 8832
rect 17531 8792 17672 8820
rect 17531 8789 17543 8792
rect 17485 8783 17543 8789
rect 17666 8780 17672 8792
rect 17724 8780 17730 8832
rect 21622 8780 21628 8832
rect 21680 8820 21686 8832
rect 21680 8792 21725 8820
rect 21680 8780 21686 8792
rect 23278 8780 23284 8832
rect 23336 8820 23342 8832
rect 23925 8823 23983 8829
rect 23925 8820 23937 8823
rect 23336 8792 23937 8820
rect 23336 8780 23342 8792
rect 23925 8789 23937 8792
rect 23971 8789 23983 8823
rect 23925 8783 23983 8789
rect 632 8730 26392 8752
rect 632 8678 5176 8730
rect 5228 8678 5240 8730
rect 5292 8678 5304 8730
rect 5356 8678 5368 8730
rect 5420 8678 14510 8730
rect 14562 8678 14574 8730
rect 14626 8678 14638 8730
rect 14690 8678 14702 8730
rect 14754 8678 23843 8730
rect 23895 8678 23907 8730
rect 23959 8678 23971 8730
rect 24023 8678 24035 8730
rect 24087 8678 26392 8730
rect 632 8656 26392 8678
rect 12882 8616 12888 8628
rect 12843 8588 12888 8616
rect 12882 8576 12888 8588
rect 12940 8576 12946 8628
rect 13526 8576 13532 8628
rect 13584 8616 13590 8628
rect 13621 8619 13679 8625
rect 13621 8616 13633 8619
rect 13584 8588 13633 8616
rect 13584 8576 13590 8588
rect 13621 8585 13633 8588
rect 13667 8616 13679 8619
rect 15274 8616 15280 8628
rect 13667 8588 15280 8616
rect 13667 8585 13679 8588
rect 13621 8579 13679 8585
rect 15274 8576 15280 8588
rect 15332 8576 15338 8628
rect 15458 8616 15464 8628
rect 15419 8588 15464 8616
rect 15458 8576 15464 8588
rect 15516 8576 15522 8628
rect 15734 8616 15740 8628
rect 15695 8588 15740 8616
rect 15734 8576 15740 8588
rect 15792 8576 15798 8628
rect 16746 8576 16752 8628
rect 16804 8616 16810 8628
rect 16933 8619 16991 8625
rect 16933 8616 16945 8619
rect 16804 8588 16945 8616
rect 16804 8576 16810 8588
rect 16933 8585 16945 8588
rect 16979 8616 16991 8619
rect 17301 8619 17359 8625
rect 17301 8616 17313 8619
rect 16979 8588 17313 8616
rect 16979 8585 16991 8588
rect 16933 8579 16991 8585
rect 17301 8585 17313 8588
rect 17347 8585 17359 8619
rect 17301 8579 17359 8585
rect 18497 8619 18555 8625
rect 18497 8585 18509 8619
rect 18543 8616 18555 8619
rect 18862 8616 18868 8628
rect 18543 8588 18868 8616
rect 18543 8585 18555 8588
rect 18497 8579 18555 8585
rect 13253 8483 13311 8489
rect 13253 8449 13265 8483
rect 13299 8480 13311 8483
rect 13618 8480 13624 8492
rect 13299 8452 13624 8480
rect 13299 8449 13311 8452
rect 13253 8443 13311 8449
rect 13618 8440 13624 8452
rect 13676 8440 13682 8492
rect 17316 8480 17344 8579
rect 18862 8576 18868 8588
rect 18920 8576 18926 8628
rect 18954 8576 18960 8628
rect 19012 8616 19018 8628
rect 19141 8619 19199 8625
rect 19141 8616 19153 8619
rect 19012 8588 19153 8616
rect 19012 8576 19018 8588
rect 19141 8585 19153 8588
rect 19187 8585 19199 8619
rect 19141 8579 19199 8585
rect 20429 8619 20487 8625
rect 20429 8585 20441 8619
rect 20475 8616 20487 8619
rect 20702 8616 20708 8628
rect 20475 8588 20708 8616
rect 20475 8585 20487 8588
rect 20429 8579 20487 8585
rect 17316 8452 17712 8480
rect 14354 8412 14360 8424
rect 14315 8384 14360 8412
rect 14354 8372 14360 8384
rect 14412 8372 14418 8424
rect 14906 8372 14912 8424
rect 14964 8412 14970 8424
rect 15001 8415 15059 8421
rect 15001 8412 15013 8415
rect 14964 8384 15013 8412
rect 14964 8372 14970 8384
rect 15001 8381 15013 8384
rect 15047 8381 15059 8415
rect 15001 8375 15059 8381
rect 15734 8372 15740 8424
rect 15792 8412 15798 8424
rect 15921 8415 15979 8421
rect 15921 8412 15933 8415
rect 15792 8384 15933 8412
rect 15792 8372 15798 8384
rect 15921 8381 15933 8384
rect 15967 8412 15979 8415
rect 16194 8412 16200 8424
rect 15967 8384 16200 8412
rect 15967 8381 15979 8384
rect 15921 8375 15979 8381
rect 16194 8372 16200 8384
rect 16252 8372 16258 8424
rect 16378 8412 16384 8424
rect 16339 8384 16384 8412
rect 16378 8372 16384 8384
rect 16436 8372 16442 8424
rect 16657 8415 16715 8421
rect 16657 8381 16669 8415
rect 16703 8412 16715 8415
rect 17574 8412 17580 8424
rect 16703 8384 17580 8412
rect 16703 8381 16715 8384
rect 16657 8375 16715 8381
rect 17574 8372 17580 8384
rect 17632 8372 17638 8424
rect 13250 8304 13256 8356
rect 13308 8344 13314 8356
rect 13713 8347 13771 8353
rect 13713 8344 13725 8347
rect 13308 8316 13725 8344
rect 13308 8304 13314 8316
rect 13713 8313 13725 8316
rect 13759 8313 13771 8347
rect 15090 8344 15096 8356
rect 13713 8307 13771 8313
rect 14740 8316 15096 8344
rect 13802 8236 13808 8288
rect 13860 8276 13866 8288
rect 14740 8276 14768 8316
rect 15090 8304 15096 8316
rect 15148 8304 15154 8356
rect 17684 8344 17712 8452
rect 17758 8344 17764 8356
rect 17671 8316 17764 8344
rect 17758 8304 17764 8316
rect 17816 8344 17822 8356
rect 17898 8347 17956 8353
rect 17898 8344 17910 8347
rect 17816 8316 17910 8344
rect 17816 8304 17822 8316
rect 17898 8313 17910 8316
rect 17944 8313 17956 8347
rect 19156 8344 19184 8579
rect 20702 8576 20708 8588
rect 20760 8576 20766 8628
rect 20797 8619 20855 8625
rect 20797 8585 20809 8619
rect 20843 8616 20855 8619
rect 21254 8616 21260 8628
rect 20843 8588 21260 8616
rect 20843 8585 20855 8588
rect 20797 8579 20855 8585
rect 21254 8576 21260 8588
rect 21312 8576 21318 8628
rect 22637 8619 22695 8625
rect 22637 8585 22649 8619
rect 22683 8616 22695 8619
rect 22818 8616 22824 8628
rect 22683 8588 22824 8616
rect 22683 8585 22695 8588
rect 22637 8579 22695 8585
rect 22818 8576 22824 8588
rect 22876 8616 22882 8628
rect 23002 8616 23008 8628
rect 22876 8588 23008 8616
rect 22876 8576 22882 8588
rect 23002 8576 23008 8588
rect 23060 8576 23066 8628
rect 24934 8616 24940 8628
rect 24895 8588 24940 8616
rect 24934 8576 24940 8588
rect 24992 8576 24998 8628
rect 19417 8483 19475 8489
rect 19417 8449 19429 8483
rect 19463 8480 19475 8483
rect 19506 8480 19512 8492
rect 19463 8452 19512 8480
rect 19463 8449 19475 8452
rect 19417 8443 19475 8449
rect 19506 8440 19512 8452
rect 19564 8440 19570 8492
rect 19690 8480 19696 8492
rect 19651 8452 19696 8480
rect 19690 8440 19696 8452
rect 19748 8440 19754 8492
rect 21349 8483 21407 8489
rect 21349 8449 21361 8483
rect 21395 8480 21407 8483
rect 21530 8480 21536 8492
rect 21395 8452 21536 8480
rect 21395 8449 21407 8452
rect 21349 8443 21407 8449
rect 21530 8440 21536 8452
rect 21588 8440 21594 8492
rect 23278 8480 23284 8492
rect 23239 8452 23284 8480
rect 23278 8440 23284 8452
rect 23336 8440 23342 8492
rect 23554 8480 23560 8492
rect 23515 8452 23560 8480
rect 23554 8440 23560 8452
rect 23612 8440 23618 8492
rect 22269 8415 22327 8421
rect 22269 8381 22281 8415
rect 22315 8381 22327 8415
rect 24750 8412 24756 8424
rect 24711 8384 24756 8412
rect 22269 8375 22327 8381
rect 19509 8347 19567 8353
rect 19509 8344 19521 8347
rect 19156 8316 19521 8344
rect 17898 8307 17956 8313
rect 19509 8313 19521 8316
rect 19555 8313 19567 8347
rect 19509 8307 19567 8313
rect 21254 8304 21260 8356
rect 21312 8344 21318 8356
rect 21670 8347 21728 8353
rect 21670 8344 21682 8347
rect 21312 8316 21682 8344
rect 21312 8304 21318 8316
rect 21670 8313 21682 8316
rect 21716 8313 21728 8347
rect 22284 8344 22312 8375
rect 24750 8372 24756 8384
rect 24808 8412 24814 8424
rect 25305 8415 25363 8421
rect 25305 8412 25317 8415
rect 24808 8384 25317 8412
rect 24808 8372 24814 8384
rect 25305 8381 25317 8384
rect 25351 8381 25363 8415
rect 25305 8375 25363 8381
rect 23370 8344 23376 8356
rect 22284 8316 23376 8344
rect 21670 8307 21728 8313
rect 23370 8304 23376 8316
rect 23428 8344 23434 8356
rect 24201 8347 24259 8353
rect 24201 8344 24213 8347
rect 23428 8316 24213 8344
rect 23428 8304 23434 8316
rect 24201 8313 24213 8316
rect 24247 8313 24259 8347
rect 24201 8307 24259 8313
rect 24382 8304 24388 8356
rect 24440 8344 24446 8356
rect 24569 8347 24627 8353
rect 24569 8344 24581 8347
rect 24440 8316 24581 8344
rect 24440 8304 24446 8316
rect 24569 8313 24581 8316
rect 24615 8313 24627 8347
rect 24569 8307 24627 8313
rect 13860 8248 14768 8276
rect 13860 8236 13866 8248
rect 17666 8236 17672 8288
rect 17724 8276 17730 8288
rect 18773 8279 18831 8285
rect 18773 8276 18785 8279
rect 17724 8248 18785 8276
rect 17724 8236 17730 8248
rect 18773 8245 18785 8248
rect 18819 8245 18831 8279
rect 18773 8239 18831 8245
rect 23005 8279 23063 8285
rect 23005 8245 23017 8279
rect 23051 8276 23063 8279
rect 23094 8276 23100 8288
rect 23051 8248 23100 8276
rect 23051 8245 23063 8248
rect 23005 8239 23063 8245
rect 23094 8236 23100 8248
rect 23152 8236 23158 8288
rect 632 8186 26392 8208
rect 632 8134 9843 8186
rect 9895 8134 9907 8186
rect 9959 8134 9971 8186
rect 10023 8134 10035 8186
rect 10087 8134 19176 8186
rect 19228 8134 19240 8186
rect 19292 8134 19304 8186
rect 19356 8134 19368 8186
rect 19420 8134 26392 8186
rect 632 8112 26392 8134
rect 13250 8072 13256 8084
rect 13211 8044 13256 8072
rect 13250 8032 13256 8044
rect 13308 8032 13314 8084
rect 13805 8075 13863 8081
rect 13805 8041 13817 8075
rect 13851 8072 13863 8075
rect 14354 8072 14360 8084
rect 13851 8044 14360 8072
rect 13851 8041 13863 8044
rect 13805 8035 13863 8041
rect 14354 8032 14360 8044
rect 14412 8032 14418 8084
rect 16562 8032 16568 8084
rect 16620 8072 16626 8084
rect 16933 8075 16991 8081
rect 16933 8072 16945 8075
rect 16620 8044 16945 8072
rect 16620 8032 16626 8044
rect 16933 8041 16945 8044
rect 16979 8041 16991 8075
rect 17574 8072 17580 8084
rect 17535 8044 17580 8072
rect 16933 8035 16991 8041
rect 17574 8032 17580 8044
rect 17632 8032 17638 8084
rect 18313 8075 18371 8081
rect 18313 8041 18325 8075
rect 18359 8072 18371 8075
rect 18402 8072 18408 8084
rect 18359 8044 18408 8072
rect 18359 8041 18371 8044
rect 18313 8035 18371 8041
rect 18402 8032 18408 8044
rect 18460 8032 18466 8084
rect 24658 8032 24664 8084
rect 24716 8072 24722 8084
rect 24753 8075 24811 8081
rect 24753 8072 24765 8075
rect 24716 8044 24765 8072
rect 24716 8032 24722 8044
rect 24753 8041 24765 8044
rect 24799 8041 24811 8075
rect 24753 8035 24811 8041
rect 14173 8007 14231 8013
rect 14173 7973 14185 8007
rect 14219 8004 14231 8007
rect 14998 8004 15004 8016
rect 14219 7976 15004 8004
rect 14219 7973 14231 7976
rect 14173 7967 14231 7973
rect 14998 7964 15004 7976
rect 15056 7964 15062 8016
rect 18586 8004 18592 8016
rect 18547 7976 18592 8004
rect 18586 7964 18592 7976
rect 18644 7964 18650 8016
rect 21622 7964 21628 8016
rect 21680 8004 21686 8016
rect 23186 8004 23192 8016
rect 21680 7976 21725 8004
rect 23147 7976 23192 8004
rect 21680 7964 21686 7976
rect 23186 7964 23192 7976
rect 23244 7964 23250 8016
rect 16102 7896 16108 7948
rect 16160 7936 16166 7948
rect 16470 7936 16476 7948
rect 16160 7908 16205 7936
rect 16431 7908 16476 7936
rect 16160 7896 16166 7908
rect 16470 7896 16476 7908
rect 16528 7896 16534 7948
rect 24566 7936 24572 7948
rect 24527 7908 24572 7936
rect 24566 7896 24572 7908
rect 24624 7896 24630 7948
rect 16657 7871 16715 7877
rect 16657 7837 16669 7871
rect 16703 7868 16715 7871
rect 17482 7868 17488 7880
rect 16703 7840 17488 7868
rect 16703 7837 16715 7840
rect 16657 7831 16715 7837
rect 17482 7828 17488 7840
rect 17540 7828 17546 7880
rect 18494 7868 18500 7880
rect 18455 7840 18500 7868
rect 18494 7828 18500 7840
rect 18552 7828 18558 7880
rect 18862 7868 18868 7880
rect 18823 7840 18868 7868
rect 18862 7828 18868 7840
rect 18920 7828 18926 7880
rect 20978 7828 20984 7880
rect 21036 7868 21042 7880
rect 21533 7871 21591 7877
rect 21533 7868 21545 7871
rect 21036 7840 21545 7868
rect 21036 7828 21042 7840
rect 21533 7837 21545 7840
rect 21579 7837 21591 7871
rect 23094 7868 23100 7880
rect 23055 7840 23100 7868
rect 21533 7831 21591 7837
rect 23094 7828 23100 7840
rect 23152 7828 23158 7880
rect 23278 7828 23284 7880
rect 23336 7868 23342 7880
rect 23373 7871 23431 7877
rect 23373 7868 23385 7871
rect 23336 7840 23385 7868
rect 23336 7828 23342 7840
rect 23373 7837 23385 7840
rect 23419 7837 23431 7871
rect 23373 7831 23431 7837
rect 22085 7803 22143 7809
rect 22085 7769 22097 7803
rect 22131 7800 22143 7803
rect 23296 7800 23324 7828
rect 22131 7772 23324 7800
rect 22131 7769 22143 7772
rect 22085 7763 22143 7769
rect 15366 7732 15372 7744
rect 15327 7704 15372 7732
rect 15366 7692 15372 7704
rect 15424 7692 15430 7744
rect 15550 7692 15556 7744
rect 15608 7732 15614 7744
rect 15737 7735 15795 7741
rect 15737 7732 15749 7735
rect 15608 7704 15749 7732
rect 15608 7692 15614 7704
rect 15737 7701 15749 7704
rect 15783 7701 15795 7735
rect 15737 7695 15795 7701
rect 632 7642 26392 7664
rect 632 7590 5176 7642
rect 5228 7590 5240 7642
rect 5292 7590 5304 7642
rect 5356 7590 5368 7642
rect 5420 7590 14510 7642
rect 14562 7590 14574 7642
rect 14626 7590 14638 7642
rect 14690 7590 14702 7642
rect 14754 7590 23843 7642
rect 23895 7590 23907 7642
rect 23959 7590 23971 7642
rect 24023 7590 24035 7642
rect 24087 7590 26392 7642
rect 632 7568 26392 7590
rect 15185 7531 15243 7537
rect 15185 7528 15197 7531
rect 14096 7500 15197 7528
rect 13618 7420 13624 7472
rect 13676 7460 13682 7472
rect 14096 7469 14124 7500
rect 15185 7497 15197 7500
rect 15231 7528 15243 7531
rect 15645 7531 15703 7537
rect 15645 7528 15657 7531
rect 15231 7500 15657 7528
rect 15231 7497 15243 7500
rect 15185 7491 15243 7497
rect 15645 7497 15657 7500
rect 15691 7497 15703 7531
rect 15645 7491 15703 7497
rect 16102 7488 16108 7540
rect 16160 7528 16166 7540
rect 16381 7531 16439 7537
rect 16381 7528 16393 7531
rect 16160 7500 16393 7528
rect 16160 7488 16166 7500
rect 16381 7497 16393 7500
rect 16427 7497 16439 7531
rect 20978 7528 20984 7540
rect 20939 7500 20984 7528
rect 16381 7491 16439 7497
rect 20978 7488 20984 7500
rect 21036 7488 21042 7540
rect 21441 7531 21499 7537
rect 21441 7497 21453 7531
rect 21487 7528 21499 7531
rect 21622 7528 21628 7540
rect 21487 7500 21628 7528
rect 21487 7497 21499 7500
rect 21441 7491 21499 7497
rect 21622 7488 21628 7500
rect 21680 7488 21686 7540
rect 21993 7531 22051 7537
rect 21993 7497 22005 7531
rect 22039 7528 22051 7531
rect 23005 7531 23063 7537
rect 23005 7528 23017 7531
rect 22039 7500 23017 7528
rect 22039 7497 22051 7500
rect 21993 7491 22051 7497
rect 23005 7497 23017 7500
rect 23051 7528 23063 7531
rect 23186 7528 23192 7540
rect 23051 7500 23192 7528
rect 23051 7497 23063 7500
rect 23005 7491 23063 7497
rect 23186 7488 23192 7500
rect 23244 7488 23250 7540
rect 24198 7488 24204 7540
rect 24256 7528 24262 7540
rect 24937 7531 24995 7537
rect 24937 7528 24949 7531
rect 24256 7500 24949 7528
rect 24256 7488 24262 7500
rect 24937 7497 24949 7500
rect 24983 7497 24995 7531
rect 24937 7491 24995 7497
rect 14081 7463 14139 7469
rect 14081 7460 14093 7463
rect 13676 7432 14093 7460
rect 13676 7420 13682 7432
rect 14081 7429 14093 7432
rect 14127 7429 14139 7463
rect 14909 7463 14967 7469
rect 14909 7460 14921 7463
rect 14081 7423 14139 7429
rect 14188 7432 14921 7460
rect 14188 7401 14216 7432
rect 14909 7429 14921 7432
rect 14955 7460 14967 7463
rect 14998 7460 15004 7472
rect 14955 7432 15004 7460
rect 14955 7429 14967 7432
rect 14909 7423 14967 7429
rect 14998 7420 15004 7432
rect 15056 7420 15062 7472
rect 15550 7469 15556 7472
rect 15534 7463 15556 7469
rect 15534 7429 15546 7463
rect 15534 7423 15556 7429
rect 15550 7420 15556 7423
rect 15608 7420 15614 7472
rect 12609 7395 12667 7401
rect 12609 7361 12621 7395
rect 12655 7392 12667 7395
rect 13253 7395 13311 7401
rect 13253 7392 13265 7395
rect 12655 7364 13265 7392
rect 12655 7361 12667 7364
rect 12609 7355 12667 7361
rect 13253 7361 13265 7364
rect 13299 7361 13311 7395
rect 13253 7355 13311 7361
rect 14173 7395 14231 7401
rect 14173 7361 14185 7395
rect 14219 7361 14231 7395
rect 15016 7392 15044 7420
rect 15737 7395 15795 7401
rect 15737 7392 15749 7395
rect 15016 7364 15749 7392
rect 14173 7355 14231 7361
rect 15737 7361 15749 7364
rect 15783 7361 15795 7395
rect 15737 7355 15795 7361
rect 18497 7395 18555 7401
rect 18497 7361 18509 7395
rect 18543 7392 18555 7395
rect 18586 7392 18592 7404
rect 18543 7364 18592 7392
rect 18543 7361 18555 7364
rect 18497 7355 18555 7361
rect 12238 7324 12244 7336
rect 12151 7296 12244 7324
rect 12238 7284 12244 7296
rect 12296 7324 12302 7336
rect 12885 7327 12943 7333
rect 12885 7324 12897 7327
rect 12296 7296 12897 7324
rect 12296 7284 12302 7296
rect 12885 7293 12897 7296
rect 12931 7293 12943 7327
rect 12885 7287 12943 7293
rect 11781 7259 11839 7265
rect 11781 7225 11793 7259
rect 11827 7256 11839 7259
rect 12054 7256 12060 7268
rect 11827 7228 12060 7256
rect 11827 7225 11839 7228
rect 11781 7219 11839 7225
rect 12054 7216 12060 7228
rect 12112 7216 12118 7268
rect 13268 7256 13296 7355
rect 18586 7352 18592 7364
rect 18644 7392 18650 7404
rect 18773 7395 18831 7401
rect 18773 7392 18785 7395
rect 18644 7364 18785 7392
rect 18644 7352 18650 7364
rect 18773 7361 18785 7364
rect 18819 7361 18831 7395
rect 18773 7355 18831 7361
rect 23002 7352 23008 7404
rect 23060 7392 23066 7404
rect 23189 7395 23247 7401
rect 23189 7392 23201 7395
rect 23060 7364 23201 7392
rect 23060 7352 23066 7364
rect 23189 7361 23201 7364
rect 23235 7361 23247 7395
rect 23189 7355 23247 7361
rect 13952 7327 14010 7333
rect 13952 7293 13964 7327
rect 13998 7324 14010 7327
rect 14078 7324 14084 7336
rect 13998 7296 14084 7324
rect 13998 7293 14010 7296
rect 13952 7287 14010 7293
rect 14078 7284 14084 7296
rect 14136 7324 14142 7336
rect 15550 7324 15556 7336
rect 14136 7296 15556 7324
rect 14136 7284 14142 7296
rect 15550 7284 15556 7296
rect 15608 7284 15614 7336
rect 17393 7327 17451 7333
rect 17393 7293 17405 7327
rect 17439 7324 17451 7327
rect 17666 7324 17672 7336
rect 17439 7296 17672 7324
rect 17439 7293 17451 7296
rect 17393 7287 17451 7293
rect 17666 7284 17672 7296
rect 17724 7324 17730 7336
rect 17853 7327 17911 7333
rect 17853 7324 17865 7327
rect 17724 7296 17865 7324
rect 17724 7284 17730 7296
rect 17853 7293 17865 7296
rect 17899 7293 17911 7327
rect 17853 7287 17911 7293
rect 21622 7284 21628 7336
rect 21680 7324 21686 7336
rect 23370 7324 23376 7336
rect 21680 7296 21725 7324
rect 23331 7296 23376 7324
rect 21680 7284 21686 7296
rect 23370 7284 23376 7296
rect 23428 7284 23434 7336
rect 24474 7284 24480 7336
rect 24532 7324 24538 7336
rect 24753 7327 24811 7333
rect 24753 7324 24765 7327
rect 24532 7296 24765 7324
rect 24532 7284 24538 7296
rect 24753 7293 24765 7296
rect 24799 7324 24811 7327
rect 25305 7327 25363 7333
rect 25305 7324 25317 7327
rect 24799 7296 25317 7324
rect 24799 7293 24811 7296
rect 24753 7287 24811 7293
rect 25305 7293 25317 7296
rect 25351 7293 25363 7327
rect 25305 7287 25363 7293
rect 13802 7256 13808 7268
rect 13268 7228 13808 7256
rect 13802 7216 13808 7228
rect 13860 7216 13866 7268
rect 15366 7256 15372 7268
rect 15327 7228 15372 7256
rect 15366 7216 15372 7228
rect 15424 7216 15430 7268
rect 16105 7259 16163 7265
rect 16105 7225 16117 7259
rect 16151 7225 16163 7259
rect 16105 7219 16163 7225
rect 22637 7259 22695 7265
rect 22637 7225 22649 7259
rect 22683 7256 22695 7259
rect 23094 7256 23100 7268
rect 22683 7228 23100 7256
rect 22683 7225 22695 7228
rect 22637 7219 22695 7225
rect 13618 7188 13624 7200
rect 13579 7160 13624 7188
rect 13618 7148 13624 7160
rect 13676 7148 13682 7200
rect 14354 7148 14360 7200
rect 14412 7188 14418 7200
rect 14449 7191 14507 7197
rect 14449 7188 14461 7191
rect 14412 7160 14461 7188
rect 14412 7148 14418 7160
rect 14449 7157 14461 7160
rect 14495 7157 14507 7191
rect 16120 7188 16148 7219
rect 23094 7216 23100 7228
rect 23152 7256 23158 7268
rect 24382 7256 24388 7268
rect 23152 7228 24388 7256
rect 23152 7216 23158 7228
rect 24382 7216 24388 7228
rect 24440 7216 24446 7268
rect 16470 7188 16476 7200
rect 16120 7160 16476 7188
rect 14449 7151 14507 7157
rect 16470 7148 16476 7160
rect 16528 7188 16534 7200
rect 16841 7191 16899 7197
rect 16841 7188 16853 7191
rect 16528 7160 16853 7188
rect 16528 7148 16534 7160
rect 16841 7157 16853 7160
rect 16887 7188 16899 7191
rect 16930 7188 16936 7200
rect 16887 7160 16936 7188
rect 16887 7157 16899 7160
rect 16841 7151 16899 7157
rect 16930 7148 16936 7160
rect 16988 7148 16994 7200
rect 18494 7148 18500 7200
rect 18552 7188 18558 7200
rect 19233 7191 19291 7197
rect 19233 7188 19245 7191
rect 18552 7160 19245 7188
rect 18552 7148 18558 7160
rect 19233 7157 19245 7160
rect 19279 7188 19291 7191
rect 19598 7188 19604 7200
rect 19279 7160 19604 7188
rect 19279 7157 19291 7160
rect 19233 7151 19291 7157
rect 19598 7148 19604 7160
rect 19656 7148 19662 7200
rect 20153 7191 20211 7197
rect 20153 7157 20165 7191
rect 20199 7188 20211 7191
rect 20242 7188 20248 7200
rect 20199 7160 20248 7188
rect 20199 7157 20211 7160
rect 20153 7151 20211 7157
rect 20242 7148 20248 7160
rect 20300 7148 20306 7200
rect 24198 7148 24204 7200
rect 24256 7188 24262 7200
rect 24566 7188 24572 7200
rect 24256 7160 24572 7188
rect 24256 7148 24262 7160
rect 24566 7148 24572 7160
rect 24624 7148 24630 7200
rect 632 7098 26392 7120
rect 632 7046 9843 7098
rect 9895 7046 9907 7098
rect 9959 7046 9971 7098
rect 10023 7046 10035 7098
rect 10087 7046 19176 7098
rect 19228 7046 19240 7098
rect 19292 7046 19304 7098
rect 19356 7046 19368 7098
rect 19420 7046 26392 7098
rect 632 7024 26392 7046
rect 15366 6984 15372 6996
rect 13268 6956 15372 6984
rect 12072 6888 12376 6916
rect 11870 6848 11876 6860
rect 11831 6820 11876 6848
rect 11870 6808 11876 6820
rect 11928 6808 11934 6860
rect 11965 6851 12023 6857
rect 11965 6817 11977 6851
rect 12011 6848 12023 6851
rect 12072 6848 12100 6888
rect 12011 6820 12100 6848
rect 12149 6851 12207 6857
rect 12011 6817 12023 6820
rect 11965 6811 12023 6817
rect 12149 6817 12161 6851
rect 12195 6848 12207 6851
rect 12238 6848 12244 6860
rect 12195 6820 12244 6848
rect 12195 6817 12207 6820
rect 12149 6811 12207 6817
rect 11594 6740 11600 6792
rect 11652 6780 11658 6792
rect 12164 6780 12192 6811
rect 12238 6808 12244 6820
rect 12296 6808 12302 6860
rect 12348 6848 12376 6888
rect 13268 6848 13296 6956
rect 15366 6944 15372 6956
rect 15424 6944 15430 6996
rect 21622 6944 21628 6996
rect 21680 6984 21686 6996
rect 23370 6984 23376 6996
rect 21680 6956 21725 6984
rect 23331 6956 23376 6984
rect 21680 6944 21686 6956
rect 23370 6944 23376 6956
rect 23428 6944 23434 6996
rect 14078 6876 14084 6928
rect 14136 6916 14142 6928
rect 14173 6919 14231 6925
rect 14173 6916 14185 6919
rect 14136 6888 14185 6916
rect 14136 6876 14142 6888
rect 14173 6885 14185 6888
rect 14219 6885 14231 6919
rect 17114 6916 17120 6928
rect 17075 6888 17120 6916
rect 14173 6879 14231 6885
rect 17114 6876 17120 6888
rect 17172 6876 17178 6928
rect 18862 6916 18868 6928
rect 18823 6888 18868 6916
rect 18862 6876 18868 6888
rect 18920 6876 18926 6928
rect 13434 6848 13440 6860
rect 12348 6820 13296 6848
rect 13395 6820 13440 6848
rect 13434 6808 13440 6820
rect 13492 6808 13498 6860
rect 13713 6851 13771 6857
rect 13713 6817 13725 6851
rect 13759 6848 13771 6851
rect 14354 6848 14360 6860
rect 13759 6820 14360 6848
rect 13759 6817 13771 6820
rect 13713 6811 13771 6817
rect 14354 6808 14360 6820
rect 14412 6808 14418 6860
rect 15090 6848 15096 6860
rect 15051 6820 15096 6848
rect 15090 6808 15096 6820
rect 15148 6808 15154 6860
rect 15182 6808 15188 6860
rect 15240 6848 15246 6860
rect 15277 6851 15335 6857
rect 15277 6848 15289 6851
rect 15240 6820 15289 6848
rect 15240 6808 15246 6820
rect 15277 6817 15289 6820
rect 15323 6817 15335 6851
rect 15277 6811 15335 6817
rect 16194 6808 16200 6860
rect 16252 6848 16258 6860
rect 16562 6848 16568 6860
rect 16252 6820 16568 6848
rect 16252 6808 16258 6820
rect 16562 6808 16568 6820
rect 16620 6808 16626 6860
rect 16930 6848 16936 6860
rect 16891 6820 16936 6848
rect 16930 6808 16936 6820
rect 16988 6808 16994 6860
rect 18494 6848 18500 6860
rect 18455 6820 18500 6848
rect 18494 6808 18500 6820
rect 18552 6808 18558 6860
rect 21070 6848 21076 6860
rect 21031 6820 21076 6848
rect 21070 6808 21076 6820
rect 21128 6808 21134 6860
rect 22818 6848 22824 6860
rect 22779 6820 22824 6848
rect 22818 6808 22824 6820
rect 22876 6808 22882 6860
rect 23554 6808 23560 6860
rect 23612 6848 23618 6860
rect 23868 6851 23926 6857
rect 23868 6848 23880 6851
rect 23612 6820 23880 6848
rect 23612 6808 23618 6820
rect 23868 6817 23880 6820
rect 23914 6817 23926 6851
rect 23868 6811 23926 6817
rect 23971 6851 24029 6857
rect 23971 6817 23983 6851
rect 24017 6848 24029 6851
rect 24290 6848 24296 6860
rect 24017 6820 24296 6848
rect 24017 6817 24029 6820
rect 23971 6811 24029 6817
rect 24290 6808 24296 6820
rect 24348 6808 24354 6860
rect 24912 6851 24970 6857
rect 24912 6817 24924 6851
rect 24958 6848 24970 6851
rect 25118 6848 25124 6860
rect 24958 6820 25124 6848
rect 24958 6817 24970 6820
rect 24912 6811 24970 6817
rect 25118 6808 25124 6820
rect 25176 6808 25182 6860
rect 13894 6780 13900 6792
rect 11652 6752 12192 6780
rect 13855 6752 13900 6780
rect 11652 6740 11658 6752
rect 13894 6740 13900 6752
rect 13952 6740 13958 6792
rect 15366 6740 15372 6792
rect 15424 6780 15430 6792
rect 15553 6783 15611 6789
rect 15553 6780 15565 6783
rect 15424 6752 15565 6780
rect 15424 6740 15430 6752
rect 15553 6749 15565 6752
rect 15599 6780 15611 6783
rect 15829 6783 15887 6789
rect 15829 6780 15841 6783
rect 15599 6752 15841 6780
rect 15599 6749 15611 6752
rect 15553 6743 15611 6749
rect 15829 6749 15841 6752
rect 15875 6749 15887 6783
rect 18512 6780 18540 6808
rect 18773 6783 18831 6789
rect 18773 6780 18785 6783
rect 18512 6752 18785 6780
rect 15829 6743 15887 6749
rect 18773 6749 18785 6752
rect 18819 6749 18831 6783
rect 18773 6743 18831 6749
rect 19417 6783 19475 6789
rect 19417 6749 19429 6783
rect 19463 6780 19475 6783
rect 19874 6780 19880 6792
rect 19463 6752 19880 6780
rect 19463 6749 19475 6752
rect 19417 6743 19475 6749
rect 19874 6740 19880 6752
rect 19932 6740 19938 6792
rect 24382 6672 24388 6724
rect 24440 6712 24446 6724
rect 24983 6715 25041 6721
rect 24983 6712 24995 6715
rect 24440 6684 24995 6712
rect 24440 6672 24446 6684
rect 24983 6681 24995 6684
rect 25029 6681 25041 6715
rect 24983 6675 25041 6681
rect 20886 6644 20892 6656
rect 20847 6616 20892 6644
rect 20886 6604 20892 6616
rect 20944 6604 20950 6656
rect 632 6554 26392 6576
rect 632 6502 5176 6554
rect 5228 6502 5240 6554
rect 5292 6502 5304 6554
rect 5356 6502 5368 6554
rect 5420 6502 14510 6554
rect 14562 6502 14574 6554
rect 14626 6502 14638 6554
rect 14690 6502 14702 6554
rect 14754 6502 23843 6554
rect 23895 6502 23907 6554
rect 23959 6502 23971 6554
rect 24023 6502 24035 6554
rect 24087 6502 26392 6554
rect 632 6480 26392 6502
rect 12054 6400 12060 6452
rect 12112 6440 12118 6452
rect 12241 6443 12299 6449
rect 12241 6440 12253 6443
rect 12112 6412 12253 6440
rect 12112 6400 12118 6412
rect 12241 6409 12253 6412
rect 12287 6409 12299 6443
rect 12241 6403 12299 6409
rect 13434 6400 13440 6452
rect 13492 6440 13498 6452
rect 13529 6443 13587 6449
rect 13529 6440 13541 6443
rect 13492 6412 13541 6440
rect 13492 6400 13498 6412
rect 13529 6409 13541 6412
rect 13575 6409 13587 6443
rect 13529 6403 13587 6409
rect 14909 6443 14967 6449
rect 14909 6409 14921 6443
rect 14955 6440 14967 6443
rect 15090 6440 15096 6452
rect 14955 6412 15096 6440
rect 14955 6409 14967 6412
rect 14909 6403 14967 6409
rect 15090 6400 15096 6412
rect 15148 6440 15154 6452
rect 16562 6440 16568 6452
rect 15148 6412 16568 6440
rect 15148 6400 15154 6412
rect 16562 6400 16568 6412
rect 16620 6400 16626 6452
rect 16930 6440 16936 6452
rect 16891 6412 16936 6440
rect 16930 6400 16936 6412
rect 16988 6400 16994 6452
rect 18497 6443 18555 6449
rect 18497 6409 18509 6443
rect 18543 6440 18555 6443
rect 18862 6440 18868 6452
rect 18543 6412 18868 6440
rect 18543 6409 18555 6412
rect 18497 6403 18555 6409
rect 18862 6400 18868 6412
rect 18920 6400 18926 6452
rect 20242 6400 20248 6452
rect 20300 6440 20306 6452
rect 20521 6443 20579 6449
rect 20521 6440 20533 6443
rect 20300 6412 20533 6440
rect 20300 6400 20306 6412
rect 20521 6409 20533 6412
rect 20567 6409 20579 6443
rect 20886 6440 20892 6452
rect 20847 6412 20892 6440
rect 20521 6403 20579 6409
rect 13253 6375 13311 6381
rect 13253 6341 13265 6375
rect 13299 6372 13311 6375
rect 14354 6372 14360 6384
rect 13299 6344 14360 6372
rect 13299 6341 13311 6344
rect 13253 6335 13311 6341
rect 14354 6332 14360 6344
rect 14412 6372 14418 6384
rect 14541 6375 14599 6381
rect 14541 6372 14553 6375
rect 14412 6344 14553 6372
rect 14412 6332 14418 6344
rect 14541 6341 14553 6344
rect 14587 6372 14599 6375
rect 15182 6372 15188 6384
rect 14587 6344 15188 6372
rect 14587 6341 14599 6344
rect 14541 6335 14599 6341
rect 15182 6332 15188 6344
rect 15240 6332 15246 6384
rect 20536 6372 20564 6403
rect 20886 6400 20892 6412
rect 20944 6400 20950 6452
rect 21070 6400 21076 6452
rect 21128 6440 21134 6452
rect 22085 6443 22143 6449
rect 22085 6440 22097 6443
rect 21128 6412 22097 6440
rect 21128 6400 21134 6412
rect 22085 6409 22097 6412
rect 22131 6409 22143 6443
rect 22085 6403 22143 6409
rect 23554 6400 23560 6452
rect 23612 6440 23618 6452
rect 23833 6443 23891 6449
rect 23833 6440 23845 6443
rect 23612 6412 23845 6440
rect 23612 6400 23618 6412
rect 23833 6409 23845 6412
rect 23879 6409 23891 6443
rect 24750 6440 24756 6452
rect 24711 6412 24756 6440
rect 23833 6403 23891 6409
rect 24750 6400 24756 6412
rect 24808 6400 24814 6452
rect 20794 6372 20800 6384
rect 20536 6344 20800 6372
rect 20794 6332 20800 6344
rect 20852 6332 20858 6384
rect 15366 6304 15372 6316
rect 15327 6276 15372 6304
rect 15366 6264 15372 6276
rect 15424 6264 15430 6316
rect 17482 6264 17488 6316
rect 17540 6304 17546 6316
rect 17577 6307 17635 6313
rect 17577 6304 17589 6307
rect 17540 6276 17589 6304
rect 17540 6264 17546 6276
rect 17577 6273 17589 6276
rect 17623 6273 17635 6307
rect 17577 6267 17635 6273
rect 19046 6264 19052 6316
rect 19104 6304 19110 6316
rect 19325 6307 19383 6313
rect 19325 6304 19337 6307
rect 19104 6276 19337 6304
rect 19104 6264 19110 6276
rect 19325 6273 19337 6276
rect 19371 6273 19383 6307
rect 19325 6267 19383 6273
rect 11321 6239 11379 6245
rect 11321 6205 11333 6239
rect 11367 6236 11379 6239
rect 11870 6236 11876 6248
rect 11367 6208 11876 6236
rect 11367 6205 11379 6208
rect 11321 6199 11379 6205
rect 11870 6196 11876 6208
rect 11928 6236 11934 6248
rect 12057 6239 12115 6245
rect 12057 6236 12069 6239
rect 11928 6208 12069 6236
rect 11928 6196 11934 6208
rect 12057 6205 12069 6208
rect 12103 6205 12115 6239
rect 12057 6199 12115 6205
rect 15690 6171 15748 6177
rect 15690 6168 15702 6171
rect 15200 6140 15702 6168
rect 11594 6100 11600 6112
rect 11555 6072 11600 6100
rect 11594 6060 11600 6072
rect 11652 6060 11658 6112
rect 15090 6060 15096 6112
rect 15148 6100 15154 6112
rect 15200 6109 15228 6140
rect 15690 6137 15702 6140
rect 15736 6168 15748 6171
rect 17393 6171 17451 6177
rect 17393 6168 17405 6171
rect 15736 6140 17405 6168
rect 15736 6137 15748 6140
rect 15690 6131 15748 6137
rect 17393 6137 17405 6140
rect 17439 6168 17451 6171
rect 17758 6168 17764 6180
rect 17439 6140 17764 6168
rect 17439 6137 17451 6140
rect 17393 6131 17451 6137
rect 17758 6128 17764 6140
rect 17816 6168 17822 6180
rect 19690 6177 19696 6180
rect 17939 6171 17997 6177
rect 17939 6168 17951 6171
rect 17816 6140 17951 6168
rect 17816 6128 17822 6140
rect 17939 6137 17951 6140
rect 17985 6168 17997 6171
rect 19233 6171 19291 6177
rect 19233 6168 19245 6171
rect 17985 6140 19245 6168
rect 17985 6137 17997 6140
rect 17939 6131 17997 6137
rect 19233 6137 19245 6140
rect 19279 6168 19291 6171
rect 19687 6168 19696 6177
rect 19279 6140 19696 6168
rect 19279 6137 19291 6140
rect 19233 6131 19291 6137
rect 19687 6131 19696 6140
rect 19690 6128 19696 6131
rect 19748 6128 19754 6180
rect 15185 6103 15243 6109
rect 15185 6100 15197 6103
rect 15148 6072 15197 6100
rect 15148 6060 15154 6072
rect 15185 6069 15197 6072
rect 15231 6069 15243 6103
rect 16286 6100 16292 6112
rect 16247 6072 16292 6100
rect 15185 6063 15243 6069
rect 16286 6060 16292 6072
rect 16344 6060 16350 6112
rect 20242 6100 20248 6112
rect 20203 6072 20248 6100
rect 20242 6060 20248 6072
rect 20300 6060 20306 6112
rect 20904 6100 20932 6400
rect 23327 6375 23385 6381
rect 23327 6341 23339 6375
rect 23373 6372 23385 6375
rect 24198 6372 24204 6384
rect 23373 6344 24204 6372
rect 23373 6341 23385 6344
rect 23327 6335 23385 6341
rect 24198 6332 24204 6344
rect 24256 6332 24262 6384
rect 20978 6264 20984 6316
rect 21036 6304 21042 6316
rect 21165 6307 21223 6313
rect 21165 6304 21177 6307
rect 21036 6276 21177 6304
rect 21036 6264 21042 6276
rect 21165 6273 21177 6276
rect 21211 6273 21223 6307
rect 21438 6304 21444 6316
rect 21399 6276 21444 6304
rect 21165 6267 21223 6273
rect 21438 6264 21444 6276
rect 21496 6304 21502 6316
rect 22913 6307 22971 6313
rect 22913 6304 22925 6307
rect 21496 6276 22925 6304
rect 21496 6264 21502 6276
rect 22913 6273 22925 6276
rect 22959 6273 22971 6307
rect 22913 6267 22971 6273
rect 22928 6236 22956 6267
rect 23002 6264 23008 6316
rect 23060 6304 23066 6316
rect 24339 6307 24397 6313
rect 24339 6304 24351 6307
rect 23060 6276 24351 6304
rect 23060 6264 23066 6276
rect 24339 6273 24351 6276
rect 24385 6273 24397 6307
rect 24339 6267 24397 6273
rect 23224 6239 23282 6245
rect 23224 6236 23236 6239
rect 22928 6208 23236 6236
rect 23224 6205 23236 6208
rect 23270 6205 23282 6239
rect 23224 6199 23282 6205
rect 24252 6239 24310 6245
rect 24252 6205 24264 6239
rect 24298 6236 24310 6239
rect 24750 6236 24756 6248
rect 24298 6208 24756 6236
rect 24298 6205 24310 6208
rect 24252 6199 24310 6205
rect 24750 6196 24756 6208
rect 24808 6196 24814 6248
rect 21257 6171 21315 6177
rect 21257 6137 21269 6171
rect 21303 6137 21315 6171
rect 21257 6131 21315 6137
rect 21272 6100 21300 6131
rect 25118 6100 25124 6112
rect 20904 6072 21300 6100
rect 25079 6072 25124 6100
rect 25118 6060 25124 6072
rect 25176 6060 25182 6112
rect 632 6010 26392 6032
rect 632 5958 9843 6010
rect 9895 5958 9907 6010
rect 9959 5958 9971 6010
rect 10023 5958 10035 6010
rect 10087 5958 19176 6010
rect 19228 5958 19240 6010
rect 19292 5958 19304 6010
rect 19356 5958 19368 6010
rect 19420 5958 26392 6010
rect 632 5936 26392 5958
rect 17482 5856 17488 5908
rect 17540 5896 17546 5908
rect 17577 5899 17635 5905
rect 17577 5896 17589 5899
rect 17540 5868 17589 5896
rect 17540 5856 17546 5868
rect 17577 5865 17589 5868
rect 17623 5865 17635 5899
rect 17577 5859 17635 5865
rect 19046 5856 19052 5908
rect 19104 5896 19110 5908
rect 19325 5899 19383 5905
rect 19325 5896 19337 5899
rect 19104 5868 19337 5896
rect 19104 5856 19110 5868
rect 19325 5865 19337 5868
rect 19371 5865 19383 5899
rect 19325 5859 19383 5865
rect 20242 5856 20248 5908
rect 20300 5896 20306 5908
rect 21070 5896 21076 5908
rect 20300 5868 21076 5896
rect 20300 5856 20306 5868
rect 15090 5788 15096 5840
rect 15148 5837 15154 5840
rect 15148 5831 15196 5837
rect 15148 5797 15150 5831
rect 15184 5797 15196 5831
rect 15148 5791 15196 5797
rect 15148 5788 15154 5791
rect 16286 5788 16292 5840
rect 16344 5828 16350 5840
rect 16749 5831 16807 5837
rect 16749 5828 16761 5831
rect 16344 5800 16761 5828
rect 16344 5788 16350 5800
rect 16749 5797 16761 5800
rect 16795 5828 16807 5831
rect 16930 5828 16936 5840
rect 16795 5800 16936 5828
rect 16795 5797 16807 5800
rect 16749 5791 16807 5797
rect 16930 5788 16936 5800
rect 16988 5828 16994 5840
rect 20628 5837 20656 5868
rect 21070 5856 21076 5868
rect 21128 5856 21134 5908
rect 23235 5899 23293 5905
rect 23235 5865 23247 5899
rect 23281 5896 23293 5899
rect 24290 5896 24296 5908
rect 23281 5868 24296 5896
rect 23281 5865 23293 5868
rect 23235 5859 23293 5865
rect 24290 5856 24296 5868
rect 24348 5856 24354 5908
rect 20613 5831 20671 5837
rect 16988 5800 18264 5828
rect 16988 5788 16994 5800
rect 13894 5720 13900 5772
rect 13952 5760 13958 5772
rect 14817 5763 14875 5769
rect 14817 5760 14829 5763
rect 13952 5732 14829 5760
rect 13952 5720 13958 5732
rect 14817 5729 14829 5732
rect 14863 5760 14875 5763
rect 14998 5760 15004 5772
rect 14863 5732 15004 5760
rect 14863 5729 14875 5732
rect 14817 5723 14875 5729
rect 14998 5720 15004 5732
rect 15056 5720 15062 5772
rect 18236 5769 18264 5800
rect 20613 5797 20625 5831
rect 20659 5797 20671 5831
rect 20613 5791 20671 5797
rect 21165 5831 21223 5837
rect 21165 5797 21177 5831
rect 21211 5828 21223 5831
rect 21438 5828 21444 5840
rect 21211 5800 21444 5828
rect 21211 5797 21223 5800
rect 21165 5791 21223 5797
rect 21438 5788 21444 5800
rect 21496 5788 21502 5840
rect 18221 5763 18279 5769
rect 18221 5729 18233 5763
rect 18267 5760 18279 5763
rect 18586 5760 18592 5772
rect 18267 5732 18592 5760
rect 18267 5729 18279 5732
rect 18221 5723 18279 5729
rect 18586 5720 18592 5732
rect 18644 5720 18650 5772
rect 23094 5720 23100 5772
rect 23152 5769 23158 5772
rect 23152 5763 23190 5769
rect 23178 5729 23190 5763
rect 23152 5723 23190 5729
rect 24176 5763 24234 5769
rect 24176 5729 24188 5763
rect 24222 5760 24234 5763
rect 25026 5760 25032 5772
rect 24222 5732 25032 5760
rect 24222 5729 24234 5732
rect 24176 5723 24234 5729
rect 23152 5720 23158 5723
rect 25026 5720 25032 5732
rect 25084 5720 25090 5772
rect 16654 5692 16660 5704
rect 16615 5664 16660 5692
rect 16654 5652 16660 5664
rect 16712 5652 16718 5704
rect 17301 5695 17359 5701
rect 17301 5661 17313 5695
rect 17347 5692 17359 5695
rect 17390 5692 17396 5704
rect 17347 5664 17396 5692
rect 17347 5661 17359 5664
rect 17301 5655 17359 5661
rect 17390 5652 17396 5664
rect 17448 5652 17454 5704
rect 18126 5692 18132 5704
rect 18087 5664 18132 5692
rect 18126 5652 18132 5664
rect 18184 5652 18190 5704
rect 19874 5652 19880 5704
rect 19932 5692 19938 5704
rect 20521 5695 20579 5701
rect 20521 5692 20533 5695
rect 19932 5664 20533 5692
rect 19932 5652 19938 5664
rect 20521 5661 20533 5664
rect 20567 5661 20579 5695
rect 20521 5655 20579 5661
rect 10582 5584 10588 5636
rect 10640 5624 10646 5636
rect 11870 5624 11876 5636
rect 10640 5596 11876 5624
rect 10640 5584 10646 5596
rect 11870 5584 11876 5596
rect 11928 5624 11934 5636
rect 11965 5627 12023 5633
rect 11965 5624 11977 5627
rect 11928 5596 11977 5624
rect 11928 5584 11934 5596
rect 11965 5593 11977 5596
rect 12011 5593 12023 5627
rect 11965 5587 12023 5593
rect 23646 5584 23652 5636
rect 23704 5624 23710 5636
rect 24247 5627 24305 5633
rect 24247 5624 24259 5627
rect 23704 5596 24259 5624
rect 23704 5584 23710 5596
rect 24247 5593 24259 5596
rect 24293 5593 24305 5627
rect 24247 5587 24305 5593
rect 15734 5556 15740 5568
rect 15695 5528 15740 5556
rect 15734 5516 15740 5528
rect 15792 5516 15798 5568
rect 632 5466 26392 5488
rect 632 5414 5176 5466
rect 5228 5414 5240 5466
rect 5292 5414 5304 5466
rect 5356 5414 5368 5466
rect 5420 5414 14510 5466
rect 14562 5414 14574 5466
rect 14626 5414 14638 5466
rect 14690 5414 14702 5466
rect 14754 5414 23843 5466
rect 23895 5414 23907 5466
rect 23959 5414 23971 5466
rect 24023 5414 24035 5466
rect 24087 5414 26392 5466
rect 632 5392 26392 5414
rect 13986 5352 13992 5364
rect 13947 5324 13992 5352
rect 13986 5312 13992 5324
rect 14044 5312 14050 5364
rect 14817 5355 14875 5361
rect 14817 5321 14829 5355
rect 14863 5352 14875 5355
rect 15090 5352 15096 5364
rect 14863 5324 15096 5352
rect 14863 5321 14875 5324
rect 14817 5315 14875 5321
rect 15090 5312 15096 5324
rect 15148 5312 15154 5364
rect 16381 5355 16439 5361
rect 16381 5352 16393 5355
rect 15476 5324 16393 5352
rect 14004 5216 14032 5312
rect 15476 5225 15504 5324
rect 16381 5321 16393 5324
rect 16427 5352 16439 5355
rect 16654 5352 16660 5364
rect 16427 5324 16660 5352
rect 16427 5321 16439 5324
rect 16381 5315 16439 5321
rect 16654 5312 16660 5324
rect 16712 5312 16718 5364
rect 16930 5352 16936 5364
rect 16891 5324 16936 5352
rect 16930 5312 16936 5324
rect 16988 5312 16994 5364
rect 18586 5352 18592 5364
rect 18547 5324 18592 5352
rect 18586 5312 18592 5324
rect 18644 5312 18650 5364
rect 20242 5312 20248 5364
rect 20300 5352 20306 5364
rect 20521 5355 20579 5361
rect 20521 5352 20533 5355
rect 20300 5324 20533 5352
rect 20300 5312 20306 5324
rect 20521 5321 20533 5324
rect 20567 5321 20579 5355
rect 20521 5315 20579 5321
rect 23094 5312 23100 5364
rect 23152 5352 23158 5364
rect 23373 5355 23431 5361
rect 23373 5352 23385 5355
rect 23152 5324 23385 5352
rect 23152 5312 23158 5324
rect 23373 5321 23385 5324
rect 23419 5321 23431 5355
rect 23373 5315 23431 5321
rect 23738 5312 23744 5364
rect 23796 5352 23802 5364
rect 24247 5355 24305 5361
rect 24247 5352 24259 5355
rect 23796 5324 24259 5352
rect 23796 5312 23802 5324
rect 24247 5321 24259 5324
rect 24293 5321 24305 5355
rect 24658 5352 24664 5364
rect 24619 5324 24664 5352
rect 24247 5315 24305 5321
rect 24658 5312 24664 5324
rect 24716 5312 24722 5364
rect 25026 5352 25032 5364
rect 24987 5324 25032 5352
rect 25026 5312 25032 5324
rect 25084 5312 25090 5364
rect 15001 5219 15059 5225
rect 15001 5216 15013 5219
rect 14004 5188 15013 5216
rect 15001 5185 15013 5188
rect 15047 5185 15059 5219
rect 15001 5179 15059 5185
rect 15461 5219 15519 5225
rect 15461 5185 15473 5219
rect 15507 5185 15519 5219
rect 15461 5179 15519 5185
rect 17482 5176 17488 5228
rect 17540 5216 17546 5228
rect 17945 5219 18003 5225
rect 17945 5216 17957 5219
rect 17540 5188 17957 5216
rect 17540 5176 17546 5188
rect 17945 5185 17957 5188
rect 17991 5185 18003 5219
rect 19874 5216 19880 5228
rect 19835 5188 19880 5216
rect 17945 5179 18003 5185
rect 19874 5176 19880 5188
rect 19932 5216 19938 5228
rect 20889 5219 20947 5225
rect 20889 5216 20901 5219
rect 19932 5188 20901 5216
rect 19932 5176 19938 5188
rect 20889 5185 20901 5188
rect 20935 5185 20947 5219
rect 20889 5179 20947 5185
rect 24176 5151 24234 5157
rect 24176 5117 24188 5151
rect 24222 5148 24234 5151
rect 24658 5148 24664 5160
rect 24222 5120 24664 5148
rect 24222 5117 24234 5120
rect 24176 5111 24234 5117
rect 24658 5108 24664 5120
rect 24716 5108 24722 5160
rect 14449 5083 14507 5089
rect 14449 5049 14461 5083
rect 14495 5080 14507 5083
rect 15093 5083 15151 5089
rect 14495 5052 14952 5080
rect 14495 5049 14507 5052
rect 14449 5043 14507 5049
rect 14924 5024 14952 5052
rect 15093 5049 15105 5083
rect 15139 5080 15151 5083
rect 15734 5080 15740 5092
rect 15139 5052 15740 5080
rect 15139 5049 15151 5052
rect 15093 5043 15151 5049
rect 14906 5012 14912 5024
rect 14819 4984 14912 5012
rect 14906 4972 14912 4984
rect 14964 5012 14970 5024
rect 15108 5012 15136 5043
rect 15734 5040 15740 5052
rect 15792 5040 15798 5092
rect 16473 5083 16531 5089
rect 16473 5049 16485 5083
rect 16519 5080 16531 5083
rect 17666 5080 17672 5092
rect 16519 5052 17672 5080
rect 16519 5049 16531 5052
rect 16473 5043 16531 5049
rect 17666 5040 17672 5052
rect 17724 5040 17730 5092
rect 17761 5083 17819 5089
rect 17761 5049 17773 5083
rect 17807 5080 17819 5083
rect 18126 5080 18132 5092
rect 17807 5052 18132 5080
rect 17807 5049 17819 5052
rect 17761 5043 17819 5049
rect 14964 4984 15136 5012
rect 17393 5015 17451 5021
rect 14964 4972 14970 4984
rect 17393 4981 17405 5015
rect 17439 5012 17451 5015
rect 17776 5012 17804 5043
rect 18126 5040 18132 5052
rect 18184 5040 18190 5092
rect 19049 5083 19107 5089
rect 19049 5049 19061 5083
rect 19095 5080 19107 5083
rect 19598 5080 19604 5092
rect 19095 5052 19604 5080
rect 19095 5049 19107 5052
rect 19049 5043 19107 5049
rect 19598 5040 19604 5052
rect 19656 5040 19662 5092
rect 19693 5083 19751 5089
rect 19693 5049 19705 5083
rect 19739 5049 19751 5083
rect 19693 5043 19751 5049
rect 17439 4984 17804 5012
rect 19417 5015 19475 5021
rect 17439 4981 17451 4984
rect 17393 4975 17451 4981
rect 19417 4981 19429 5015
rect 19463 5012 19475 5015
rect 19506 5012 19512 5024
rect 19463 4984 19512 5012
rect 19463 4981 19475 4984
rect 19417 4975 19475 4981
rect 19506 4972 19512 4984
rect 19564 5012 19570 5024
rect 19708 5012 19736 5043
rect 19564 4984 19736 5012
rect 19564 4972 19570 4984
rect 632 4922 26392 4944
rect 632 4870 9843 4922
rect 9895 4870 9907 4922
rect 9959 4870 9971 4922
rect 10023 4870 10035 4922
rect 10087 4870 19176 4922
rect 19228 4870 19240 4922
rect 19292 4870 19304 4922
rect 19356 4870 19368 4922
rect 19420 4870 26392 4922
rect 632 4848 26392 4870
rect 14998 4808 15004 4820
rect 14959 4780 15004 4808
rect 14998 4768 15004 4780
rect 15056 4768 15062 4820
rect 17666 4808 17672 4820
rect 17627 4780 17672 4808
rect 17666 4768 17672 4780
rect 17724 4768 17730 4820
rect 23186 4768 23192 4820
rect 23244 4808 23250 4820
rect 24247 4811 24305 4817
rect 24247 4808 24259 4811
rect 23244 4780 24259 4808
rect 23244 4768 23250 4780
rect 24247 4777 24259 4780
rect 24293 4777 24305 4811
rect 24247 4771 24305 4777
rect 15918 4740 15924 4752
rect 15879 4712 15924 4740
rect 15918 4700 15924 4712
rect 15976 4700 15982 4752
rect 16473 4743 16531 4749
rect 16473 4709 16485 4743
rect 16519 4740 16531 4743
rect 16654 4740 16660 4752
rect 16519 4712 16660 4740
rect 16519 4709 16531 4712
rect 16473 4703 16531 4709
rect 16654 4700 16660 4712
rect 16712 4700 16718 4752
rect 19506 4740 19512 4752
rect 19467 4712 19512 4740
rect 19506 4700 19512 4712
rect 19564 4700 19570 4752
rect 18862 4672 18868 4684
rect 18823 4644 18868 4672
rect 18862 4632 18868 4644
rect 18920 4632 18926 4684
rect 24198 4681 24204 4684
rect 24176 4675 24204 4681
rect 24176 4641 24188 4675
rect 24176 4635 24204 4641
rect 24198 4632 24204 4635
rect 24256 4632 24262 4684
rect 15829 4607 15887 4613
rect 15829 4573 15841 4607
rect 15875 4604 15887 4607
rect 16194 4604 16200 4616
rect 15875 4576 16200 4604
rect 15875 4573 15887 4576
rect 15829 4567 15887 4573
rect 16194 4564 16200 4576
rect 16252 4564 16258 4616
rect 632 4378 26392 4400
rect 632 4326 5176 4378
rect 5228 4326 5240 4378
rect 5292 4326 5304 4378
rect 5356 4326 5368 4378
rect 5420 4326 14510 4378
rect 14562 4326 14574 4378
rect 14626 4326 14638 4378
rect 14690 4326 14702 4378
rect 14754 4326 23843 4378
rect 23895 4326 23907 4378
rect 23959 4326 23971 4378
rect 24023 4326 24035 4378
rect 24087 4326 26392 4378
rect 632 4304 26392 4326
rect 14906 4264 14912 4276
rect 14867 4236 14912 4264
rect 14906 4224 14912 4236
rect 14964 4224 14970 4276
rect 18862 4264 18868 4276
rect 18823 4236 18868 4264
rect 18862 4224 18868 4236
rect 18920 4224 18926 4276
rect 15829 4131 15887 4137
rect 15829 4097 15841 4131
rect 15875 4128 15887 4131
rect 15918 4128 15924 4140
rect 15875 4100 15924 4128
rect 15875 4097 15887 4100
rect 15829 4091 15887 4097
rect 15918 4088 15924 4100
rect 15976 4128 15982 4140
rect 16105 4131 16163 4137
rect 16105 4128 16117 4131
rect 15976 4100 16117 4128
rect 15976 4088 15982 4100
rect 16105 4097 16117 4100
rect 16151 4097 16163 4131
rect 16105 4091 16163 4097
rect 16194 4088 16200 4140
rect 16252 4128 16258 4140
rect 16473 4131 16531 4137
rect 16473 4128 16485 4131
rect 16252 4100 16485 4128
rect 16252 4088 16258 4100
rect 16473 4097 16485 4100
rect 16519 4097 16531 4131
rect 25026 4128 25032 4140
rect 24987 4100 25032 4128
rect 16473 4091 16531 4097
rect 25026 4088 25032 4100
rect 25084 4088 25090 4140
rect 14906 4020 14912 4072
rect 14964 4060 14970 4072
rect 15185 4063 15243 4069
rect 15185 4060 15197 4063
rect 14964 4032 15197 4060
rect 14964 4020 14970 4032
rect 15185 4029 15197 4032
rect 15231 4029 15243 4063
rect 15185 4023 15243 4029
rect 24160 4063 24218 4069
rect 24160 4029 24172 4063
rect 24206 4060 24218 4063
rect 24206 4032 24704 4060
rect 24206 4029 24218 4032
rect 24160 4023 24218 4029
rect 23002 3952 23008 4004
rect 23060 3992 23066 4004
rect 24247 3995 24305 4001
rect 24247 3992 24259 3995
rect 23060 3964 24259 3992
rect 23060 3952 23066 3964
rect 24247 3961 24259 3964
rect 24293 3961 24305 3995
rect 24247 3955 24305 3961
rect 24676 3936 24704 4032
rect 24658 3924 24664 3936
rect 24619 3896 24664 3924
rect 24658 3884 24664 3896
rect 24716 3884 24722 3936
rect 632 3834 26392 3856
rect 632 3782 9843 3834
rect 9895 3782 9907 3834
rect 9959 3782 9971 3834
rect 10023 3782 10035 3834
rect 10087 3782 19176 3834
rect 19228 3782 19240 3834
rect 19292 3782 19304 3834
rect 19356 3782 19368 3834
rect 19420 3782 26392 3834
rect 632 3760 26392 3782
rect 16194 3680 16200 3732
rect 16252 3720 16258 3732
rect 16335 3723 16393 3729
rect 16335 3720 16347 3723
rect 16252 3692 16347 3720
rect 16252 3680 16258 3692
rect 16335 3689 16347 3692
rect 16381 3689 16393 3723
rect 16335 3683 16393 3689
rect 16286 3593 16292 3596
rect 16264 3587 16292 3593
rect 16264 3553 16276 3587
rect 16264 3547 16292 3553
rect 16286 3544 16292 3547
rect 16344 3544 16350 3596
rect 632 3290 26392 3312
rect 632 3238 5176 3290
rect 5228 3238 5240 3290
rect 5292 3238 5304 3290
rect 5356 3238 5368 3290
rect 5420 3238 14510 3290
rect 14562 3238 14574 3290
rect 14626 3238 14638 3290
rect 14690 3238 14702 3290
rect 14754 3238 23843 3290
rect 23895 3238 23907 3290
rect 23959 3238 23971 3290
rect 24023 3238 24035 3290
rect 24087 3238 26392 3290
rect 632 3216 26392 3238
rect 16286 2972 16292 2984
rect 16247 2944 16292 2972
rect 16286 2932 16292 2944
rect 16344 2932 16350 2984
rect 632 2746 26392 2768
rect 632 2694 9843 2746
rect 9895 2694 9907 2746
rect 9959 2694 9971 2746
rect 10023 2694 10035 2746
rect 10087 2694 19176 2746
rect 19228 2694 19240 2746
rect 19292 2694 19304 2746
rect 19356 2694 19368 2746
rect 19420 2694 26392 2746
rect 632 2672 26392 2694
rect 23462 2592 23468 2644
rect 23520 2632 23526 2644
rect 24247 2635 24305 2641
rect 24247 2632 24259 2635
rect 23520 2604 24259 2632
rect 23520 2592 23526 2604
rect 24247 2601 24259 2604
rect 24293 2601 24305 2635
rect 24247 2595 24305 2601
rect 24176 2499 24234 2505
rect 24176 2465 24188 2499
rect 24222 2496 24234 2499
rect 24658 2496 24664 2508
rect 24222 2468 24664 2496
rect 24222 2465 24234 2468
rect 24176 2459 24234 2465
rect 24658 2456 24664 2468
rect 24716 2456 24722 2508
rect 24658 2292 24664 2304
rect 24619 2264 24664 2292
rect 24658 2252 24664 2264
rect 24716 2252 24722 2304
rect 632 2202 26392 2224
rect 632 2150 5176 2202
rect 5228 2150 5240 2202
rect 5292 2150 5304 2202
rect 5356 2150 5368 2202
rect 5420 2150 14510 2202
rect 14562 2150 14574 2202
rect 14626 2150 14638 2202
rect 14690 2150 14702 2202
rect 14754 2150 23843 2202
rect 23895 2150 23907 2202
rect 23959 2150 23971 2202
rect 24023 2150 24035 2202
rect 24087 2150 26392 2202
rect 632 2128 26392 2150
<< via1 >>
rect 9843 25542 9895 25594
rect 9907 25542 9959 25594
rect 9971 25542 10023 25594
rect 10035 25542 10087 25594
rect 19176 25542 19228 25594
rect 19240 25542 19292 25594
rect 19304 25542 19356 25594
rect 19368 25542 19420 25594
rect 13256 25304 13308 25356
rect 20800 25347 20852 25356
rect 20800 25313 20818 25347
rect 20818 25313 20852 25347
rect 20800 25304 20852 25313
rect 17120 25100 17172 25152
rect 21996 25100 22048 25152
rect 5176 24998 5228 25050
rect 5240 24998 5292 25050
rect 5304 24998 5356 25050
rect 5368 24998 5420 25050
rect 14510 24998 14562 25050
rect 14574 24998 14626 25050
rect 14638 24998 14690 25050
rect 14702 24998 14754 25050
rect 23843 24998 23895 25050
rect 23907 24998 23959 25050
rect 23971 24998 24023 25050
rect 24035 24998 24087 25050
rect 13256 24896 13308 24948
rect 20800 24939 20852 24948
rect 20800 24905 20809 24939
rect 20809 24905 20843 24939
rect 20843 24905 20852 24939
rect 20800 24896 20852 24905
rect 11324 24803 11376 24812
rect 11324 24769 11333 24803
rect 11333 24769 11367 24803
rect 11367 24769 11376 24803
rect 11324 24760 11376 24769
rect 24296 24803 24348 24812
rect 24296 24769 24305 24803
rect 24305 24769 24339 24803
rect 24339 24769 24348 24803
rect 24296 24760 24348 24769
rect 25400 24803 25452 24812
rect 25400 24769 25409 24803
rect 25409 24769 25443 24803
rect 25443 24769 25452 24803
rect 25400 24760 25452 24769
rect 12612 24735 12664 24744
rect 12612 24701 12656 24735
rect 12656 24701 12664 24735
rect 12612 24692 12664 24701
rect 14084 24692 14136 24744
rect 15464 24735 15516 24744
rect 15464 24701 15482 24735
rect 15482 24701 15516 24735
rect 15464 24692 15516 24701
rect 20156 24735 20208 24744
rect 20156 24701 20165 24735
rect 20165 24701 20199 24735
rect 20199 24701 20208 24735
rect 20156 24692 20208 24701
rect 21352 24692 21404 24744
rect 14176 24624 14228 24676
rect 20524 24667 20576 24676
rect 20524 24633 20533 24667
rect 20533 24633 20567 24667
rect 20567 24633 20576 24667
rect 20524 24624 20576 24633
rect 11048 24556 11100 24608
rect 14452 24599 14504 24608
rect 14452 24565 14461 24599
rect 14461 24565 14495 24599
rect 14495 24565 14504 24599
rect 14452 24556 14504 24565
rect 16016 24556 16068 24608
rect 18040 24556 18092 24608
rect 21812 24556 21864 24608
rect 24204 24556 24256 24608
rect 25032 24556 25084 24608
rect 9843 24454 9895 24506
rect 9907 24454 9959 24506
rect 9971 24454 10023 24506
rect 10035 24454 10087 24506
rect 19176 24454 19228 24506
rect 19240 24454 19292 24506
rect 19304 24454 19356 24506
rect 19368 24454 19420 24506
rect 15004 24395 15056 24404
rect 15004 24361 15013 24395
rect 15013 24361 15047 24395
rect 15047 24361 15056 24395
rect 15004 24352 15056 24361
rect 18500 24395 18552 24404
rect 18500 24361 18509 24395
rect 18509 24361 18543 24395
rect 18543 24361 18552 24395
rect 18500 24352 18552 24361
rect 22272 24395 22324 24404
rect 22272 24361 22281 24395
rect 22281 24361 22315 24395
rect 22315 24361 22324 24395
rect 22272 24352 22324 24361
rect 24848 24352 24900 24404
rect 20524 24284 20576 24336
rect 6172 24216 6224 24268
rect 8288 24216 8340 24268
rect 9300 24259 9352 24268
rect 9300 24225 9318 24259
rect 9318 24225 9352 24259
rect 9300 24216 9352 24225
rect 12888 24216 12940 24268
rect 13808 24259 13860 24268
rect 13808 24225 13826 24259
rect 13826 24225 13860 24259
rect 13808 24216 13860 24225
rect 14360 24216 14412 24268
rect 11692 24148 11744 24200
rect 12152 24191 12204 24200
rect 12152 24157 12161 24191
rect 12161 24157 12195 24191
rect 12195 24157 12204 24191
rect 12152 24148 12204 24157
rect 14176 24148 14228 24200
rect 16752 24216 16804 24268
rect 18316 24259 18368 24268
rect 18316 24225 18325 24259
rect 18325 24225 18359 24259
rect 18359 24225 18368 24259
rect 18316 24216 18368 24225
rect 21812 24216 21864 24268
rect 22640 24216 22692 24268
rect 24296 24216 24348 24268
rect 24572 24259 24624 24268
rect 24572 24225 24590 24259
rect 24590 24225 24624 24259
rect 24572 24216 24624 24225
rect 20616 24148 20668 24200
rect 24480 24080 24532 24132
rect 6264 24012 6316 24064
rect 8196 24012 8248 24064
rect 9392 24012 9444 24064
rect 14268 24012 14320 24064
rect 17212 24055 17264 24064
rect 17212 24021 17221 24055
rect 17221 24021 17255 24055
rect 17255 24021 17264 24055
rect 17212 24012 17264 24021
rect 17764 24055 17816 24064
rect 17764 24021 17773 24055
rect 17773 24021 17807 24055
rect 17807 24021 17816 24055
rect 17764 24012 17816 24021
rect 20800 24012 20852 24064
rect 5176 23910 5228 23962
rect 5240 23910 5292 23962
rect 5304 23910 5356 23962
rect 5368 23910 5420 23962
rect 14510 23910 14562 23962
rect 14574 23910 14626 23962
rect 14638 23910 14690 23962
rect 14702 23910 14754 23962
rect 23843 23910 23895 23962
rect 23907 23910 23959 23962
rect 23971 23910 24023 23962
rect 24035 23910 24087 23962
rect 1940 23808 1992 23860
rect 2032 23808 2084 23860
rect 3044 23808 3096 23860
rect 5068 23808 5120 23860
rect 6172 23808 6224 23860
rect 7184 23808 7236 23860
rect 8380 23851 8432 23860
rect 8380 23817 8389 23851
rect 8389 23817 8423 23851
rect 8423 23817 8432 23851
rect 8380 23808 8432 23817
rect 9300 23851 9352 23860
rect 9300 23817 9309 23851
rect 9309 23817 9343 23851
rect 9343 23817 9352 23851
rect 9300 23808 9352 23817
rect 10312 23851 10364 23860
rect 10312 23817 10321 23851
rect 10321 23817 10355 23851
rect 10355 23817 10364 23851
rect 10312 23808 10364 23817
rect 10956 23851 11008 23860
rect 10956 23817 10965 23851
rect 10965 23817 10999 23851
rect 10999 23817 11008 23851
rect 10956 23808 11008 23817
rect 11692 23851 11744 23860
rect 11692 23817 11701 23851
rect 11701 23817 11735 23851
rect 11735 23817 11744 23851
rect 11692 23808 11744 23817
rect 12152 23851 12204 23860
rect 12152 23817 12161 23851
rect 12161 23817 12195 23851
rect 12195 23817 12204 23851
rect 12152 23808 12204 23817
rect 13808 23851 13860 23860
rect 13808 23817 13817 23851
rect 13817 23817 13851 23851
rect 13851 23817 13860 23851
rect 13808 23808 13860 23817
rect 14084 23808 14136 23860
rect 14176 23808 14228 23860
rect 19696 23851 19748 23860
rect 19696 23817 19705 23851
rect 19705 23817 19739 23851
rect 19739 23817 19748 23851
rect 19696 23808 19748 23817
rect 20524 23851 20576 23860
rect 20524 23817 20533 23851
rect 20533 23817 20567 23851
rect 20567 23817 20576 23851
rect 20524 23808 20576 23817
rect 21812 23808 21864 23860
rect 22640 23851 22692 23860
rect 22640 23817 22649 23851
rect 22649 23817 22683 23851
rect 22683 23817 22692 23851
rect 22640 23808 22692 23817
rect 24572 23851 24624 23860
rect 24572 23817 24581 23851
rect 24581 23817 24615 23851
rect 24615 23817 24624 23851
rect 24572 23808 24624 23817
rect 25308 23851 25360 23860
rect 25308 23817 25317 23851
rect 25317 23817 25351 23851
rect 25351 23817 25360 23851
rect 25308 23808 25360 23817
rect 8288 23740 8340 23792
rect 18316 23740 18368 23792
rect 20800 23672 20852 23724
rect 2032 23604 2084 23656
rect 3044 23604 3096 23656
rect 5068 23604 5120 23656
rect 7184 23604 7236 23656
rect 8380 23604 8432 23656
rect 10312 23604 10364 23656
rect 10956 23604 11008 23656
rect 12152 23536 12204 23588
rect 13072 23579 13124 23588
rect 13072 23545 13081 23579
rect 13081 23545 13115 23579
rect 13115 23545 13124 23579
rect 13072 23536 13124 23545
rect 15832 23536 15884 23588
rect 23008 23647 23060 23656
rect 17764 23579 17816 23588
rect 17764 23545 17773 23579
rect 17773 23545 17807 23579
rect 17807 23545 17816 23579
rect 17764 23536 17816 23545
rect 3596 23468 3648 23520
rect 4976 23468 5028 23520
rect 7736 23468 7788 23520
rect 8932 23468 8984 23520
rect 10312 23468 10364 23520
rect 15188 23511 15240 23520
rect 15188 23477 15197 23511
rect 15197 23477 15231 23511
rect 15231 23477 15240 23511
rect 15188 23468 15240 23477
rect 16292 23511 16344 23520
rect 16292 23477 16301 23511
rect 16301 23477 16335 23511
rect 16335 23477 16344 23511
rect 16292 23468 16344 23477
rect 16752 23468 16804 23520
rect 17396 23511 17448 23520
rect 17396 23477 17405 23511
rect 17405 23477 17439 23511
rect 17439 23477 17448 23511
rect 18500 23536 18552 23588
rect 23008 23613 23017 23647
rect 23017 23613 23051 23647
rect 23051 23613 23060 23647
rect 23008 23604 23060 23613
rect 25308 23604 25360 23656
rect 21352 23579 21404 23588
rect 17396 23468 17448 23477
rect 19512 23468 19564 23520
rect 20156 23511 20208 23520
rect 20156 23477 20165 23511
rect 20165 23477 20199 23511
rect 20199 23477 20208 23511
rect 21352 23545 21361 23579
rect 21361 23545 21395 23579
rect 21395 23545 21404 23579
rect 21352 23536 21404 23545
rect 23192 23579 23244 23588
rect 23192 23545 23201 23579
rect 23201 23545 23235 23579
rect 23235 23545 23244 23579
rect 23192 23536 23244 23545
rect 20156 23468 20208 23477
rect 24480 23468 24532 23520
rect 9843 23366 9895 23418
rect 9907 23366 9959 23418
rect 9971 23366 10023 23418
rect 10035 23366 10087 23418
rect 19176 23366 19228 23418
rect 19240 23366 19292 23418
rect 19304 23366 19356 23418
rect 19368 23366 19420 23418
rect 20616 23264 20668 23316
rect 22916 23264 22968 23316
rect 10864 23239 10916 23248
rect 10864 23205 10873 23239
rect 10873 23205 10907 23239
rect 10907 23205 10916 23239
rect 10864 23196 10916 23205
rect 11324 23196 11376 23248
rect 12888 23196 12940 23248
rect 13072 23239 13124 23248
rect 13072 23205 13081 23239
rect 13081 23205 13115 23239
rect 13115 23205 13124 23239
rect 13072 23196 13124 23205
rect 15188 23239 15240 23248
rect 15188 23205 15197 23239
rect 15197 23205 15231 23239
rect 15231 23205 15240 23239
rect 15188 23196 15240 23205
rect 16752 23239 16804 23248
rect 16752 23205 16761 23239
rect 16761 23205 16795 23239
rect 16795 23205 16804 23239
rect 16752 23196 16804 23205
rect 18224 23196 18276 23248
rect 21444 23239 21496 23248
rect 21444 23205 21453 23239
rect 21453 23205 21487 23239
rect 21487 23205 21496 23239
rect 21444 23196 21496 23205
rect 21628 23196 21680 23248
rect 24204 23264 24256 23316
rect 24388 23264 24440 23316
rect 23192 23196 23244 23248
rect 9852 23171 9904 23180
rect 9852 23137 9861 23171
rect 9861 23137 9895 23171
rect 9895 23137 9904 23171
rect 9852 23128 9904 23137
rect 24572 23171 24624 23180
rect 24572 23137 24590 23171
rect 24590 23137 24624 23171
rect 24572 23128 24624 23137
rect 9208 23103 9260 23112
rect 9208 23069 9217 23103
rect 9217 23069 9251 23103
rect 9251 23069 9260 23103
rect 9208 23060 9260 23069
rect 12428 23103 12480 23112
rect 12428 23069 12437 23103
rect 12437 23069 12471 23103
rect 12471 23069 12480 23103
rect 12428 23060 12480 23069
rect 15096 23103 15148 23112
rect 15096 23069 15105 23103
rect 15105 23069 15139 23103
rect 15139 23069 15148 23103
rect 15096 23060 15148 23069
rect 15924 23060 15976 23112
rect 16292 23060 16344 23112
rect 16660 23103 16712 23112
rect 16660 23069 16669 23103
rect 16669 23069 16703 23103
rect 16703 23069 16712 23103
rect 16660 23060 16712 23069
rect 17304 23103 17356 23112
rect 17304 23069 17313 23103
rect 17313 23069 17347 23103
rect 17347 23069 17356 23103
rect 17304 23060 17356 23069
rect 17764 23060 17816 23112
rect 18040 23060 18092 23112
rect 18500 23103 18552 23112
rect 18500 23069 18509 23103
rect 18509 23069 18543 23103
rect 18543 23069 18552 23103
rect 18500 23060 18552 23069
rect 23284 23103 23336 23112
rect 23284 23069 23293 23103
rect 23293 23069 23327 23103
rect 23327 23069 23336 23103
rect 23284 23060 23336 23069
rect 17672 23035 17724 23044
rect 17672 23001 17681 23035
rect 17681 23001 17715 23035
rect 17715 23001 17724 23035
rect 17672 22992 17724 23001
rect 15648 22924 15700 22976
rect 20708 22967 20760 22976
rect 20708 22933 20717 22967
rect 20717 22933 20751 22967
rect 20751 22933 20760 22967
rect 20708 22924 20760 22933
rect 5176 22822 5228 22874
rect 5240 22822 5292 22874
rect 5304 22822 5356 22874
rect 5368 22822 5420 22874
rect 14510 22822 14562 22874
rect 14574 22822 14626 22874
rect 14638 22822 14690 22874
rect 14702 22822 14754 22874
rect 23843 22822 23895 22874
rect 23907 22822 23959 22874
rect 23971 22822 24023 22874
rect 24035 22822 24087 22874
rect 9208 22763 9260 22772
rect 9208 22729 9217 22763
rect 9217 22729 9251 22763
rect 9251 22729 9260 22763
rect 9208 22720 9260 22729
rect 9576 22720 9628 22772
rect 9852 22720 9904 22772
rect 10956 22720 11008 22772
rect 11324 22763 11376 22772
rect 11324 22729 11333 22763
rect 11333 22729 11367 22763
rect 11367 22729 11376 22763
rect 11324 22720 11376 22729
rect 15096 22720 15148 22772
rect 16660 22720 16712 22772
rect 17212 22720 17264 22772
rect 18040 22720 18092 22772
rect 19512 22720 19564 22772
rect 21628 22763 21680 22772
rect 21628 22729 21637 22763
rect 21637 22729 21671 22763
rect 21671 22729 21680 22763
rect 21628 22720 21680 22729
rect 23192 22720 23244 22772
rect 24204 22763 24256 22772
rect 24204 22729 24213 22763
rect 24213 22729 24247 22763
rect 24247 22729 24256 22763
rect 24204 22720 24256 22729
rect 21444 22652 21496 22704
rect 12428 22627 12480 22636
rect 12428 22593 12437 22627
rect 12437 22593 12471 22627
rect 12471 22593 12480 22627
rect 12428 22584 12480 22593
rect 14084 22627 14136 22636
rect 14084 22593 14093 22627
rect 14093 22593 14127 22627
rect 14127 22593 14136 22627
rect 14084 22584 14136 22593
rect 15188 22584 15240 22636
rect 15648 22627 15700 22636
rect 9208 22380 9260 22432
rect 10220 22448 10272 22500
rect 15648 22593 15657 22627
rect 15657 22593 15691 22627
rect 15691 22593 15700 22627
rect 15648 22584 15700 22593
rect 15924 22627 15976 22636
rect 15924 22593 15933 22627
rect 15933 22593 15967 22627
rect 15967 22593 15976 22627
rect 15924 22584 15976 22593
rect 17304 22584 17356 22636
rect 21352 22627 21404 22636
rect 21352 22593 21361 22627
rect 21361 22593 21395 22627
rect 21395 22593 21404 22627
rect 21352 22584 21404 22593
rect 23284 22627 23336 22636
rect 23284 22593 23293 22627
rect 23293 22593 23327 22627
rect 23327 22593 23336 22627
rect 23284 22584 23336 22593
rect 23560 22627 23612 22636
rect 23560 22593 23569 22627
rect 23569 22593 23603 22627
rect 23603 22593 23612 22627
rect 24572 22627 24624 22636
rect 23560 22584 23612 22593
rect 24572 22593 24581 22627
rect 24581 22593 24615 22627
rect 24615 22593 24624 22627
rect 24572 22584 24624 22593
rect 18500 22516 18552 22568
rect 12060 22491 12112 22500
rect 12060 22457 12069 22491
rect 12069 22457 12103 22491
rect 12103 22457 12112 22491
rect 12060 22448 12112 22457
rect 11876 22380 11928 22432
rect 12888 22380 12940 22432
rect 13348 22380 13400 22432
rect 15832 22448 15884 22500
rect 17672 22491 17724 22500
rect 17672 22457 17681 22491
rect 17681 22457 17715 22491
rect 17715 22457 17724 22491
rect 17672 22448 17724 22457
rect 20708 22491 20760 22500
rect 16660 22423 16712 22432
rect 16660 22389 16669 22423
rect 16669 22389 16703 22423
rect 16703 22389 16712 22423
rect 16660 22380 16712 22389
rect 17212 22380 17264 22432
rect 20708 22457 20717 22491
rect 20717 22457 20751 22491
rect 20751 22457 20760 22491
rect 20708 22448 20760 22457
rect 18132 22380 18184 22432
rect 20616 22380 20668 22432
rect 23192 22380 23244 22432
rect 9843 22278 9895 22330
rect 9907 22278 9959 22330
rect 9971 22278 10023 22330
rect 10035 22278 10087 22330
rect 19176 22278 19228 22330
rect 19240 22278 19292 22330
rect 19304 22278 19356 22330
rect 19368 22278 19420 22330
rect 10864 22219 10916 22228
rect 10864 22185 10873 22219
rect 10873 22185 10907 22219
rect 10907 22185 10916 22219
rect 10864 22176 10916 22185
rect 11876 22219 11928 22228
rect 11876 22185 11885 22219
rect 11885 22185 11919 22219
rect 11919 22185 11928 22219
rect 11876 22176 11928 22185
rect 14084 22176 14136 22228
rect 20708 22176 20760 22228
rect 23284 22176 23336 22228
rect 9576 22151 9628 22160
rect 9576 22117 9585 22151
rect 9585 22117 9619 22151
rect 9619 22117 9628 22151
rect 9576 22108 9628 22117
rect 10220 22108 10272 22160
rect 1020 22083 1072 22092
rect 1020 22049 1038 22083
rect 1038 22049 1072 22083
rect 1020 22040 1072 22049
rect 11324 22040 11376 22092
rect 13256 22040 13308 22092
rect 13808 22083 13860 22092
rect 13808 22049 13817 22083
rect 13817 22049 13851 22083
rect 13851 22049 13860 22083
rect 13808 22040 13860 22049
rect 14912 22108 14964 22160
rect 15648 22108 15700 22160
rect 18132 22151 18184 22160
rect 18132 22117 18141 22151
rect 18141 22117 18175 22151
rect 18175 22117 18184 22151
rect 18132 22108 18184 22117
rect 20248 22108 20300 22160
rect 23008 22151 23060 22160
rect 23008 22117 23017 22151
rect 23017 22117 23051 22151
rect 23051 22117 23060 22151
rect 23008 22108 23060 22117
rect 23560 22151 23612 22160
rect 23560 22117 23569 22151
rect 23569 22117 23603 22151
rect 23603 22117 23612 22151
rect 23560 22108 23612 22117
rect 17396 22040 17448 22092
rect 17764 22083 17816 22092
rect 17764 22049 17773 22083
rect 17773 22049 17807 22083
rect 17807 22049 17816 22083
rect 17764 22040 17816 22049
rect 24480 22083 24532 22092
rect 24480 22049 24498 22083
rect 24498 22049 24532 22083
rect 24480 22040 24532 22049
rect 9484 22015 9536 22024
rect 9484 21981 9493 22015
rect 9493 21981 9527 22015
rect 9527 21981 9536 22015
rect 9484 21972 9536 21981
rect 15924 21972 15976 22024
rect 20524 22015 20576 22024
rect 20524 21981 20533 22015
rect 20533 21981 20567 22015
rect 20567 21981 20576 22015
rect 20524 21972 20576 21981
rect 20800 22015 20852 22024
rect 20800 21981 20809 22015
rect 20809 21981 20843 22015
rect 20843 21981 20852 22015
rect 20800 21972 20852 21981
rect 22548 21972 22600 22024
rect 2216 21836 2268 21888
rect 12060 21836 12112 21888
rect 12704 21879 12756 21888
rect 12704 21845 12713 21879
rect 12713 21845 12747 21879
rect 12747 21845 12756 21879
rect 12704 21836 12756 21845
rect 15832 21879 15884 21888
rect 15832 21845 15841 21879
rect 15841 21845 15875 21879
rect 15875 21845 15884 21879
rect 15832 21836 15884 21845
rect 18500 21879 18552 21888
rect 18500 21845 18509 21879
rect 18509 21845 18543 21879
rect 18543 21845 18552 21879
rect 18500 21836 18552 21845
rect 24388 21836 24440 21888
rect 5176 21734 5228 21786
rect 5240 21734 5292 21786
rect 5304 21734 5356 21786
rect 5368 21734 5420 21786
rect 14510 21734 14562 21786
rect 14574 21734 14626 21786
rect 14638 21734 14690 21786
rect 14702 21734 14754 21786
rect 23843 21734 23895 21786
rect 23907 21734 23959 21786
rect 23971 21734 24023 21786
rect 24035 21734 24087 21786
rect 1020 21632 1072 21684
rect 4148 21632 4200 21684
rect 9576 21632 9628 21684
rect 10220 21632 10272 21684
rect 11324 21632 11376 21684
rect 12520 21675 12572 21684
rect 12520 21641 12529 21675
rect 12529 21641 12563 21675
rect 12563 21641 12572 21675
rect 12520 21632 12572 21641
rect 13808 21632 13860 21684
rect 14912 21675 14964 21684
rect 14912 21641 14921 21675
rect 14921 21641 14955 21675
rect 14955 21641 14964 21675
rect 14912 21632 14964 21641
rect 17764 21675 17816 21684
rect 17764 21641 17773 21675
rect 17773 21641 17807 21675
rect 17807 21641 17816 21675
rect 17764 21632 17816 21641
rect 20616 21675 20668 21684
rect 20616 21641 20625 21675
rect 20625 21641 20659 21675
rect 20659 21641 20668 21675
rect 20616 21632 20668 21641
rect 21720 21632 21772 21684
rect 22548 21675 22600 21684
rect 22548 21641 22557 21675
rect 22557 21641 22591 21675
rect 22591 21641 22600 21675
rect 22548 21632 22600 21641
rect 24480 21675 24532 21684
rect 24480 21641 24489 21675
rect 24489 21641 24523 21675
rect 24523 21641 24532 21675
rect 24480 21632 24532 21641
rect 25308 21675 25360 21684
rect 25308 21641 25317 21675
rect 25317 21641 25351 21675
rect 25351 21641 25360 21675
rect 25308 21632 25360 21641
rect 15924 21564 15976 21616
rect 20524 21564 20576 21616
rect 7460 21539 7512 21548
rect 7460 21505 7469 21539
rect 7469 21505 7503 21539
rect 7503 21505 7512 21539
rect 7460 21496 7512 21505
rect 9484 21496 9536 21548
rect 15096 21496 15148 21548
rect 18960 21539 19012 21548
rect 18960 21505 18969 21539
rect 18969 21505 19003 21539
rect 19003 21505 19012 21539
rect 18960 21496 19012 21505
rect 23008 21496 23060 21548
rect 4148 21428 4200 21480
rect 12520 21428 12572 21480
rect 13624 21428 13676 21480
rect 20156 21428 20208 21480
rect 20708 21471 20760 21480
rect 20708 21437 20717 21471
rect 20717 21437 20751 21471
rect 20751 21437 20760 21471
rect 20708 21428 20760 21437
rect 7644 21360 7696 21412
rect 9024 21403 9076 21412
rect 9024 21369 9033 21403
rect 9033 21369 9067 21403
rect 9067 21369 9076 21403
rect 9024 21360 9076 21369
rect 4976 21292 5028 21344
rect 8748 21335 8800 21344
rect 8748 21301 8757 21335
rect 8757 21301 8791 21335
rect 8791 21301 8800 21335
rect 11692 21360 11744 21412
rect 18500 21403 18552 21412
rect 18500 21369 18509 21403
rect 18509 21369 18543 21403
rect 18543 21369 18552 21403
rect 18500 21360 18552 21369
rect 18592 21403 18644 21412
rect 18592 21369 18601 21403
rect 18601 21369 18635 21403
rect 18635 21369 18644 21403
rect 18592 21360 18644 21369
rect 8748 21292 8800 21301
rect 12244 21292 12296 21344
rect 20248 21335 20300 21344
rect 20248 21301 20257 21335
rect 20257 21301 20291 21335
rect 20291 21301 20300 21335
rect 20248 21292 20300 21301
rect 21628 21292 21680 21344
rect 23284 21471 23336 21480
rect 23284 21437 23293 21471
rect 23293 21437 23327 21471
rect 23327 21437 23336 21471
rect 23284 21428 23336 21437
rect 25308 21428 25360 21480
rect 24480 21292 24532 21344
rect 9843 21190 9895 21242
rect 9907 21190 9959 21242
rect 9971 21190 10023 21242
rect 10035 21190 10087 21242
rect 19176 21190 19228 21242
rect 19240 21190 19292 21242
rect 19304 21190 19356 21242
rect 19368 21190 19420 21242
rect 7460 21131 7512 21140
rect 7460 21097 7469 21131
rect 7469 21097 7503 21131
rect 7503 21097 7512 21131
rect 7460 21088 7512 21097
rect 10220 21131 10272 21140
rect 10220 21097 10229 21131
rect 10229 21097 10263 21131
rect 10263 21097 10272 21131
rect 10220 21088 10272 21097
rect 11324 21088 11376 21140
rect 17764 21088 17816 21140
rect 22548 21088 22600 21140
rect 24204 21088 24256 21140
rect 8748 21020 8800 21072
rect 9668 21063 9720 21072
rect 9668 21029 9671 21063
rect 9671 21029 9705 21063
rect 9705 21029 9720 21063
rect 9668 21020 9720 21029
rect 11692 21063 11744 21072
rect 11692 21029 11695 21063
rect 11695 21029 11729 21063
rect 11729 21029 11744 21063
rect 11692 21020 11744 21029
rect 16752 21063 16804 21072
rect 16752 21029 16755 21063
rect 16755 21029 16789 21063
rect 16789 21029 16804 21063
rect 16752 21020 16804 21029
rect 18868 21020 18920 21072
rect 20432 21063 20484 21072
rect 20432 21029 20441 21063
rect 20441 21029 20475 21063
rect 20475 21029 20484 21063
rect 20432 21020 20484 21029
rect 7644 20952 7696 21004
rect 9116 20952 9168 21004
rect 15372 20995 15424 21004
rect 9300 20927 9352 20936
rect 9300 20893 9309 20927
rect 9309 20893 9343 20927
rect 9343 20893 9352 20927
rect 9300 20884 9352 20893
rect 11232 20884 11284 20936
rect 15372 20961 15381 20995
rect 15381 20961 15415 20995
rect 15415 20961 15424 20995
rect 15372 20952 15424 20961
rect 20524 20995 20576 21004
rect 20524 20961 20533 20995
rect 20533 20961 20567 20995
rect 20567 20961 20576 20995
rect 20524 20952 20576 20961
rect 24388 20952 24440 21004
rect 15280 20884 15332 20936
rect 15740 20884 15792 20936
rect 16384 20927 16436 20936
rect 16384 20893 16393 20927
rect 16393 20893 16427 20927
rect 16427 20893 16436 20927
rect 16384 20884 16436 20893
rect 18960 20884 19012 20936
rect 19512 20927 19564 20936
rect 19512 20893 19521 20927
rect 19521 20893 19555 20927
rect 19555 20893 19564 20927
rect 19512 20884 19564 20893
rect 9024 20791 9076 20800
rect 9024 20757 9033 20791
rect 9033 20757 9067 20791
rect 9067 20757 9076 20791
rect 9024 20748 9076 20757
rect 13624 20791 13676 20800
rect 13624 20757 13633 20791
rect 13633 20757 13667 20791
rect 13667 20757 13676 20791
rect 13624 20748 13676 20757
rect 13900 20748 13952 20800
rect 17672 20791 17724 20800
rect 17672 20757 17681 20791
rect 17681 20757 17715 20791
rect 17715 20757 17724 20791
rect 17672 20748 17724 20757
rect 23008 20748 23060 20800
rect 23284 20748 23336 20800
rect 5176 20646 5228 20698
rect 5240 20646 5292 20698
rect 5304 20646 5356 20698
rect 5368 20646 5420 20698
rect 14510 20646 14562 20698
rect 14574 20646 14626 20698
rect 14638 20646 14690 20698
rect 14702 20646 14754 20698
rect 23843 20646 23895 20698
rect 23907 20646 23959 20698
rect 23971 20646 24023 20698
rect 24035 20646 24087 20698
rect 7644 20587 7696 20596
rect 7644 20553 7653 20587
rect 7653 20553 7687 20587
rect 7687 20553 7696 20587
rect 7644 20544 7696 20553
rect 9208 20544 9260 20596
rect 12888 20587 12940 20596
rect 12888 20553 12897 20587
rect 12897 20553 12931 20587
rect 12931 20553 12940 20587
rect 12888 20544 12940 20553
rect 15832 20544 15884 20596
rect 16660 20587 16712 20596
rect 16660 20553 16669 20587
rect 16669 20553 16703 20587
rect 16703 20553 16712 20587
rect 16660 20544 16712 20553
rect 20524 20587 20576 20596
rect 20524 20553 20533 20587
rect 20533 20553 20567 20587
rect 20567 20553 20576 20587
rect 20524 20544 20576 20553
rect 21720 20544 21772 20596
rect 24388 20544 24440 20596
rect 24296 20476 24348 20528
rect 9300 20408 9352 20460
rect 15740 20451 15792 20460
rect 15740 20417 15749 20451
rect 15749 20417 15783 20451
rect 15783 20417 15792 20451
rect 15740 20408 15792 20417
rect 18592 20408 18644 20460
rect 18960 20408 19012 20460
rect 19512 20451 19564 20460
rect 19512 20417 19521 20451
rect 19521 20417 19555 20451
rect 19555 20417 19564 20451
rect 19512 20408 19564 20417
rect 9116 20340 9168 20392
rect 12060 20340 12112 20392
rect 9668 20272 9720 20324
rect 11232 20272 11284 20324
rect 11876 20272 11928 20324
rect 11692 20247 11744 20256
rect 11692 20213 11701 20247
rect 11701 20213 11735 20247
rect 11735 20213 11744 20247
rect 13900 20340 13952 20392
rect 16752 20340 16804 20392
rect 21168 20340 21220 20392
rect 24480 20340 24532 20392
rect 16200 20272 16252 20324
rect 16384 20272 16436 20324
rect 15280 20247 15332 20256
rect 11692 20204 11744 20213
rect 15280 20213 15289 20247
rect 15289 20213 15323 20247
rect 15323 20213 15332 20247
rect 15280 20204 15332 20213
rect 17580 20204 17632 20256
rect 17764 20315 17816 20324
rect 17764 20281 17773 20315
rect 17773 20281 17807 20315
rect 17807 20281 17816 20315
rect 17764 20272 17816 20281
rect 18500 20204 18552 20256
rect 18960 20247 19012 20256
rect 18960 20213 18969 20247
rect 18969 20213 19003 20247
rect 19003 20213 19012 20247
rect 21076 20247 21128 20256
rect 18960 20204 19012 20213
rect 21076 20213 21085 20247
rect 21085 20213 21119 20247
rect 21119 20213 21128 20247
rect 21076 20204 21128 20213
rect 23008 20204 23060 20256
rect 9843 20102 9895 20154
rect 9907 20102 9959 20154
rect 9971 20102 10023 20154
rect 10035 20102 10087 20154
rect 19176 20102 19228 20154
rect 19240 20102 19292 20154
rect 19304 20102 19356 20154
rect 19368 20102 19420 20154
rect 9300 20000 9352 20052
rect 17672 20000 17724 20052
rect 18592 20043 18644 20052
rect 18592 20009 18601 20043
rect 18601 20009 18635 20043
rect 18635 20009 18644 20043
rect 18592 20000 18644 20009
rect 18960 20043 19012 20052
rect 18960 20009 18969 20043
rect 18969 20009 19003 20043
rect 19003 20009 19012 20043
rect 18960 20000 19012 20009
rect 21536 20000 21588 20052
rect 22916 20000 22968 20052
rect 13900 19975 13952 19984
rect 13900 19941 13909 19975
rect 13909 19941 13943 19975
rect 13943 19941 13952 19975
rect 13900 19932 13952 19941
rect 16384 19932 16436 19984
rect 16752 19932 16804 19984
rect 21076 19932 21128 19984
rect 9576 19864 9628 19916
rect 11508 19907 11560 19916
rect 11508 19873 11517 19907
rect 11517 19873 11551 19907
rect 11551 19873 11560 19907
rect 11508 19864 11560 19873
rect 12152 19864 12204 19916
rect 13348 19907 13400 19916
rect 13348 19873 13357 19907
rect 13357 19873 13391 19907
rect 13391 19873 13400 19907
rect 13348 19864 13400 19873
rect 13992 19864 14044 19916
rect 14912 19907 14964 19916
rect 14912 19873 14921 19907
rect 14921 19873 14955 19907
rect 14955 19873 14964 19907
rect 14912 19864 14964 19873
rect 15372 19907 15424 19916
rect 15372 19873 15381 19907
rect 15381 19873 15415 19907
rect 15415 19873 15424 19907
rect 15372 19864 15424 19873
rect 17672 19907 17724 19916
rect 17672 19873 17681 19907
rect 17681 19873 17715 19907
rect 17715 19873 17724 19907
rect 17672 19864 17724 19873
rect 18868 19907 18920 19916
rect 18868 19873 18877 19907
rect 18877 19873 18911 19907
rect 18911 19873 18920 19907
rect 18868 19864 18920 19873
rect 19512 19864 19564 19916
rect 20984 19864 21036 19916
rect 23652 19907 23704 19916
rect 23652 19873 23661 19907
rect 23661 19873 23695 19907
rect 23695 19873 23704 19907
rect 23652 19864 23704 19873
rect 25400 19864 25452 19916
rect 10312 19796 10364 19848
rect 12060 19839 12112 19848
rect 12060 19805 12069 19839
rect 12069 19805 12103 19839
rect 12103 19805 12112 19839
rect 12060 19796 12112 19805
rect 16476 19839 16528 19848
rect 16476 19805 16485 19839
rect 16485 19805 16519 19839
rect 16519 19805 16528 19839
rect 16476 19796 16528 19805
rect 21536 19839 21588 19848
rect 21536 19805 21545 19839
rect 21545 19805 21579 19839
rect 21579 19805 21588 19839
rect 21536 19796 21588 19805
rect 24388 19728 24440 19780
rect 14820 19660 14872 19712
rect 21168 19660 21220 19712
rect 23560 19703 23612 19712
rect 23560 19669 23569 19703
rect 23569 19669 23603 19703
rect 23603 19669 23612 19703
rect 23560 19660 23612 19669
rect 5176 19558 5228 19610
rect 5240 19558 5292 19610
rect 5304 19558 5356 19610
rect 5368 19558 5420 19610
rect 14510 19558 14562 19610
rect 14574 19558 14626 19610
rect 14638 19558 14690 19610
rect 14702 19558 14754 19610
rect 23843 19558 23895 19610
rect 23907 19558 23959 19610
rect 23971 19558 24023 19610
rect 24035 19558 24087 19610
rect 16200 19456 16252 19508
rect 16752 19456 16804 19508
rect 18868 19499 18920 19508
rect 18868 19465 18877 19499
rect 18877 19465 18911 19499
rect 18911 19465 18920 19499
rect 18868 19456 18920 19465
rect 20984 19499 21036 19508
rect 20984 19465 20993 19499
rect 20993 19465 21027 19499
rect 21027 19465 21036 19499
rect 20984 19456 21036 19465
rect 25400 19499 25452 19508
rect 25400 19465 25409 19499
rect 25409 19465 25443 19499
rect 25443 19465 25452 19499
rect 25400 19456 25452 19465
rect 13348 19388 13400 19440
rect 14912 19431 14964 19440
rect 14912 19397 14921 19431
rect 14921 19397 14955 19431
rect 14955 19397 14964 19431
rect 14912 19388 14964 19397
rect 16752 19320 16804 19372
rect 9484 19295 9536 19304
rect 9484 19261 9493 19295
rect 9493 19261 9527 19295
rect 9527 19261 9536 19295
rect 9484 19252 9536 19261
rect 9576 19252 9628 19304
rect 11508 19295 11560 19304
rect 11508 19261 11517 19295
rect 11517 19261 11551 19295
rect 11551 19261 11560 19295
rect 11508 19252 11560 19261
rect 12060 19295 12112 19304
rect 12060 19261 12069 19295
rect 12069 19261 12103 19295
rect 12103 19261 12112 19295
rect 12060 19252 12112 19261
rect 9208 19116 9260 19168
rect 10312 19159 10364 19168
rect 10312 19125 10321 19159
rect 10321 19125 10355 19159
rect 10355 19125 10364 19159
rect 10312 19116 10364 19125
rect 12152 19184 12204 19236
rect 13256 19252 13308 19304
rect 13716 19295 13768 19304
rect 13716 19261 13725 19295
rect 13725 19261 13759 19295
rect 13759 19261 13768 19295
rect 13716 19252 13768 19261
rect 13992 19295 14044 19304
rect 13992 19261 14001 19295
rect 14001 19261 14035 19295
rect 14035 19261 14044 19295
rect 13992 19252 14044 19261
rect 15280 19295 15332 19304
rect 15280 19261 15289 19295
rect 15289 19261 15323 19295
rect 15323 19261 15332 19295
rect 15280 19252 15332 19261
rect 15556 19252 15608 19304
rect 16476 19252 16528 19304
rect 13164 19227 13216 19236
rect 13164 19193 13173 19227
rect 13173 19193 13207 19227
rect 13207 19193 13216 19227
rect 13164 19184 13216 19193
rect 17580 19295 17632 19304
rect 17580 19261 17589 19295
rect 17589 19261 17623 19295
rect 17623 19261 17632 19295
rect 17580 19252 17632 19261
rect 18868 19252 18920 19304
rect 19788 19295 19840 19304
rect 19788 19261 19797 19295
rect 19797 19261 19831 19295
rect 19831 19261 19840 19295
rect 19788 19252 19840 19261
rect 20708 19295 20760 19304
rect 20708 19261 20717 19295
rect 20717 19261 20751 19295
rect 20751 19261 20760 19295
rect 20708 19252 20760 19261
rect 22272 19252 22324 19304
rect 23652 19320 23704 19372
rect 24204 19320 24256 19372
rect 24480 19320 24532 19372
rect 26872 19252 26924 19304
rect 18960 19184 19012 19236
rect 21076 19184 21128 19236
rect 23376 19227 23428 19236
rect 23376 19193 23385 19227
rect 23385 19193 23419 19227
rect 23419 19193 23428 19227
rect 23376 19184 23428 19193
rect 11968 19116 12020 19168
rect 13624 19159 13676 19168
rect 13624 19125 13633 19159
rect 13633 19125 13667 19159
rect 13667 19125 13676 19159
rect 13624 19116 13676 19125
rect 21628 19116 21680 19168
rect 23560 19184 23612 19236
rect 24296 19116 24348 19168
rect 9843 19014 9895 19066
rect 9907 19014 9959 19066
rect 9971 19014 10023 19066
rect 10035 19014 10087 19066
rect 19176 19014 19228 19066
rect 19240 19014 19292 19066
rect 19304 19014 19356 19066
rect 19368 19014 19420 19066
rect 13992 18912 14044 18964
rect 18500 18912 18552 18964
rect 23376 18955 23428 18964
rect 23376 18921 23385 18955
rect 23385 18921 23419 18955
rect 23419 18921 23428 18955
rect 23376 18912 23428 18921
rect 9208 18844 9260 18896
rect 9852 18887 9904 18896
rect 9852 18853 9861 18887
rect 9861 18853 9895 18887
rect 9895 18853 9904 18887
rect 9852 18844 9904 18853
rect 10220 18844 10272 18896
rect 14912 18844 14964 18896
rect 17580 18887 17632 18896
rect 17580 18853 17589 18887
rect 17589 18853 17623 18887
rect 17623 18853 17632 18887
rect 17580 18844 17632 18853
rect 19788 18887 19840 18896
rect 19788 18853 19797 18887
rect 19797 18853 19831 18887
rect 19831 18853 19840 18887
rect 19788 18844 19840 18853
rect 21168 18887 21220 18896
rect 21168 18853 21177 18887
rect 21177 18853 21211 18887
rect 21211 18853 21220 18887
rect 21168 18844 21220 18853
rect 23652 18887 23704 18896
rect 23652 18853 23661 18887
rect 23661 18853 23695 18887
rect 23695 18853 23704 18887
rect 23652 18844 23704 18853
rect 24204 18887 24256 18896
rect 24204 18853 24213 18887
rect 24213 18853 24247 18887
rect 24247 18853 24256 18887
rect 24204 18844 24256 18853
rect 15280 18819 15332 18828
rect 10680 18708 10732 18760
rect 11324 18751 11376 18760
rect 11324 18717 11333 18751
rect 11333 18717 11367 18751
rect 11367 18717 11376 18751
rect 11324 18708 11376 18717
rect 11968 18751 12020 18760
rect 11968 18717 11977 18751
rect 11977 18717 12011 18751
rect 12011 18717 12020 18751
rect 11968 18708 12020 18717
rect 13716 18708 13768 18760
rect 15280 18785 15289 18819
rect 15289 18785 15323 18819
rect 15323 18785 15332 18819
rect 15280 18776 15332 18785
rect 15832 18819 15884 18828
rect 15832 18785 15841 18819
rect 15841 18785 15875 18819
rect 15875 18785 15884 18819
rect 15832 18776 15884 18785
rect 18868 18819 18920 18828
rect 14636 18751 14688 18760
rect 14636 18717 14645 18751
rect 14645 18717 14679 18751
rect 14679 18717 14688 18751
rect 14636 18708 14688 18717
rect 18868 18785 18877 18819
rect 18877 18785 18911 18819
rect 18911 18785 18920 18819
rect 18868 18776 18920 18785
rect 19052 18776 19104 18828
rect 20708 18819 20760 18828
rect 20708 18785 20717 18819
rect 20717 18785 20751 18819
rect 20751 18785 20760 18819
rect 20708 18776 20760 18785
rect 20984 18819 21036 18828
rect 20984 18785 20993 18819
rect 20993 18785 21027 18819
rect 21027 18785 21036 18819
rect 20984 18776 21036 18785
rect 9576 18615 9628 18624
rect 9576 18581 9585 18615
rect 9585 18581 9619 18615
rect 9619 18581 9628 18615
rect 9576 18572 9628 18581
rect 10588 18572 10640 18624
rect 12060 18572 12112 18624
rect 13624 18615 13676 18624
rect 13624 18581 13633 18615
rect 13633 18581 13667 18615
rect 13667 18581 13676 18615
rect 13624 18572 13676 18581
rect 15556 18572 15608 18624
rect 16568 18708 16620 18760
rect 23560 18751 23612 18760
rect 23560 18717 23569 18751
rect 23569 18717 23603 18751
rect 23603 18717 23612 18751
rect 23560 18708 23612 18717
rect 21352 18572 21404 18624
rect 5176 18470 5228 18522
rect 5240 18470 5292 18522
rect 5304 18470 5356 18522
rect 5368 18470 5420 18522
rect 14510 18470 14562 18522
rect 14574 18470 14626 18522
rect 14638 18470 14690 18522
rect 14702 18470 14754 18522
rect 23843 18470 23895 18522
rect 23907 18470 23959 18522
rect 23971 18470 24023 18522
rect 24035 18470 24087 18522
rect 9852 18368 9904 18420
rect 13624 18368 13676 18420
rect 13992 18411 14044 18420
rect 13992 18377 14001 18411
rect 14001 18377 14035 18411
rect 14035 18377 14044 18411
rect 13992 18368 14044 18377
rect 15832 18411 15884 18420
rect 15832 18377 15841 18411
rect 15841 18377 15875 18411
rect 15875 18377 15884 18411
rect 15832 18368 15884 18377
rect 16108 18368 16160 18420
rect 16568 18411 16620 18420
rect 16568 18377 16577 18411
rect 16577 18377 16611 18411
rect 16611 18377 16620 18411
rect 16568 18368 16620 18377
rect 18960 18368 19012 18420
rect 20156 18411 20208 18420
rect 20156 18377 20165 18411
rect 20165 18377 20199 18411
rect 20199 18377 20208 18411
rect 20156 18368 20208 18377
rect 21076 18368 21128 18420
rect 21628 18368 21680 18420
rect 22272 18411 22324 18420
rect 22272 18377 22281 18411
rect 22281 18377 22315 18411
rect 22315 18377 22324 18411
rect 22272 18368 22324 18377
rect 23560 18368 23612 18420
rect 10588 18300 10640 18352
rect 12612 18343 12664 18352
rect 12612 18309 12621 18343
rect 12621 18309 12655 18343
rect 12655 18309 12664 18343
rect 12612 18300 12664 18309
rect 10680 18275 10732 18284
rect 10680 18241 10689 18275
rect 10689 18241 10723 18275
rect 10723 18241 10732 18275
rect 12060 18275 12112 18284
rect 10680 18232 10732 18241
rect 12060 18241 12069 18275
rect 12069 18241 12103 18275
rect 12103 18241 12112 18275
rect 12060 18232 12112 18241
rect 13440 18232 13492 18284
rect 13992 18232 14044 18284
rect 19512 18232 19564 18284
rect 24388 18232 24440 18284
rect 10220 18164 10272 18216
rect 18224 18207 18276 18216
rect 18224 18173 18233 18207
rect 18233 18173 18267 18207
rect 18267 18173 18276 18207
rect 18224 18164 18276 18173
rect 21352 18207 21404 18216
rect 21352 18173 21361 18207
rect 21361 18173 21395 18207
rect 21395 18173 21404 18207
rect 21352 18164 21404 18173
rect 11784 18139 11836 18148
rect 11784 18105 11793 18139
rect 11793 18105 11827 18139
rect 11827 18105 11836 18139
rect 11784 18096 11836 18105
rect 13716 18096 13768 18148
rect 18960 18096 19012 18148
rect 21628 18096 21680 18148
rect 23928 18139 23980 18148
rect 23928 18105 23937 18139
rect 23937 18105 23971 18139
rect 23971 18105 23980 18139
rect 23928 18096 23980 18105
rect 13440 18071 13492 18080
rect 13440 18037 13449 18071
rect 13449 18037 13483 18071
rect 13483 18037 13492 18071
rect 13440 18028 13492 18037
rect 14544 18071 14596 18080
rect 14544 18037 14553 18071
rect 14553 18037 14587 18071
rect 14587 18037 14596 18071
rect 14544 18028 14596 18037
rect 15188 18028 15240 18080
rect 16200 18071 16252 18080
rect 16200 18037 16209 18071
rect 16209 18037 16243 18071
rect 16243 18037 16252 18071
rect 16200 18028 16252 18037
rect 18868 18028 18920 18080
rect 19052 18028 19104 18080
rect 20708 18028 20760 18080
rect 23652 18071 23704 18080
rect 23652 18037 23661 18071
rect 23661 18037 23695 18071
rect 23695 18037 23704 18071
rect 23652 18028 23704 18037
rect 9843 17926 9895 17978
rect 9907 17926 9959 17978
rect 9971 17926 10023 17978
rect 10035 17926 10087 17978
rect 19176 17926 19228 17978
rect 19240 17926 19292 17978
rect 19304 17926 19356 17978
rect 19368 17926 19420 17978
rect 10220 17824 10272 17876
rect 13808 17867 13860 17876
rect 13808 17833 13817 17867
rect 13817 17833 13851 17867
rect 13851 17833 13860 17867
rect 13808 17824 13860 17833
rect 13992 17824 14044 17876
rect 14544 17867 14596 17876
rect 14544 17833 14553 17867
rect 14553 17833 14587 17867
rect 14587 17833 14596 17867
rect 14544 17824 14596 17833
rect 16108 17824 16160 17876
rect 23560 17867 23612 17876
rect 23560 17833 23569 17867
rect 23569 17833 23603 17867
rect 23603 17833 23612 17867
rect 23560 17824 23612 17833
rect 9668 17756 9720 17808
rect 11600 17756 11652 17808
rect 12612 17756 12664 17808
rect 9484 17663 9536 17672
rect 9484 17629 9493 17663
rect 9493 17629 9527 17663
rect 9527 17629 9536 17663
rect 9484 17620 9536 17629
rect 11324 17620 11376 17672
rect 10680 17527 10732 17536
rect 10680 17493 10689 17527
rect 10689 17493 10723 17527
rect 10723 17493 10732 17527
rect 10680 17484 10732 17493
rect 12704 17527 12756 17536
rect 12704 17493 12713 17527
rect 12713 17493 12747 17527
rect 12747 17493 12756 17527
rect 12704 17484 12756 17493
rect 12980 17484 13032 17536
rect 13624 17756 13676 17808
rect 15556 17799 15608 17808
rect 15556 17765 15565 17799
rect 15565 17765 15599 17799
rect 15599 17765 15608 17799
rect 15556 17756 15608 17765
rect 18868 17756 18920 17808
rect 13716 17688 13768 17740
rect 13256 17620 13308 17672
rect 13440 17620 13492 17672
rect 13440 17527 13492 17536
rect 13440 17493 13449 17527
rect 13449 17493 13483 17527
rect 13483 17493 13492 17527
rect 13440 17484 13492 17493
rect 14176 17484 14228 17536
rect 15004 17731 15056 17740
rect 15004 17697 15010 17731
rect 15010 17697 15056 17731
rect 16384 17731 16436 17740
rect 15004 17688 15056 17697
rect 16384 17697 16393 17731
rect 16393 17697 16427 17731
rect 16427 17697 16436 17731
rect 16384 17688 16436 17697
rect 18684 17731 18736 17740
rect 18684 17697 18693 17731
rect 18693 17697 18727 17731
rect 18727 17697 18736 17731
rect 18684 17688 18736 17697
rect 19144 17731 19196 17740
rect 19144 17697 19153 17731
rect 19153 17697 19187 17731
rect 19187 17697 19196 17731
rect 19144 17688 19196 17697
rect 19512 17756 19564 17808
rect 21536 17756 21588 17808
rect 21628 17756 21680 17808
rect 20800 17688 20852 17740
rect 20984 17731 21036 17740
rect 20984 17697 20993 17731
rect 20993 17697 21027 17731
rect 21027 17697 21036 17731
rect 24204 17756 24256 17808
rect 20984 17688 21036 17697
rect 15188 17663 15240 17672
rect 15188 17629 15197 17663
rect 15197 17629 15231 17663
rect 15231 17629 15240 17663
rect 15188 17620 15240 17629
rect 14912 17552 14964 17604
rect 22364 17620 22416 17672
rect 24296 17620 24348 17672
rect 21536 17552 21588 17604
rect 24388 17595 24440 17604
rect 24388 17561 24397 17595
rect 24397 17561 24431 17595
rect 24431 17561 24440 17595
rect 24388 17552 24440 17561
rect 14360 17484 14412 17536
rect 15372 17484 15424 17536
rect 16844 17527 16896 17536
rect 16844 17493 16853 17527
rect 16853 17493 16887 17527
rect 16887 17493 16896 17527
rect 16844 17484 16896 17493
rect 17856 17484 17908 17536
rect 20156 17527 20208 17536
rect 20156 17493 20165 17527
rect 20165 17493 20199 17527
rect 20199 17493 20208 17527
rect 20156 17484 20208 17493
rect 21444 17527 21496 17536
rect 21444 17493 21453 17527
rect 21453 17493 21487 17527
rect 21487 17493 21496 17527
rect 21444 17484 21496 17493
rect 5176 17382 5228 17434
rect 5240 17382 5292 17434
rect 5304 17382 5356 17434
rect 5368 17382 5420 17434
rect 14510 17382 14562 17434
rect 14574 17382 14626 17434
rect 14638 17382 14690 17434
rect 14702 17382 14754 17434
rect 23843 17382 23895 17434
rect 23907 17382 23959 17434
rect 23971 17382 24023 17434
rect 24035 17382 24087 17434
rect 9668 17323 9720 17332
rect 9668 17289 9677 17323
rect 9677 17289 9711 17323
rect 9711 17289 9720 17323
rect 9668 17280 9720 17289
rect 11600 17323 11652 17332
rect 11600 17289 11609 17323
rect 11609 17289 11643 17323
rect 11643 17289 11652 17323
rect 11600 17280 11652 17289
rect 12980 17323 13032 17332
rect 12980 17289 13004 17323
rect 13004 17289 13032 17323
rect 12980 17280 13032 17289
rect 13348 17280 13400 17332
rect 14268 17280 14320 17332
rect 12520 17212 12572 17264
rect 13992 17212 14044 17264
rect 14636 17255 14688 17264
rect 14636 17221 14645 17255
rect 14645 17221 14679 17255
rect 14679 17221 14688 17255
rect 14636 17212 14688 17221
rect 15924 17280 15976 17332
rect 19144 17280 19196 17332
rect 21536 17280 21588 17332
rect 23652 17323 23704 17332
rect 23652 17289 23661 17323
rect 23661 17289 23695 17323
rect 23695 17289 23704 17323
rect 23652 17280 23704 17289
rect 24480 17280 24532 17332
rect 25492 17323 25544 17332
rect 25492 17289 25501 17323
rect 25501 17289 25535 17323
rect 25535 17289 25544 17323
rect 25492 17280 25544 17289
rect 15372 17255 15424 17264
rect 15372 17221 15381 17255
rect 15381 17221 15415 17255
rect 15415 17221 15424 17255
rect 15372 17212 15424 17221
rect 16200 17255 16252 17264
rect 16200 17221 16209 17255
rect 16209 17221 16243 17255
rect 16243 17221 16252 17255
rect 16200 17212 16252 17221
rect 16384 17212 16436 17264
rect 17212 17212 17264 17264
rect 18224 17212 18276 17264
rect 9484 17144 9536 17196
rect 9024 17076 9076 17128
rect 10404 17144 10456 17196
rect 13256 17144 13308 17196
rect 15188 17144 15240 17196
rect 16844 17144 16896 17196
rect 17856 17144 17908 17196
rect 17948 17187 18000 17196
rect 17948 17153 17957 17187
rect 17957 17153 17991 17187
rect 17991 17153 18000 17187
rect 21352 17187 21404 17196
rect 17948 17144 18000 17153
rect 21352 17153 21361 17187
rect 21361 17153 21395 17187
rect 21395 17153 21404 17187
rect 21352 17144 21404 17153
rect 10680 17076 10732 17128
rect 11784 17076 11836 17128
rect 13440 17076 13492 17128
rect 12704 17008 12756 17060
rect 13164 17008 13216 17060
rect 20800 17119 20852 17128
rect 14360 17051 14412 17060
rect 14360 17017 14369 17051
rect 14369 17017 14403 17051
rect 14403 17017 14412 17051
rect 14360 17008 14412 17017
rect 15648 17008 15700 17060
rect 13256 16940 13308 16992
rect 14176 16983 14228 16992
rect 14176 16949 14185 16983
rect 14185 16949 14219 16983
rect 14219 16949 14228 16983
rect 14176 16940 14228 16949
rect 17304 16983 17356 16992
rect 17304 16949 17313 16983
rect 17313 16949 17347 16983
rect 17347 16949 17356 16983
rect 18040 17008 18092 17060
rect 20800 17085 20809 17119
rect 20809 17085 20843 17119
rect 20843 17085 20852 17119
rect 20800 17076 20852 17085
rect 20892 17076 20944 17128
rect 21444 17076 21496 17128
rect 21628 17076 21680 17128
rect 24204 17076 24256 17128
rect 25492 17076 25544 17128
rect 17304 16940 17356 16949
rect 18684 16940 18736 16992
rect 20708 16940 20760 16992
rect 22364 16983 22416 16992
rect 22364 16949 22373 16983
rect 22373 16949 22407 16983
rect 22407 16949 22416 16983
rect 22364 16940 22416 16949
rect 9843 16838 9895 16890
rect 9907 16838 9959 16890
rect 9971 16838 10023 16890
rect 10035 16838 10087 16890
rect 19176 16838 19228 16890
rect 19240 16838 19292 16890
rect 19304 16838 19356 16890
rect 19368 16838 19420 16890
rect 9024 16736 9076 16788
rect 9484 16779 9536 16788
rect 9484 16745 9493 16779
rect 9493 16745 9527 16779
rect 9527 16745 9536 16779
rect 9484 16736 9536 16745
rect 11324 16779 11376 16788
rect 11324 16745 11333 16779
rect 11333 16745 11367 16779
rect 11367 16745 11376 16779
rect 11324 16736 11376 16745
rect 11600 16736 11652 16788
rect 12980 16736 13032 16788
rect 13808 16779 13860 16788
rect 13808 16745 13817 16779
rect 13817 16745 13851 16779
rect 13851 16745 13860 16779
rect 13808 16736 13860 16745
rect 15004 16779 15056 16788
rect 15004 16745 15013 16779
rect 15013 16745 15047 16779
rect 15047 16745 15056 16779
rect 15004 16736 15056 16745
rect 18684 16779 18736 16788
rect 18684 16745 18693 16779
rect 18693 16745 18727 16779
rect 18727 16745 18736 16779
rect 18684 16736 18736 16745
rect 24296 16736 24348 16788
rect 10680 16711 10732 16720
rect 10680 16677 10689 16711
rect 10689 16677 10723 16711
rect 10723 16677 10732 16711
rect 10680 16668 10732 16677
rect 12612 16668 12664 16720
rect 14176 16668 14228 16720
rect 10220 16643 10272 16652
rect 10220 16609 10229 16643
rect 10229 16609 10263 16643
rect 10263 16609 10272 16643
rect 10220 16600 10272 16609
rect 10404 16643 10456 16652
rect 10404 16609 10413 16643
rect 10413 16609 10447 16643
rect 10447 16609 10456 16643
rect 10404 16600 10456 16609
rect 11784 16643 11836 16652
rect 11784 16609 11793 16643
rect 11793 16609 11827 16643
rect 11827 16609 11836 16643
rect 11784 16600 11836 16609
rect 13164 16643 13216 16652
rect 13164 16609 13173 16643
rect 13173 16609 13207 16643
rect 13207 16609 13216 16643
rect 13164 16600 13216 16609
rect 14912 16668 14964 16720
rect 15648 16711 15700 16720
rect 15648 16677 15657 16711
rect 15657 16677 15691 16711
rect 15691 16677 15700 16711
rect 15648 16668 15700 16677
rect 16016 16711 16068 16720
rect 16016 16677 16025 16711
rect 16025 16677 16059 16711
rect 16059 16677 16068 16711
rect 16016 16668 16068 16677
rect 16200 16668 16252 16720
rect 15004 16600 15056 16652
rect 13256 16532 13308 16584
rect 17948 16668 18000 16720
rect 18776 16668 18828 16720
rect 22364 16668 22416 16720
rect 24388 16668 24440 16720
rect 17580 16643 17632 16652
rect 17580 16609 17589 16643
rect 17589 16609 17623 16643
rect 17623 16609 17632 16643
rect 17580 16600 17632 16609
rect 18040 16600 18092 16652
rect 18224 16643 18276 16652
rect 18224 16609 18233 16643
rect 18233 16609 18267 16643
rect 18267 16609 18276 16643
rect 18224 16600 18276 16609
rect 19052 16643 19104 16652
rect 19052 16609 19061 16643
rect 19061 16609 19095 16643
rect 19095 16609 19104 16643
rect 19052 16600 19104 16609
rect 20708 16643 20760 16652
rect 20708 16609 20717 16643
rect 20717 16609 20751 16643
rect 20751 16609 20760 16643
rect 20708 16600 20760 16609
rect 20892 16600 20944 16652
rect 23192 16643 23244 16652
rect 23192 16609 23236 16643
rect 23236 16609 23244 16643
rect 23192 16600 23244 16609
rect 23744 16600 23796 16652
rect 24296 16643 24348 16652
rect 24296 16609 24314 16643
rect 24314 16609 24348 16643
rect 24296 16600 24348 16609
rect 14268 16464 14320 16516
rect 12980 16396 13032 16448
rect 14360 16439 14412 16448
rect 14360 16405 14369 16439
rect 14369 16405 14403 16439
rect 14403 16405 14412 16439
rect 14360 16396 14412 16405
rect 23008 16396 23060 16448
rect 5176 16294 5228 16346
rect 5240 16294 5292 16346
rect 5304 16294 5356 16346
rect 5368 16294 5420 16346
rect 14510 16294 14562 16346
rect 14574 16294 14626 16346
rect 14638 16294 14690 16346
rect 14702 16294 14754 16346
rect 23843 16294 23895 16346
rect 23907 16294 23959 16346
rect 23971 16294 24023 16346
rect 24035 16294 24087 16346
rect 9208 16192 9260 16244
rect 10220 16192 10272 16244
rect 10772 16235 10824 16244
rect 10772 16201 10781 16235
rect 10781 16201 10815 16235
rect 10815 16201 10824 16235
rect 10772 16192 10824 16201
rect 11784 16192 11836 16244
rect 12980 16192 13032 16244
rect 14084 16192 14136 16244
rect 14820 16192 14872 16244
rect 15004 16192 15056 16244
rect 18868 16235 18920 16244
rect 18868 16201 18877 16235
rect 18877 16201 18911 16235
rect 18911 16201 18920 16235
rect 24296 16235 24348 16244
rect 18868 16192 18920 16201
rect 13440 16056 13492 16108
rect 14268 16056 14320 16108
rect 15188 16056 15240 16108
rect 17304 16056 17356 16108
rect 24296 16201 24305 16235
rect 24305 16201 24339 16235
rect 24339 16201 24348 16235
rect 24296 16192 24348 16201
rect 24940 16235 24992 16244
rect 24940 16201 24949 16235
rect 24949 16201 24983 16235
rect 24983 16201 24992 16235
rect 24940 16192 24992 16201
rect 20156 16099 20208 16108
rect 20156 16065 20165 16099
rect 20165 16065 20199 16099
rect 20199 16065 20208 16099
rect 20156 16056 20208 16065
rect 25032 16056 25084 16108
rect 16200 15988 16252 16040
rect 17948 15988 18000 16040
rect 14360 15920 14412 15972
rect 18592 15963 18644 15972
rect 18592 15929 18601 15963
rect 18601 15929 18635 15963
rect 18635 15929 18644 15963
rect 18592 15920 18644 15929
rect 10220 15852 10272 15904
rect 12520 15895 12572 15904
rect 12520 15861 12529 15895
rect 12529 15861 12563 15895
rect 12563 15861 12572 15895
rect 12520 15852 12572 15861
rect 13256 15895 13308 15904
rect 13256 15861 13265 15895
rect 13265 15861 13299 15895
rect 13299 15861 13308 15895
rect 13256 15852 13308 15861
rect 15188 15852 15240 15904
rect 17304 15895 17356 15904
rect 17304 15861 17313 15895
rect 17313 15861 17347 15895
rect 17347 15861 17356 15895
rect 17304 15852 17356 15861
rect 24388 15988 24440 16040
rect 20708 15963 20760 15972
rect 20708 15929 20717 15963
rect 20717 15929 20751 15963
rect 20751 15929 20760 15963
rect 20708 15920 20760 15929
rect 21444 15920 21496 15972
rect 23376 15963 23428 15972
rect 23376 15929 23385 15963
rect 23385 15929 23419 15963
rect 23419 15929 23428 15963
rect 23928 15963 23980 15972
rect 23376 15920 23428 15929
rect 23928 15929 23937 15963
rect 23937 15929 23971 15963
rect 23971 15929 23980 15963
rect 23928 15920 23980 15929
rect 20892 15852 20944 15904
rect 9843 15750 9895 15802
rect 9907 15750 9959 15802
rect 9971 15750 10023 15802
rect 10035 15750 10087 15802
rect 19176 15750 19228 15802
rect 19240 15750 19292 15802
rect 19304 15750 19356 15802
rect 19368 15750 19420 15802
rect 14084 15691 14136 15700
rect 14084 15657 14093 15691
rect 14093 15657 14127 15691
rect 14127 15657 14136 15691
rect 14084 15648 14136 15657
rect 16200 15691 16252 15700
rect 16200 15657 16209 15691
rect 16209 15657 16243 15691
rect 16243 15657 16252 15691
rect 16200 15648 16252 15657
rect 17948 15691 18000 15700
rect 17948 15657 17957 15691
rect 17957 15657 17991 15691
rect 17991 15657 18000 15691
rect 17948 15648 18000 15657
rect 18224 15691 18276 15700
rect 18224 15657 18233 15691
rect 18233 15657 18267 15691
rect 18267 15657 18276 15691
rect 18224 15648 18276 15657
rect 23376 15648 23428 15700
rect 15740 15580 15792 15632
rect 16108 15580 16160 15632
rect 18592 15623 18644 15632
rect 18592 15589 18601 15623
rect 18601 15589 18635 15623
rect 18635 15589 18644 15623
rect 18592 15580 18644 15589
rect 20156 15580 20208 15632
rect 21904 15623 21956 15632
rect 21904 15589 21913 15623
rect 21913 15589 21947 15623
rect 21947 15589 21956 15623
rect 21904 15580 21956 15589
rect 23192 15580 23244 15632
rect 23928 15580 23980 15632
rect 16752 15512 16804 15564
rect 23376 15555 23428 15564
rect 23376 15521 23385 15555
rect 23385 15521 23419 15555
rect 23419 15521 23428 15555
rect 23376 15512 23428 15521
rect 24848 15555 24900 15564
rect 24848 15521 24892 15555
rect 24892 15521 24900 15555
rect 24848 15512 24900 15521
rect 14912 15487 14964 15496
rect 14912 15453 14921 15487
rect 14921 15453 14955 15487
rect 14955 15453 14964 15487
rect 14912 15444 14964 15453
rect 16660 15487 16712 15496
rect 16660 15453 16669 15487
rect 16669 15453 16703 15487
rect 16703 15453 16712 15487
rect 16660 15444 16712 15453
rect 18776 15444 18828 15496
rect 20524 15444 20576 15496
rect 21812 15487 21864 15496
rect 21812 15453 21821 15487
rect 21821 15453 21855 15487
rect 21855 15453 21864 15487
rect 21812 15444 21864 15453
rect 13164 15308 13216 15360
rect 13348 15308 13400 15360
rect 14360 15308 14412 15360
rect 18960 15308 19012 15360
rect 20984 15351 21036 15360
rect 20984 15317 20993 15351
rect 20993 15317 21027 15351
rect 21027 15317 21036 15351
rect 20984 15308 21036 15317
rect 24296 15308 24348 15360
rect 5176 15206 5228 15258
rect 5240 15206 5292 15258
rect 5304 15206 5356 15258
rect 5368 15206 5420 15258
rect 14510 15206 14562 15258
rect 14574 15206 14626 15258
rect 14638 15206 14690 15258
rect 14702 15206 14754 15258
rect 23843 15206 23895 15258
rect 23907 15206 23959 15258
rect 23971 15206 24023 15258
rect 24035 15206 24087 15258
rect 15740 15147 15792 15156
rect 15740 15113 15749 15147
rect 15749 15113 15783 15147
rect 15783 15113 15792 15147
rect 15740 15104 15792 15113
rect 16752 15147 16804 15156
rect 16752 15113 16761 15147
rect 16761 15113 16795 15147
rect 16795 15113 16804 15147
rect 16752 15104 16804 15113
rect 17212 15147 17264 15156
rect 17212 15113 17221 15147
rect 17221 15113 17255 15147
rect 17255 15113 17264 15147
rect 17212 15104 17264 15113
rect 18592 15147 18644 15156
rect 18592 15113 18601 15147
rect 18601 15113 18635 15147
rect 18635 15113 18644 15147
rect 18592 15104 18644 15113
rect 19052 15147 19104 15156
rect 19052 15113 19061 15147
rect 19061 15113 19095 15147
rect 19095 15113 19104 15147
rect 19052 15104 19104 15113
rect 21904 15147 21956 15156
rect 21904 15113 21913 15147
rect 21913 15113 21947 15147
rect 21947 15113 21956 15147
rect 21904 15104 21956 15113
rect 23376 15147 23428 15156
rect 23376 15113 23385 15147
rect 23385 15113 23419 15147
rect 23419 15113 23428 15147
rect 23376 15104 23428 15113
rect 21812 15036 21864 15088
rect 17672 15011 17724 15020
rect 17672 14977 17681 15011
rect 17681 14977 17715 15011
rect 17715 14977 17724 15011
rect 17672 14968 17724 14977
rect 14360 14900 14412 14952
rect 14636 14943 14688 14952
rect 14636 14909 14645 14943
rect 14645 14909 14679 14943
rect 14679 14909 14688 14943
rect 14636 14900 14688 14909
rect 15004 14900 15056 14952
rect 15188 14943 15240 14952
rect 15188 14909 15197 14943
rect 15197 14909 15231 14943
rect 15231 14909 15240 14943
rect 15188 14900 15240 14909
rect 14912 14832 14964 14884
rect 13900 14807 13952 14816
rect 13900 14773 13909 14807
rect 13909 14773 13943 14807
rect 13943 14773 13952 14807
rect 13900 14764 13952 14773
rect 15464 14807 15516 14816
rect 15464 14773 15473 14807
rect 15473 14773 15507 14807
rect 15507 14773 15516 14807
rect 15464 14764 15516 14773
rect 17212 14900 17264 14952
rect 20984 14943 21036 14952
rect 20984 14909 20993 14943
rect 20993 14909 21027 14943
rect 21027 14909 21036 14943
rect 20984 14900 21036 14909
rect 22088 14900 22140 14952
rect 24296 15104 24348 15156
rect 17764 14875 17816 14884
rect 17764 14841 17773 14875
rect 17773 14841 17807 14875
rect 17807 14841 17816 14875
rect 17764 14832 17816 14841
rect 18960 14832 19012 14884
rect 19052 14764 19104 14816
rect 20708 14832 20760 14884
rect 21536 14832 21588 14884
rect 24204 14764 24256 14816
rect 24848 14807 24900 14816
rect 24848 14773 24857 14807
rect 24857 14773 24891 14807
rect 24891 14773 24900 14807
rect 24848 14764 24900 14773
rect 9843 14662 9895 14714
rect 9907 14662 9959 14714
rect 9971 14662 10023 14714
rect 10035 14662 10087 14714
rect 19176 14662 19228 14714
rect 19240 14662 19292 14714
rect 19304 14662 19356 14714
rect 19368 14662 19420 14714
rect 13900 14560 13952 14612
rect 14912 14603 14964 14612
rect 14912 14569 14921 14603
rect 14921 14569 14955 14603
rect 14955 14569 14964 14603
rect 14912 14560 14964 14569
rect 15464 14560 15516 14612
rect 16660 14603 16712 14612
rect 16660 14569 16669 14603
rect 16669 14569 16703 14603
rect 16703 14569 16712 14603
rect 16660 14560 16712 14569
rect 17764 14560 17816 14612
rect 22088 14603 22140 14612
rect 22088 14569 22097 14603
rect 22097 14569 22131 14603
rect 22131 14569 22140 14603
rect 22088 14560 22140 14569
rect 23192 14603 23244 14612
rect 23192 14569 23201 14603
rect 23201 14569 23235 14603
rect 23235 14569 23244 14603
rect 23192 14560 23244 14569
rect 15188 14492 15240 14544
rect 16752 14492 16804 14544
rect 17948 14492 18000 14544
rect 20616 14535 20668 14544
rect 20616 14501 20625 14535
rect 20625 14501 20659 14535
rect 20659 14501 20668 14535
rect 20616 14492 20668 14501
rect 14636 14424 14688 14476
rect 15004 14424 15056 14476
rect 15648 14467 15700 14476
rect 15648 14433 15657 14467
rect 15657 14433 15691 14467
rect 15691 14433 15700 14467
rect 15648 14424 15700 14433
rect 21444 14424 21496 14476
rect 22364 14424 22416 14476
rect 24204 14467 24256 14476
rect 15740 14356 15792 14408
rect 18132 14356 18184 14408
rect 20524 14399 20576 14408
rect 20524 14365 20533 14399
rect 20533 14365 20567 14399
rect 20567 14365 20576 14399
rect 20524 14356 20576 14365
rect 20708 14356 20760 14408
rect 21812 14356 21864 14408
rect 24204 14433 24213 14467
rect 24213 14433 24247 14467
rect 24247 14433 24256 14467
rect 24204 14424 24256 14433
rect 23560 14399 23612 14408
rect 23560 14365 23569 14399
rect 23569 14365 23603 14399
rect 23603 14365 23612 14399
rect 23560 14356 23612 14365
rect 19144 14263 19196 14272
rect 19144 14229 19153 14263
rect 19153 14229 19187 14263
rect 19187 14229 19196 14263
rect 19144 14220 19196 14229
rect 21352 14220 21404 14272
rect 5176 14118 5228 14170
rect 5240 14118 5292 14170
rect 5304 14118 5356 14170
rect 5368 14118 5420 14170
rect 14510 14118 14562 14170
rect 14574 14118 14626 14170
rect 14638 14118 14690 14170
rect 14702 14118 14754 14170
rect 23843 14118 23895 14170
rect 23907 14118 23959 14170
rect 23971 14118 24023 14170
rect 24035 14118 24087 14170
rect 14360 14016 14412 14068
rect 15740 14059 15792 14068
rect 15740 14025 15749 14059
rect 15749 14025 15783 14059
rect 15783 14025 15792 14059
rect 15740 14016 15792 14025
rect 17948 14016 18000 14068
rect 20524 14016 20576 14068
rect 23376 14016 23428 14068
rect 24204 14059 24256 14068
rect 24204 14025 24213 14059
rect 24213 14025 24247 14059
rect 24247 14025 24256 14059
rect 24204 14016 24256 14025
rect 13348 13948 13400 14000
rect 13164 13812 13216 13864
rect 12336 13744 12388 13796
rect 14268 13948 14320 14000
rect 22364 13948 22416 14000
rect 23192 13948 23244 14000
rect 14084 13812 14136 13864
rect 14268 13812 14320 13864
rect 14728 13812 14780 13864
rect 15004 13855 15056 13864
rect 15004 13821 15013 13855
rect 15013 13821 15047 13855
rect 15047 13821 15056 13855
rect 15004 13812 15056 13821
rect 20616 13880 20668 13932
rect 15648 13812 15700 13864
rect 18132 13855 18184 13864
rect 18132 13821 18141 13855
rect 18141 13821 18175 13855
rect 18175 13821 18184 13855
rect 18132 13812 18184 13821
rect 19144 13855 19196 13864
rect 19144 13821 19153 13855
rect 19153 13821 19187 13855
rect 19187 13821 19196 13855
rect 19144 13812 19196 13821
rect 21352 13855 21404 13864
rect 21352 13821 21361 13855
rect 21361 13821 21395 13855
rect 21395 13821 21404 13855
rect 21352 13812 21404 13821
rect 21536 13744 21588 13796
rect 23376 13787 23428 13796
rect 23376 13753 23385 13787
rect 23385 13753 23419 13787
rect 23419 13753 23428 13787
rect 23928 13787 23980 13796
rect 23376 13744 23428 13753
rect 23928 13753 23937 13787
rect 23937 13753 23971 13787
rect 23971 13753 23980 13787
rect 23928 13744 23980 13753
rect 15464 13719 15516 13728
rect 15464 13685 15473 13719
rect 15473 13685 15507 13719
rect 15507 13685 15516 13719
rect 15464 13676 15516 13685
rect 23468 13676 23520 13728
rect 9843 13574 9895 13626
rect 9907 13574 9959 13626
rect 9971 13574 10023 13626
rect 10035 13574 10087 13626
rect 19176 13574 19228 13626
rect 19240 13574 19292 13626
rect 19304 13574 19356 13626
rect 19368 13574 19420 13626
rect 12336 13515 12388 13524
rect 12336 13481 12345 13515
rect 12345 13481 12379 13515
rect 12379 13481 12388 13515
rect 12336 13472 12388 13481
rect 15464 13472 15516 13524
rect 24940 13515 24992 13524
rect 13900 13447 13952 13456
rect 13900 13413 13909 13447
rect 13909 13413 13943 13447
rect 13943 13413 13952 13447
rect 13900 13404 13952 13413
rect 15924 13447 15976 13456
rect 15924 13413 15933 13447
rect 15933 13413 15967 13447
rect 15967 13413 15976 13447
rect 15924 13404 15976 13413
rect 18776 13404 18828 13456
rect 21352 13447 21404 13456
rect 21352 13413 21361 13447
rect 21361 13413 21395 13447
rect 21395 13413 21404 13447
rect 21352 13404 21404 13413
rect 23560 13404 23612 13456
rect 23928 13447 23980 13456
rect 23928 13413 23937 13447
rect 23937 13413 23971 13447
rect 23971 13413 23980 13447
rect 23928 13404 23980 13413
rect 24204 13404 24256 13456
rect 24940 13481 24949 13515
rect 24949 13481 24983 13515
rect 24983 13481 24992 13515
rect 24940 13472 24992 13481
rect 12152 13379 12204 13388
rect 12152 13345 12161 13379
rect 12161 13345 12195 13379
rect 12195 13345 12204 13379
rect 12152 13336 12204 13345
rect 13164 13379 13216 13388
rect 13164 13345 13173 13379
rect 13173 13345 13207 13379
rect 13207 13345 13216 13379
rect 13164 13336 13216 13345
rect 14728 13336 14780 13388
rect 15188 13336 15240 13388
rect 15740 13336 15792 13388
rect 17764 13379 17816 13388
rect 17764 13345 17773 13379
rect 17773 13345 17807 13379
rect 17807 13345 17816 13379
rect 17764 13336 17816 13345
rect 20800 13379 20852 13388
rect 20800 13345 20809 13379
rect 20809 13345 20843 13379
rect 20843 13345 20852 13379
rect 20800 13336 20852 13345
rect 21076 13379 21128 13388
rect 21076 13345 21085 13379
rect 21085 13345 21119 13379
rect 21119 13345 21128 13379
rect 21076 13336 21128 13345
rect 21812 13336 21864 13388
rect 22180 13379 22232 13388
rect 22180 13345 22224 13379
rect 22224 13345 22232 13379
rect 24756 13379 24808 13388
rect 22180 13336 22232 13345
rect 24756 13345 24765 13379
rect 24765 13345 24799 13379
rect 24799 13345 24808 13379
rect 24756 13336 24808 13345
rect 13532 13311 13584 13320
rect 13532 13277 13541 13311
rect 13541 13277 13575 13311
rect 13575 13277 13584 13311
rect 13532 13268 13584 13277
rect 15004 13268 15056 13320
rect 18960 13268 19012 13320
rect 23468 13268 23520 13320
rect 18684 13200 18736 13252
rect 13440 13175 13492 13184
rect 13440 13141 13449 13175
rect 13449 13141 13483 13175
rect 13483 13141 13492 13175
rect 13440 13132 13492 13141
rect 13808 13132 13860 13184
rect 14268 13132 14320 13184
rect 5176 13030 5228 13082
rect 5240 13030 5292 13082
rect 5304 13030 5356 13082
rect 5368 13030 5420 13082
rect 14510 13030 14562 13082
rect 14574 13030 14626 13082
rect 14638 13030 14690 13082
rect 14702 13030 14754 13082
rect 23843 13030 23895 13082
rect 23907 13030 23959 13082
rect 23971 13030 24023 13082
rect 24035 13030 24087 13082
rect 13072 12928 13124 12980
rect 13440 12928 13492 12980
rect 13900 12971 13952 12980
rect 13900 12937 13924 12971
rect 13924 12937 13952 12971
rect 13900 12928 13952 12937
rect 14268 12928 14320 12980
rect 14360 12971 14412 12980
rect 14360 12937 14369 12971
rect 14369 12937 14403 12971
rect 14403 12937 14412 12971
rect 14820 12971 14872 12980
rect 14360 12928 14412 12937
rect 14820 12937 14829 12971
rect 14829 12937 14863 12971
rect 14863 12937 14872 12971
rect 14820 12928 14872 12937
rect 15556 12971 15608 12980
rect 15556 12937 15565 12971
rect 15565 12937 15599 12971
rect 15599 12937 15608 12971
rect 15556 12928 15608 12937
rect 17764 12928 17816 12980
rect 18776 12971 18828 12980
rect 18776 12937 18785 12971
rect 18785 12937 18819 12971
rect 18819 12937 18828 12971
rect 18776 12928 18828 12937
rect 21812 12971 21864 12980
rect 21812 12937 21821 12971
rect 21821 12937 21855 12971
rect 21855 12937 21864 12971
rect 21812 12928 21864 12937
rect 23560 12928 23612 12980
rect 24204 12971 24256 12980
rect 24204 12937 24213 12971
rect 24213 12937 24247 12971
rect 24247 12937 24256 12971
rect 24204 12928 24256 12937
rect 24756 12971 24808 12980
rect 24756 12937 24765 12971
rect 24765 12937 24799 12971
rect 24799 12937 24808 12971
rect 24756 12928 24808 12937
rect 14176 12860 14228 12912
rect 12152 12724 12204 12776
rect 13808 12724 13860 12776
rect 13256 12631 13308 12640
rect 13256 12597 13265 12631
rect 13265 12597 13299 12631
rect 13299 12597 13308 12631
rect 13532 12631 13584 12640
rect 13256 12588 13308 12597
rect 13532 12597 13541 12631
rect 13541 12597 13575 12631
rect 13575 12597 13584 12631
rect 15464 12792 15516 12844
rect 19512 12792 19564 12844
rect 17488 12724 17540 12776
rect 20524 12724 20576 12776
rect 21444 12860 21496 12912
rect 21352 12835 21404 12844
rect 21352 12801 21361 12835
rect 21361 12801 21395 12835
rect 21395 12801 21404 12835
rect 21352 12792 21404 12801
rect 23468 12792 23520 12844
rect 21168 12724 21220 12776
rect 24204 12724 24256 12776
rect 15556 12656 15608 12708
rect 16108 12656 16160 12708
rect 18316 12699 18368 12708
rect 18316 12665 18325 12699
rect 18325 12665 18359 12699
rect 18359 12665 18368 12699
rect 18316 12656 18368 12665
rect 19972 12699 20024 12708
rect 13532 12588 13584 12597
rect 18960 12588 19012 12640
rect 19972 12665 19981 12699
rect 19981 12665 20015 12699
rect 20015 12665 20024 12699
rect 22180 12699 22232 12708
rect 19972 12656 20024 12665
rect 22180 12665 22189 12699
rect 22189 12665 22223 12699
rect 22223 12665 22232 12699
rect 22180 12656 22232 12665
rect 20524 12588 20576 12640
rect 20800 12588 20852 12640
rect 23376 12588 23428 12640
rect 9843 12486 9895 12538
rect 9907 12486 9959 12538
rect 9971 12486 10023 12538
rect 10035 12486 10087 12538
rect 19176 12486 19228 12538
rect 19240 12486 19292 12538
rect 19304 12486 19356 12538
rect 19368 12486 19420 12538
rect 13256 12384 13308 12436
rect 14176 12427 14228 12436
rect 14176 12393 14185 12427
rect 14185 12393 14219 12427
rect 14219 12393 14228 12427
rect 14176 12384 14228 12393
rect 14912 12384 14964 12436
rect 15740 12316 15792 12368
rect 17488 12359 17540 12368
rect 17488 12325 17497 12359
rect 17497 12325 17531 12359
rect 17531 12325 17540 12359
rect 17488 12316 17540 12325
rect 19512 12316 19564 12368
rect 12704 12291 12756 12300
rect 12704 12257 12713 12291
rect 12713 12257 12747 12291
rect 12747 12257 12756 12291
rect 12704 12248 12756 12257
rect 13716 12291 13768 12300
rect 13716 12257 13725 12291
rect 13725 12257 13759 12291
rect 13759 12257 13768 12291
rect 13716 12248 13768 12257
rect 14176 12248 14228 12300
rect 14820 12291 14872 12300
rect 14820 12257 14829 12291
rect 14829 12257 14863 12291
rect 14863 12257 14872 12291
rect 14820 12248 14872 12257
rect 20800 12291 20852 12300
rect 20800 12257 20809 12291
rect 20809 12257 20843 12291
rect 20843 12257 20852 12291
rect 20800 12248 20852 12257
rect 13992 12180 14044 12232
rect 17396 12223 17448 12232
rect 17396 12189 17405 12223
rect 17405 12189 17439 12223
rect 17439 12189 17448 12223
rect 17396 12180 17448 12189
rect 18500 12180 18552 12232
rect 20616 12180 20668 12232
rect 21168 12248 21220 12300
rect 22916 12291 22968 12300
rect 22916 12257 22925 12291
rect 22925 12257 22959 12291
rect 22959 12257 22968 12291
rect 22916 12248 22968 12257
rect 21260 12223 21312 12232
rect 21260 12189 21269 12223
rect 21269 12189 21303 12223
rect 21303 12189 21312 12223
rect 21260 12180 21312 12189
rect 23468 12223 23520 12232
rect 23468 12189 23477 12223
rect 23477 12189 23511 12223
rect 23511 12189 23520 12223
rect 23468 12180 23520 12189
rect 13164 12112 13216 12164
rect 14084 12044 14136 12096
rect 14360 12044 14412 12096
rect 15372 12044 15424 12096
rect 18776 12087 18828 12096
rect 18776 12053 18785 12087
rect 18785 12053 18819 12087
rect 18819 12053 18828 12087
rect 18776 12044 18828 12053
rect 5176 11942 5228 11994
rect 5240 11942 5292 11994
rect 5304 11942 5356 11994
rect 5368 11942 5420 11994
rect 14510 11942 14562 11994
rect 14574 11942 14626 11994
rect 14638 11942 14690 11994
rect 14702 11942 14754 11994
rect 23843 11942 23895 11994
rect 23907 11942 23959 11994
rect 23971 11942 24023 11994
rect 24035 11942 24087 11994
rect 13072 11883 13124 11892
rect 13072 11849 13081 11883
rect 13081 11849 13115 11883
rect 13115 11849 13124 11883
rect 13072 11840 13124 11849
rect 14820 11840 14872 11892
rect 17488 11840 17540 11892
rect 20800 11840 20852 11892
rect 21536 11840 21588 11892
rect 22916 11883 22968 11892
rect 22916 11849 22925 11883
rect 22925 11849 22959 11883
rect 22959 11849 22968 11883
rect 22916 11840 22968 11849
rect 12520 11772 12572 11824
rect 14360 11772 14412 11824
rect 16108 11772 16160 11824
rect 16752 11772 16804 11824
rect 19972 11815 20024 11824
rect 12704 11704 12756 11756
rect 14268 11747 14320 11756
rect 14268 11713 14277 11747
rect 14277 11713 14311 11747
rect 14311 11713 14320 11747
rect 14268 11704 14320 11713
rect 13992 11636 14044 11688
rect 13624 11568 13676 11620
rect 13808 11568 13860 11620
rect 13716 11543 13768 11552
rect 13716 11509 13725 11543
rect 13725 11509 13759 11543
rect 13759 11509 13768 11543
rect 13716 11500 13768 11509
rect 14360 11500 14412 11552
rect 15188 11500 15240 11552
rect 15648 11679 15700 11688
rect 15648 11645 15654 11679
rect 15654 11645 15700 11679
rect 15648 11636 15700 11645
rect 15372 11568 15424 11620
rect 16200 11611 16252 11620
rect 16200 11577 16209 11611
rect 16209 11577 16243 11611
rect 16243 11577 16252 11611
rect 16200 11568 16252 11577
rect 19972 11781 19981 11815
rect 19981 11781 20015 11815
rect 20015 11781 20024 11815
rect 19972 11772 20024 11781
rect 18500 11704 18552 11756
rect 21352 11747 21404 11756
rect 21352 11713 21361 11747
rect 21361 11713 21395 11747
rect 21395 11713 21404 11747
rect 21352 11704 21404 11713
rect 17580 11679 17632 11688
rect 17580 11645 17589 11679
rect 17589 11645 17623 11679
rect 17623 11645 17632 11679
rect 17580 11636 17632 11645
rect 18592 11500 18644 11552
rect 21536 11568 21588 11620
rect 23284 11611 23336 11620
rect 23284 11577 23293 11611
rect 23293 11577 23327 11611
rect 23327 11577 23336 11611
rect 23284 11568 23336 11577
rect 22916 11500 22968 11552
rect 24204 11568 24256 11620
rect 9843 11398 9895 11450
rect 9907 11398 9959 11450
rect 9971 11398 10023 11450
rect 10035 11398 10087 11450
rect 19176 11398 19228 11450
rect 19240 11398 19292 11450
rect 19304 11398 19356 11450
rect 19368 11398 19420 11450
rect 12520 11296 12572 11348
rect 14084 11296 14136 11348
rect 14820 11296 14872 11348
rect 17488 11296 17540 11348
rect 21352 11339 21404 11348
rect 21352 11305 21361 11339
rect 21361 11305 21395 11339
rect 21395 11305 21404 11339
rect 21352 11296 21404 11305
rect 23284 11339 23336 11348
rect 23284 11305 23293 11339
rect 23293 11305 23327 11339
rect 23327 11305 23336 11339
rect 23284 11296 23336 11305
rect 13992 11228 14044 11280
rect 15648 11228 15700 11280
rect 16752 11271 16804 11280
rect 16752 11237 16755 11271
rect 16755 11237 16789 11271
rect 16789 11237 16804 11271
rect 16752 11228 16804 11237
rect 17396 11228 17448 11280
rect 18316 11271 18368 11280
rect 18316 11237 18325 11271
rect 18325 11237 18359 11271
rect 18359 11237 18368 11271
rect 18316 11228 18368 11237
rect 20616 11271 20668 11280
rect 20616 11237 20625 11271
rect 20625 11237 20659 11271
rect 20659 11237 20668 11271
rect 20616 11228 20668 11237
rect 21536 11228 21588 11280
rect 21812 11228 21864 11280
rect 23468 11228 23520 11280
rect 24388 11228 24440 11280
rect 12520 11203 12572 11212
rect 12520 11169 12529 11203
rect 12529 11169 12563 11203
rect 12563 11169 12572 11203
rect 12520 11160 12572 11169
rect 14084 11160 14136 11212
rect 14820 11203 14872 11212
rect 14820 11169 14829 11203
rect 14829 11169 14863 11203
rect 14863 11169 14872 11203
rect 14820 11160 14872 11169
rect 15280 11203 15332 11212
rect 15280 11169 15289 11203
rect 15289 11169 15323 11203
rect 15323 11169 15332 11203
rect 15280 11160 15332 11169
rect 21260 11160 21312 11212
rect 13808 11092 13860 11144
rect 16384 11135 16436 11144
rect 16384 11101 16393 11135
rect 16393 11101 16427 11135
rect 16427 11101 16436 11135
rect 16384 11092 16436 11101
rect 17948 11092 18000 11144
rect 18500 11135 18552 11144
rect 18500 11101 18509 11135
rect 18509 11101 18543 11135
rect 18543 11101 18552 11135
rect 22548 11160 22600 11212
rect 18500 11092 18552 11101
rect 23468 11092 23520 11144
rect 13532 11024 13584 11076
rect 14268 11024 14320 11076
rect 15188 11024 15240 11076
rect 17580 11067 17632 11076
rect 16568 10956 16620 11008
rect 17580 11033 17589 11067
rect 17589 11033 17623 11067
rect 17623 11033 17632 11067
rect 17580 11024 17632 11033
rect 24204 11067 24256 11076
rect 24204 11033 24213 11067
rect 24213 11033 24247 11067
rect 24247 11033 24256 11067
rect 24204 11024 24256 11033
rect 23008 10956 23060 11008
rect 24756 10956 24808 11008
rect 5176 10854 5228 10906
rect 5240 10854 5292 10906
rect 5304 10854 5356 10906
rect 5368 10854 5420 10906
rect 14510 10854 14562 10906
rect 14574 10854 14626 10906
rect 14638 10854 14690 10906
rect 14702 10854 14754 10906
rect 23843 10854 23895 10906
rect 23907 10854 23959 10906
rect 23971 10854 24023 10906
rect 24035 10854 24087 10906
rect 12520 10795 12572 10804
rect 12520 10761 12529 10795
rect 12529 10761 12563 10795
rect 12563 10761 12572 10795
rect 13348 10795 13400 10804
rect 12520 10752 12572 10761
rect 13348 10761 13357 10795
rect 13357 10761 13391 10795
rect 13391 10761 13400 10795
rect 13348 10752 13400 10761
rect 14084 10795 14136 10804
rect 14084 10761 14093 10795
rect 14093 10761 14127 10795
rect 14127 10761 14136 10795
rect 14084 10752 14136 10761
rect 15004 10752 15056 10804
rect 15740 10795 15792 10804
rect 15740 10761 15749 10795
rect 15749 10761 15783 10795
rect 15783 10761 15792 10795
rect 15740 10752 15792 10761
rect 16384 10752 16436 10804
rect 18316 10752 18368 10804
rect 18592 10795 18644 10804
rect 18592 10761 18601 10795
rect 18601 10761 18635 10795
rect 18635 10761 18644 10795
rect 18592 10752 18644 10761
rect 18960 10795 19012 10804
rect 18960 10761 18969 10795
rect 18969 10761 19003 10795
rect 19003 10761 19012 10795
rect 18960 10752 19012 10761
rect 22548 10795 22600 10804
rect 22548 10761 22557 10795
rect 22557 10761 22591 10795
rect 22591 10761 22600 10795
rect 22548 10752 22600 10761
rect 24388 10795 24440 10804
rect 24388 10761 24397 10795
rect 24397 10761 24431 10795
rect 24431 10761 24440 10795
rect 24388 10752 24440 10761
rect 24756 10795 24808 10804
rect 24756 10761 24765 10795
rect 24765 10761 24799 10795
rect 24799 10761 24808 10795
rect 24756 10752 24808 10761
rect 25124 10795 25176 10804
rect 25124 10761 25133 10795
rect 25133 10761 25167 10795
rect 25167 10761 25176 10795
rect 25124 10752 25176 10761
rect 16752 10684 16804 10736
rect 16568 10659 16620 10668
rect 16568 10625 16577 10659
rect 16577 10625 16611 10659
rect 16611 10625 16620 10659
rect 16568 10616 16620 10625
rect 19696 10659 19748 10668
rect 19696 10625 19705 10659
rect 19705 10625 19739 10659
rect 19739 10625 19748 10659
rect 19696 10616 19748 10625
rect 13900 10548 13952 10600
rect 15188 10548 15240 10600
rect 15740 10548 15792 10600
rect 16292 10591 16344 10600
rect 16292 10557 16301 10591
rect 16301 10557 16335 10591
rect 16335 10557 16344 10591
rect 16292 10548 16344 10557
rect 18592 10548 18644 10600
rect 20800 10616 20852 10668
rect 24204 10616 24256 10668
rect 24940 10591 24992 10600
rect 24940 10557 24949 10591
rect 24949 10557 24983 10591
rect 24983 10557 24992 10591
rect 24940 10548 24992 10557
rect 20892 10480 20944 10532
rect 21536 10480 21588 10532
rect 13624 10412 13676 10464
rect 14636 10412 14688 10464
rect 17948 10412 18000 10464
rect 21812 10455 21864 10464
rect 21812 10421 21821 10455
rect 21821 10421 21855 10455
rect 21855 10421 21864 10455
rect 21812 10412 21864 10421
rect 22088 10455 22140 10464
rect 22088 10421 22097 10455
rect 22097 10421 22131 10455
rect 22131 10421 22140 10455
rect 22088 10412 22140 10421
rect 23008 10455 23060 10464
rect 23008 10421 23017 10455
rect 23017 10421 23051 10455
rect 23051 10421 23060 10455
rect 23008 10412 23060 10421
rect 23284 10412 23336 10464
rect 23928 10480 23980 10532
rect 9843 10310 9895 10362
rect 9907 10310 9959 10362
rect 9971 10310 10023 10362
rect 10035 10310 10087 10362
rect 19176 10310 19228 10362
rect 19240 10310 19292 10362
rect 19304 10310 19356 10362
rect 19368 10310 19420 10362
rect 14084 10208 14136 10260
rect 16292 10251 16344 10260
rect 13900 10183 13952 10192
rect 13900 10149 13909 10183
rect 13909 10149 13943 10183
rect 13943 10149 13952 10183
rect 13900 10140 13952 10149
rect 13532 10115 13584 10124
rect 13532 10081 13541 10115
rect 13541 10081 13575 10115
rect 13575 10081 13584 10115
rect 13532 10072 13584 10081
rect 16292 10217 16301 10251
rect 16301 10217 16335 10251
rect 16335 10217 16344 10251
rect 16292 10208 16344 10217
rect 20708 10251 20760 10260
rect 20708 10217 20717 10251
rect 20717 10217 20751 10251
rect 20751 10217 20760 10251
rect 20708 10208 20760 10217
rect 22916 10208 22968 10260
rect 24204 10208 24256 10260
rect 23652 10140 23704 10192
rect 14820 10115 14872 10124
rect 14820 10081 14829 10115
rect 14829 10081 14863 10115
rect 14863 10081 14872 10115
rect 14820 10072 14872 10081
rect 18868 10115 18920 10124
rect 18868 10081 18877 10115
rect 18877 10081 18911 10115
rect 18911 10081 18920 10115
rect 18868 10072 18920 10081
rect 20524 10115 20576 10124
rect 20524 10081 20533 10115
rect 20533 10081 20567 10115
rect 20567 10081 20576 10115
rect 20524 10072 20576 10081
rect 20892 10115 20944 10124
rect 20892 10081 20901 10115
rect 20901 10081 20935 10115
rect 20935 10081 20944 10115
rect 20892 10072 20944 10081
rect 22640 10115 22692 10124
rect 22640 10081 22658 10115
rect 22658 10081 22692 10115
rect 22640 10072 22692 10081
rect 15188 10047 15240 10056
rect 15188 10013 15197 10047
rect 15197 10013 15231 10047
rect 15231 10013 15240 10047
rect 15188 10004 15240 10013
rect 22916 10004 22968 10056
rect 23928 10047 23980 10056
rect 23928 10013 23937 10047
rect 23937 10013 23971 10047
rect 23971 10013 23980 10047
rect 23928 10004 23980 10013
rect 15280 9979 15332 9988
rect 15280 9945 15289 9979
rect 15289 9945 15323 9979
rect 15323 9945 15332 9979
rect 15280 9936 15332 9945
rect 16292 9936 16344 9988
rect 22640 9936 22692 9988
rect 13348 9868 13400 9920
rect 15556 9868 15608 9920
rect 15832 9911 15884 9920
rect 15832 9877 15841 9911
rect 15841 9877 15875 9911
rect 15875 9877 15884 9911
rect 15832 9868 15884 9877
rect 18960 9911 19012 9920
rect 18960 9877 18969 9911
rect 18969 9877 19003 9911
rect 19003 9877 19012 9911
rect 18960 9868 19012 9877
rect 23284 9911 23336 9920
rect 23284 9877 23293 9911
rect 23293 9877 23327 9911
rect 23327 9877 23336 9911
rect 23284 9868 23336 9877
rect 5176 9766 5228 9818
rect 5240 9766 5292 9818
rect 5304 9766 5356 9818
rect 5368 9766 5420 9818
rect 14510 9766 14562 9818
rect 14574 9766 14626 9818
rect 14638 9766 14690 9818
rect 14702 9766 14754 9818
rect 23843 9766 23895 9818
rect 23907 9766 23959 9818
rect 23971 9766 24023 9818
rect 24035 9766 24087 9818
rect 12612 9707 12664 9716
rect 12612 9673 12621 9707
rect 12621 9673 12655 9707
rect 12655 9673 12664 9707
rect 12612 9664 12664 9673
rect 15188 9664 15240 9716
rect 15556 9639 15608 9648
rect 15556 9605 15565 9639
rect 15565 9605 15599 9639
rect 15599 9605 15608 9639
rect 15556 9596 15608 9605
rect 14084 9571 14136 9580
rect 14084 9537 14093 9571
rect 14093 9537 14127 9571
rect 14127 9537 14136 9571
rect 20892 9664 20944 9716
rect 22088 9664 22140 9716
rect 22916 9707 22968 9716
rect 22916 9673 22925 9707
rect 22925 9673 22959 9707
rect 22959 9673 22968 9707
rect 22916 9664 22968 9673
rect 24204 9664 24256 9716
rect 25768 9664 25820 9716
rect 15832 9596 15884 9648
rect 18868 9596 18920 9648
rect 24388 9596 24440 9648
rect 14084 9528 14136 9537
rect 13716 9503 13768 9512
rect 12336 9435 12388 9444
rect 12336 9401 12345 9435
rect 12345 9401 12379 9435
rect 12379 9401 12388 9435
rect 12336 9392 12388 9401
rect 13716 9469 13725 9503
rect 13725 9469 13759 9503
rect 13759 9469 13768 9503
rect 13716 9460 13768 9469
rect 14268 9503 14320 9512
rect 14268 9469 14277 9503
rect 14277 9469 14311 9503
rect 14311 9469 14320 9503
rect 14268 9460 14320 9469
rect 14820 9503 14872 9512
rect 14820 9469 14829 9503
rect 14829 9469 14863 9503
rect 14863 9469 14872 9503
rect 20524 9528 20576 9580
rect 23744 9528 23796 9580
rect 14820 9460 14872 9469
rect 22088 9503 22140 9512
rect 22088 9469 22132 9503
rect 22132 9469 22140 9503
rect 22088 9460 22140 9469
rect 23284 9503 23336 9512
rect 23284 9469 23293 9503
rect 23293 9469 23327 9503
rect 23327 9469 23336 9503
rect 23284 9460 23336 9469
rect 13532 9324 13584 9376
rect 15096 9367 15148 9376
rect 15096 9333 15105 9367
rect 15105 9333 15139 9367
rect 15139 9333 15148 9367
rect 15372 9392 15424 9444
rect 18776 9392 18828 9444
rect 15924 9367 15976 9376
rect 15096 9324 15148 9333
rect 15924 9333 15933 9367
rect 15933 9333 15967 9367
rect 15967 9333 15976 9367
rect 15924 9324 15976 9333
rect 18868 9324 18920 9376
rect 19696 9392 19748 9444
rect 20432 9367 20484 9376
rect 20432 9333 20441 9367
rect 20441 9333 20475 9367
rect 20475 9333 20484 9367
rect 20432 9324 20484 9333
rect 9843 9222 9895 9274
rect 9907 9222 9959 9274
rect 9971 9222 10023 9274
rect 10035 9222 10087 9274
rect 19176 9222 19228 9274
rect 19240 9222 19292 9274
rect 19304 9222 19356 9274
rect 19368 9222 19420 9274
rect 14176 9120 14228 9172
rect 15188 9120 15240 9172
rect 19512 9120 19564 9172
rect 20432 9120 20484 9172
rect 21536 9120 21588 9172
rect 22640 9163 22692 9172
rect 22640 9129 22649 9163
rect 22649 9129 22683 9163
rect 22683 9129 22692 9163
rect 22640 9120 22692 9129
rect 24664 9163 24716 9172
rect 24664 9129 24673 9163
rect 24673 9129 24707 9163
rect 24707 9129 24716 9163
rect 24664 9120 24716 9129
rect 12336 9052 12388 9104
rect 14360 9052 14412 9104
rect 16752 9052 16804 9104
rect 17672 9052 17724 9104
rect 21260 9052 21312 9104
rect 21812 9052 21864 9104
rect 23100 9095 23152 9104
rect 23100 9061 23109 9095
rect 23109 9061 23143 9095
rect 23143 9061 23152 9095
rect 23100 9052 23152 9061
rect 13256 8984 13308 9036
rect 13716 8984 13768 9036
rect 14912 8984 14964 9036
rect 15464 8984 15516 9036
rect 15924 8984 15976 9036
rect 16384 8984 16436 9036
rect 20708 9027 20760 9036
rect 20708 8993 20717 9027
rect 20717 8993 20751 9027
rect 20751 8993 20760 9027
rect 20708 8984 20760 8993
rect 24388 8984 24440 9036
rect 13532 8959 13584 8968
rect 13532 8925 13541 8959
rect 13541 8925 13575 8959
rect 13575 8925 13584 8959
rect 13532 8916 13584 8925
rect 16568 8959 16620 8968
rect 16568 8925 16577 8959
rect 16577 8925 16611 8959
rect 16611 8925 16620 8959
rect 16568 8916 16620 8925
rect 18408 8959 18460 8968
rect 18408 8925 18417 8959
rect 18417 8925 18451 8959
rect 18451 8925 18460 8959
rect 18408 8916 18460 8925
rect 18776 8959 18828 8968
rect 18776 8925 18785 8959
rect 18785 8925 18819 8959
rect 18819 8925 18828 8959
rect 18776 8916 18828 8925
rect 23008 8959 23060 8968
rect 23008 8925 23017 8959
rect 23017 8925 23051 8959
rect 23051 8925 23060 8959
rect 23008 8916 23060 8925
rect 12888 8848 12940 8900
rect 14268 8848 14320 8900
rect 23560 8891 23612 8900
rect 23560 8857 23569 8891
rect 23569 8857 23603 8891
rect 23603 8857 23612 8891
rect 23560 8848 23612 8857
rect 13624 8780 13676 8832
rect 16384 8823 16436 8832
rect 16384 8789 16393 8823
rect 16393 8789 16427 8823
rect 16427 8789 16436 8823
rect 16384 8780 16436 8789
rect 17672 8780 17724 8832
rect 21628 8823 21680 8832
rect 21628 8789 21637 8823
rect 21637 8789 21671 8823
rect 21671 8789 21680 8823
rect 21628 8780 21680 8789
rect 23284 8780 23336 8832
rect 5176 8678 5228 8730
rect 5240 8678 5292 8730
rect 5304 8678 5356 8730
rect 5368 8678 5420 8730
rect 14510 8678 14562 8730
rect 14574 8678 14626 8730
rect 14638 8678 14690 8730
rect 14702 8678 14754 8730
rect 23843 8678 23895 8730
rect 23907 8678 23959 8730
rect 23971 8678 24023 8730
rect 24035 8678 24087 8730
rect 12888 8619 12940 8628
rect 12888 8585 12897 8619
rect 12897 8585 12931 8619
rect 12931 8585 12940 8619
rect 12888 8576 12940 8585
rect 13532 8576 13584 8628
rect 15280 8576 15332 8628
rect 15464 8619 15516 8628
rect 15464 8585 15473 8619
rect 15473 8585 15507 8619
rect 15507 8585 15516 8619
rect 15464 8576 15516 8585
rect 15740 8619 15792 8628
rect 15740 8585 15749 8619
rect 15749 8585 15783 8619
rect 15783 8585 15792 8619
rect 15740 8576 15792 8585
rect 16752 8576 16804 8628
rect 13624 8440 13676 8492
rect 18868 8576 18920 8628
rect 18960 8576 19012 8628
rect 14360 8415 14412 8424
rect 14360 8381 14369 8415
rect 14369 8381 14403 8415
rect 14403 8381 14412 8415
rect 14360 8372 14412 8381
rect 14912 8372 14964 8424
rect 15740 8372 15792 8424
rect 16200 8372 16252 8424
rect 16384 8415 16436 8424
rect 16384 8381 16393 8415
rect 16393 8381 16427 8415
rect 16427 8381 16436 8415
rect 16384 8372 16436 8381
rect 17580 8415 17632 8424
rect 17580 8381 17589 8415
rect 17589 8381 17623 8415
rect 17623 8381 17632 8415
rect 17580 8372 17632 8381
rect 13256 8304 13308 8356
rect 13808 8236 13860 8288
rect 15096 8304 15148 8356
rect 17764 8304 17816 8356
rect 20708 8576 20760 8628
rect 21260 8619 21312 8628
rect 21260 8585 21269 8619
rect 21269 8585 21303 8619
rect 21303 8585 21312 8619
rect 21260 8576 21312 8585
rect 22824 8576 22876 8628
rect 23008 8576 23060 8628
rect 24940 8619 24992 8628
rect 24940 8585 24949 8619
rect 24949 8585 24983 8619
rect 24983 8585 24992 8619
rect 24940 8576 24992 8585
rect 19512 8440 19564 8492
rect 19696 8483 19748 8492
rect 19696 8449 19705 8483
rect 19705 8449 19739 8483
rect 19739 8449 19748 8483
rect 19696 8440 19748 8449
rect 21536 8440 21588 8492
rect 23284 8483 23336 8492
rect 23284 8449 23293 8483
rect 23293 8449 23327 8483
rect 23327 8449 23336 8483
rect 23284 8440 23336 8449
rect 23560 8483 23612 8492
rect 23560 8449 23569 8483
rect 23569 8449 23603 8483
rect 23603 8449 23612 8483
rect 23560 8440 23612 8449
rect 24756 8415 24808 8424
rect 21260 8304 21312 8356
rect 24756 8381 24765 8415
rect 24765 8381 24799 8415
rect 24799 8381 24808 8415
rect 24756 8372 24808 8381
rect 23376 8347 23428 8356
rect 23376 8313 23385 8347
rect 23385 8313 23419 8347
rect 23419 8313 23428 8347
rect 23376 8304 23428 8313
rect 24388 8304 24440 8356
rect 17672 8236 17724 8288
rect 23100 8236 23152 8288
rect 9843 8134 9895 8186
rect 9907 8134 9959 8186
rect 9971 8134 10023 8186
rect 10035 8134 10087 8186
rect 19176 8134 19228 8186
rect 19240 8134 19292 8186
rect 19304 8134 19356 8186
rect 19368 8134 19420 8186
rect 13256 8075 13308 8084
rect 13256 8041 13265 8075
rect 13265 8041 13299 8075
rect 13299 8041 13308 8075
rect 13256 8032 13308 8041
rect 14360 8032 14412 8084
rect 16568 8032 16620 8084
rect 17580 8075 17632 8084
rect 17580 8041 17589 8075
rect 17589 8041 17623 8075
rect 17623 8041 17632 8075
rect 17580 8032 17632 8041
rect 18408 8032 18460 8084
rect 24664 8032 24716 8084
rect 15004 7964 15056 8016
rect 18592 8007 18644 8016
rect 18592 7973 18601 8007
rect 18601 7973 18635 8007
rect 18635 7973 18644 8007
rect 18592 7964 18644 7973
rect 21628 8007 21680 8016
rect 21628 7973 21637 8007
rect 21637 7973 21671 8007
rect 21671 7973 21680 8007
rect 23192 8007 23244 8016
rect 21628 7964 21680 7973
rect 23192 7973 23201 8007
rect 23201 7973 23235 8007
rect 23235 7973 23244 8007
rect 23192 7964 23244 7973
rect 16108 7939 16160 7948
rect 16108 7905 16117 7939
rect 16117 7905 16151 7939
rect 16151 7905 16160 7939
rect 16476 7939 16528 7948
rect 16108 7896 16160 7905
rect 16476 7905 16485 7939
rect 16485 7905 16519 7939
rect 16519 7905 16528 7939
rect 16476 7896 16528 7905
rect 24572 7939 24624 7948
rect 24572 7905 24581 7939
rect 24581 7905 24615 7939
rect 24615 7905 24624 7939
rect 24572 7896 24624 7905
rect 17488 7828 17540 7880
rect 18500 7871 18552 7880
rect 18500 7837 18509 7871
rect 18509 7837 18543 7871
rect 18543 7837 18552 7871
rect 18500 7828 18552 7837
rect 18868 7871 18920 7880
rect 18868 7837 18877 7871
rect 18877 7837 18911 7871
rect 18911 7837 18920 7871
rect 18868 7828 18920 7837
rect 20984 7828 21036 7880
rect 23100 7871 23152 7880
rect 23100 7837 23109 7871
rect 23109 7837 23143 7871
rect 23143 7837 23152 7871
rect 23100 7828 23152 7837
rect 23284 7828 23336 7880
rect 15372 7735 15424 7744
rect 15372 7701 15381 7735
rect 15381 7701 15415 7735
rect 15415 7701 15424 7735
rect 15372 7692 15424 7701
rect 15556 7692 15608 7744
rect 5176 7590 5228 7642
rect 5240 7590 5292 7642
rect 5304 7590 5356 7642
rect 5368 7590 5420 7642
rect 14510 7590 14562 7642
rect 14574 7590 14626 7642
rect 14638 7590 14690 7642
rect 14702 7590 14754 7642
rect 23843 7590 23895 7642
rect 23907 7590 23959 7642
rect 23971 7590 24023 7642
rect 24035 7590 24087 7642
rect 13624 7420 13676 7472
rect 16108 7488 16160 7540
rect 20984 7531 21036 7540
rect 20984 7497 20993 7531
rect 20993 7497 21027 7531
rect 21027 7497 21036 7531
rect 20984 7488 21036 7497
rect 21628 7488 21680 7540
rect 23192 7488 23244 7540
rect 24204 7488 24256 7540
rect 15004 7420 15056 7472
rect 15556 7463 15608 7472
rect 15556 7429 15580 7463
rect 15580 7429 15608 7463
rect 15556 7420 15608 7429
rect 12244 7327 12296 7336
rect 12244 7293 12253 7327
rect 12253 7293 12287 7327
rect 12287 7293 12296 7327
rect 12244 7284 12296 7293
rect 12060 7259 12112 7268
rect 12060 7225 12069 7259
rect 12069 7225 12103 7259
rect 12103 7225 12112 7259
rect 12060 7216 12112 7225
rect 18592 7352 18644 7404
rect 23008 7352 23060 7404
rect 14084 7284 14136 7336
rect 15556 7284 15608 7336
rect 17672 7284 17724 7336
rect 21628 7327 21680 7336
rect 21628 7293 21637 7327
rect 21637 7293 21671 7327
rect 21671 7293 21680 7327
rect 23376 7327 23428 7336
rect 21628 7284 21680 7293
rect 23376 7293 23385 7327
rect 23385 7293 23419 7327
rect 23419 7293 23428 7327
rect 23376 7284 23428 7293
rect 24480 7284 24532 7336
rect 13808 7259 13860 7268
rect 13808 7225 13817 7259
rect 13817 7225 13851 7259
rect 13851 7225 13860 7259
rect 13808 7216 13860 7225
rect 15372 7259 15424 7268
rect 15372 7225 15381 7259
rect 15381 7225 15415 7259
rect 15415 7225 15424 7259
rect 15372 7216 15424 7225
rect 13624 7191 13676 7200
rect 13624 7157 13633 7191
rect 13633 7157 13667 7191
rect 13667 7157 13676 7191
rect 13624 7148 13676 7157
rect 14360 7148 14412 7200
rect 23100 7216 23152 7268
rect 24388 7216 24440 7268
rect 16476 7148 16528 7200
rect 16936 7148 16988 7200
rect 18500 7148 18552 7200
rect 19604 7148 19656 7200
rect 20248 7148 20300 7200
rect 24204 7148 24256 7200
rect 24572 7191 24624 7200
rect 24572 7157 24581 7191
rect 24581 7157 24615 7191
rect 24615 7157 24624 7191
rect 24572 7148 24624 7157
rect 9843 7046 9895 7098
rect 9907 7046 9959 7098
rect 9971 7046 10023 7098
rect 10035 7046 10087 7098
rect 19176 7046 19228 7098
rect 19240 7046 19292 7098
rect 19304 7046 19356 7098
rect 19368 7046 19420 7098
rect 11876 6851 11928 6860
rect 11876 6817 11885 6851
rect 11885 6817 11919 6851
rect 11919 6817 11928 6851
rect 11876 6808 11928 6817
rect 11600 6740 11652 6792
rect 12244 6808 12296 6860
rect 15372 6944 15424 6996
rect 21628 6987 21680 6996
rect 21628 6953 21637 6987
rect 21637 6953 21671 6987
rect 21671 6953 21680 6987
rect 23376 6987 23428 6996
rect 21628 6944 21680 6953
rect 23376 6953 23385 6987
rect 23385 6953 23419 6987
rect 23419 6953 23428 6987
rect 23376 6944 23428 6953
rect 14084 6876 14136 6928
rect 17120 6919 17172 6928
rect 17120 6885 17129 6919
rect 17129 6885 17163 6919
rect 17163 6885 17172 6919
rect 17120 6876 17172 6885
rect 18868 6919 18920 6928
rect 18868 6885 18877 6919
rect 18877 6885 18911 6919
rect 18911 6885 18920 6919
rect 18868 6876 18920 6885
rect 13440 6851 13492 6860
rect 13440 6817 13449 6851
rect 13449 6817 13483 6851
rect 13483 6817 13492 6851
rect 13440 6808 13492 6817
rect 14360 6808 14412 6860
rect 15096 6851 15148 6860
rect 15096 6817 15105 6851
rect 15105 6817 15139 6851
rect 15139 6817 15148 6851
rect 15096 6808 15148 6817
rect 15188 6808 15240 6860
rect 16200 6808 16252 6860
rect 16568 6851 16620 6860
rect 16568 6817 16577 6851
rect 16577 6817 16611 6851
rect 16611 6817 16620 6851
rect 16568 6808 16620 6817
rect 16936 6851 16988 6860
rect 16936 6817 16945 6851
rect 16945 6817 16979 6851
rect 16979 6817 16988 6851
rect 16936 6808 16988 6817
rect 18500 6851 18552 6860
rect 18500 6817 18509 6851
rect 18509 6817 18543 6851
rect 18543 6817 18552 6851
rect 18500 6808 18552 6817
rect 21076 6851 21128 6860
rect 21076 6817 21085 6851
rect 21085 6817 21119 6851
rect 21119 6817 21128 6851
rect 21076 6808 21128 6817
rect 22824 6851 22876 6860
rect 22824 6817 22833 6851
rect 22833 6817 22867 6851
rect 22867 6817 22876 6851
rect 22824 6808 22876 6817
rect 23560 6808 23612 6860
rect 24296 6808 24348 6860
rect 25124 6808 25176 6860
rect 13900 6783 13952 6792
rect 13900 6749 13909 6783
rect 13909 6749 13943 6783
rect 13943 6749 13952 6783
rect 13900 6740 13952 6749
rect 15372 6740 15424 6792
rect 19880 6740 19932 6792
rect 24388 6672 24440 6724
rect 20892 6647 20944 6656
rect 20892 6613 20901 6647
rect 20901 6613 20935 6647
rect 20935 6613 20944 6647
rect 20892 6604 20944 6613
rect 5176 6502 5228 6554
rect 5240 6502 5292 6554
rect 5304 6502 5356 6554
rect 5368 6502 5420 6554
rect 14510 6502 14562 6554
rect 14574 6502 14626 6554
rect 14638 6502 14690 6554
rect 14702 6502 14754 6554
rect 23843 6502 23895 6554
rect 23907 6502 23959 6554
rect 23971 6502 24023 6554
rect 24035 6502 24087 6554
rect 12060 6400 12112 6452
rect 13440 6400 13492 6452
rect 15096 6400 15148 6452
rect 16568 6443 16620 6452
rect 16568 6409 16577 6443
rect 16577 6409 16611 6443
rect 16611 6409 16620 6443
rect 16568 6400 16620 6409
rect 16936 6443 16988 6452
rect 16936 6409 16945 6443
rect 16945 6409 16979 6443
rect 16979 6409 16988 6443
rect 16936 6400 16988 6409
rect 18868 6443 18920 6452
rect 18868 6409 18877 6443
rect 18877 6409 18911 6443
rect 18911 6409 18920 6443
rect 18868 6400 18920 6409
rect 20248 6400 20300 6452
rect 20892 6443 20944 6452
rect 14360 6332 14412 6384
rect 15188 6332 15240 6384
rect 20892 6409 20901 6443
rect 20901 6409 20935 6443
rect 20935 6409 20944 6443
rect 20892 6400 20944 6409
rect 21076 6400 21128 6452
rect 23560 6400 23612 6452
rect 24756 6443 24808 6452
rect 24756 6409 24765 6443
rect 24765 6409 24799 6443
rect 24799 6409 24808 6443
rect 24756 6400 24808 6409
rect 20800 6332 20852 6384
rect 15372 6307 15424 6316
rect 15372 6273 15381 6307
rect 15381 6273 15415 6307
rect 15415 6273 15424 6307
rect 15372 6264 15424 6273
rect 17488 6264 17540 6316
rect 19052 6264 19104 6316
rect 11876 6196 11928 6248
rect 11600 6103 11652 6112
rect 11600 6069 11609 6103
rect 11609 6069 11643 6103
rect 11643 6069 11652 6103
rect 11600 6060 11652 6069
rect 15096 6060 15148 6112
rect 17764 6128 17816 6180
rect 19696 6171 19748 6180
rect 19696 6137 19699 6171
rect 19699 6137 19733 6171
rect 19733 6137 19748 6171
rect 19696 6128 19748 6137
rect 16292 6103 16344 6112
rect 16292 6069 16301 6103
rect 16301 6069 16335 6103
rect 16335 6069 16344 6103
rect 16292 6060 16344 6069
rect 20248 6103 20300 6112
rect 20248 6069 20257 6103
rect 20257 6069 20291 6103
rect 20291 6069 20300 6103
rect 20248 6060 20300 6069
rect 24204 6332 24256 6384
rect 20984 6264 21036 6316
rect 21444 6307 21496 6316
rect 21444 6273 21453 6307
rect 21453 6273 21487 6307
rect 21487 6273 21496 6307
rect 21444 6264 21496 6273
rect 23008 6264 23060 6316
rect 24756 6196 24808 6248
rect 25124 6103 25176 6112
rect 25124 6069 25133 6103
rect 25133 6069 25167 6103
rect 25167 6069 25176 6103
rect 25124 6060 25176 6069
rect 9843 5958 9895 6010
rect 9907 5958 9959 6010
rect 9971 5958 10023 6010
rect 10035 5958 10087 6010
rect 19176 5958 19228 6010
rect 19240 5958 19292 6010
rect 19304 5958 19356 6010
rect 19368 5958 19420 6010
rect 17488 5856 17540 5908
rect 19052 5856 19104 5908
rect 20248 5856 20300 5908
rect 15096 5788 15148 5840
rect 16292 5788 16344 5840
rect 16936 5788 16988 5840
rect 21076 5856 21128 5908
rect 24296 5856 24348 5908
rect 13900 5720 13952 5772
rect 15004 5720 15056 5772
rect 21444 5788 21496 5840
rect 18592 5720 18644 5772
rect 23100 5763 23152 5772
rect 23100 5729 23144 5763
rect 23144 5729 23152 5763
rect 23100 5720 23152 5729
rect 25032 5720 25084 5772
rect 16660 5695 16712 5704
rect 16660 5661 16669 5695
rect 16669 5661 16703 5695
rect 16703 5661 16712 5695
rect 16660 5652 16712 5661
rect 17396 5652 17448 5704
rect 18132 5695 18184 5704
rect 18132 5661 18141 5695
rect 18141 5661 18175 5695
rect 18175 5661 18184 5695
rect 18132 5652 18184 5661
rect 19880 5652 19932 5704
rect 10588 5584 10640 5636
rect 11876 5584 11928 5636
rect 23652 5584 23704 5636
rect 15740 5559 15792 5568
rect 15740 5525 15749 5559
rect 15749 5525 15783 5559
rect 15783 5525 15792 5559
rect 15740 5516 15792 5525
rect 5176 5414 5228 5466
rect 5240 5414 5292 5466
rect 5304 5414 5356 5466
rect 5368 5414 5420 5466
rect 14510 5414 14562 5466
rect 14574 5414 14626 5466
rect 14638 5414 14690 5466
rect 14702 5414 14754 5466
rect 23843 5414 23895 5466
rect 23907 5414 23959 5466
rect 23971 5414 24023 5466
rect 24035 5414 24087 5466
rect 13992 5355 14044 5364
rect 13992 5321 14001 5355
rect 14001 5321 14035 5355
rect 14035 5321 14044 5355
rect 13992 5312 14044 5321
rect 15096 5312 15148 5364
rect 16660 5312 16712 5364
rect 16936 5355 16988 5364
rect 16936 5321 16945 5355
rect 16945 5321 16979 5355
rect 16979 5321 16988 5355
rect 16936 5312 16988 5321
rect 18592 5355 18644 5364
rect 18592 5321 18601 5355
rect 18601 5321 18635 5355
rect 18635 5321 18644 5355
rect 18592 5312 18644 5321
rect 20248 5312 20300 5364
rect 23100 5312 23152 5364
rect 23744 5312 23796 5364
rect 24664 5355 24716 5364
rect 24664 5321 24673 5355
rect 24673 5321 24707 5355
rect 24707 5321 24716 5355
rect 24664 5312 24716 5321
rect 25032 5355 25084 5364
rect 25032 5321 25041 5355
rect 25041 5321 25075 5355
rect 25075 5321 25084 5355
rect 25032 5312 25084 5321
rect 17488 5176 17540 5228
rect 19880 5219 19932 5228
rect 19880 5185 19889 5219
rect 19889 5185 19923 5219
rect 19923 5185 19932 5219
rect 19880 5176 19932 5185
rect 24664 5108 24716 5160
rect 14912 4972 14964 5024
rect 15740 5040 15792 5092
rect 17672 5083 17724 5092
rect 17672 5049 17681 5083
rect 17681 5049 17715 5083
rect 17715 5049 17724 5083
rect 17672 5040 17724 5049
rect 18132 5040 18184 5092
rect 19604 5083 19656 5092
rect 19604 5049 19613 5083
rect 19613 5049 19647 5083
rect 19647 5049 19656 5083
rect 19604 5040 19656 5049
rect 19512 4972 19564 5024
rect 9843 4870 9895 4922
rect 9907 4870 9959 4922
rect 9971 4870 10023 4922
rect 10035 4870 10087 4922
rect 19176 4870 19228 4922
rect 19240 4870 19292 4922
rect 19304 4870 19356 4922
rect 19368 4870 19420 4922
rect 15004 4811 15056 4820
rect 15004 4777 15013 4811
rect 15013 4777 15047 4811
rect 15047 4777 15056 4811
rect 15004 4768 15056 4777
rect 17672 4811 17724 4820
rect 17672 4777 17681 4811
rect 17681 4777 17715 4811
rect 17715 4777 17724 4811
rect 17672 4768 17724 4777
rect 23192 4768 23244 4820
rect 15924 4743 15976 4752
rect 15924 4709 15933 4743
rect 15933 4709 15967 4743
rect 15967 4709 15976 4743
rect 15924 4700 15976 4709
rect 16660 4700 16712 4752
rect 19512 4743 19564 4752
rect 19512 4709 19521 4743
rect 19521 4709 19555 4743
rect 19555 4709 19564 4743
rect 19512 4700 19564 4709
rect 18868 4675 18920 4684
rect 18868 4641 18877 4675
rect 18877 4641 18911 4675
rect 18911 4641 18920 4675
rect 18868 4632 18920 4641
rect 24204 4675 24256 4684
rect 24204 4641 24222 4675
rect 24222 4641 24256 4675
rect 24204 4632 24256 4641
rect 16200 4564 16252 4616
rect 5176 4326 5228 4378
rect 5240 4326 5292 4378
rect 5304 4326 5356 4378
rect 5368 4326 5420 4378
rect 14510 4326 14562 4378
rect 14574 4326 14626 4378
rect 14638 4326 14690 4378
rect 14702 4326 14754 4378
rect 23843 4326 23895 4378
rect 23907 4326 23959 4378
rect 23971 4326 24023 4378
rect 24035 4326 24087 4378
rect 14912 4267 14964 4276
rect 14912 4233 14921 4267
rect 14921 4233 14955 4267
rect 14955 4233 14964 4267
rect 14912 4224 14964 4233
rect 18868 4267 18920 4276
rect 18868 4233 18877 4267
rect 18877 4233 18911 4267
rect 18911 4233 18920 4267
rect 18868 4224 18920 4233
rect 15924 4088 15976 4140
rect 16200 4088 16252 4140
rect 25032 4131 25084 4140
rect 25032 4097 25041 4131
rect 25041 4097 25075 4131
rect 25075 4097 25084 4131
rect 25032 4088 25084 4097
rect 14912 4020 14964 4072
rect 23008 3952 23060 4004
rect 24664 3927 24716 3936
rect 24664 3893 24673 3927
rect 24673 3893 24707 3927
rect 24707 3893 24716 3927
rect 24664 3884 24716 3893
rect 9843 3782 9895 3834
rect 9907 3782 9959 3834
rect 9971 3782 10023 3834
rect 10035 3782 10087 3834
rect 19176 3782 19228 3834
rect 19240 3782 19292 3834
rect 19304 3782 19356 3834
rect 19368 3782 19420 3834
rect 16200 3680 16252 3732
rect 16292 3587 16344 3596
rect 16292 3553 16310 3587
rect 16310 3553 16344 3587
rect 16292 3544 16344 3553
rect 5176 3238 5228 3290
rect 5240 3238 5292 3290
rect 5304 3238 5356 3290
rect 5368 3238 5420 3290
rect 14510 3238 14562 3290
rect 14574 3238 14626 3290
rect 14638 3238 14690 3290
rect 14702 3238 14754 3290
rect 23843 3238 23895 3290
rect 23907 3238 23959 3290
rect 23971 3238 24023 3290
rect 24035 3238 24087 3290
rect 16292 2975 16344 2984
rect 16292 2941 16301 2975
rect 16301 2941 16335 2975
rect 16335 2941 16344 2975
rect 16292 2932 16344 2941
rect 9843 2694 9895 2746
rect 9907 2694 9959 2746
rect 9971 2694 10023 2746
rect 10035 2694 10087 2746
rect 19176 2694 19228 2746
rect 19240 2694 19292 2746
rect 19304 2694 19356 2746
rect 19368 2694 19420 2746
rect 23468 2592 23520 2644
rect 24664 2456 24716 2508
rect 24664 2295 24716 2304
rect 24664 2261 24673 2295
rect 24673 2261 24707 2295
rect 24707 2261 24716 2295
rect 24664 2252 24716 2261
rect 5176 2150 5228 2202
rect 5240 2150 5292 2202
rect 5304 2150 5356 2202
rect 5368 2150 5420 2202
rect 14510 2150 14562 2202
rect 14574 2150 14626 2202
rect 14638 2150 14690 2202
rect 14702 2150 14754 2202
rect 23843 2150 23895 2202
rect 23907 2150 23959 2202
rect 23971 2150 24023 2202
rect 24035 2150 24087 2202
<< metal2 >>
rect 6 27520 62 28000
rect 1018 27520 1074 28000
rect 2030 27520 2086 28000
rect 3042 27520 3098 28000
rect 4146 27520 4202 28000
rect 5158 27520 5214 28000
rect 6170 27520 6226 28000
rect 7182 27520 7238 28000
rect 8286 27520 8342 28000
rect 9298 27520 9354 28000
rect 10310 27520 10366 28000
rect 11322 27520 11378 28000
rect 12426 27520 12482 28000
rect 13438 27520 13494 28000
rect 14450 27520 14506 28000
rect 15462 27520 15518 28000
rect 16566 27520 16622 28000
rect 17578 27520 17634 28000
rect 18590 27520 18646 28000
rect 19602 27520 19658 28000
rect 20706 27520 20762 28000
rect 21718 27520 21774 28000
rect 22730 27520 22786 28000
rect 23742 27520 23798 28000
rect 24846 27520 24902 28000
rect 25858 27520 25914 28000
rect 26870 27520 26926 28000
rect 20 24313 48 27520
rect 6 24304 62 24313
rect 6 24239 62 24248
rect 1032 22098 1060 27520
rect 1938 24168 1994 24177
rect 1938 24103 1994 24112
rect 1952 23866 1980 24103
rect 2044 23866 2072 27520
rect 3056 23866 3084 27520
rect 1940 23860 1992 23866
rect 1940 23802 1992 23808
rect 2032 23860 2084 23866
rect 2032 23802 2084 23808
rect 3044 23860 3096 23866
rect 3044 23802 3096 23808
rect 2044 23662 2072 23802
rect 3056 23662 3084 23802
rect 2032 23656 2084 23662
rect 2032 23598 2084 23604
rect 3044 23656 3096 23662
rect 3044 23598 3096 23604
rect 3594 23624 3650 23633
rect 3594 23559 3650 23568
rect 3608 23526 3636 23559
rect 3596 23520 3648 23526
rect 3596 23462 3648 23468
rect 1020 22092 1072 22098
rect 1020 22034 1072 22040
rect 1032 21690 1060 22034
rect 2216 21888 2268 21894
rect 2216 21830 2268 21836
rect 1020 21684 1072 21690
rect 1020 21626 1072 21632
rect 2228 21593 2256 21830
rect 4160 21690 4188 27520
rect 5172 25242 5200 27520
rect 5080 25214 5200 25242
rect 5080 23866 5108 25214
rect 5150 25052 5446 25072
rect 5206 25050 5230 25052
rect 5286 25050 5310 25052
rect 5366 25050 5390 25052
rect 5228 24998 5230 25050
rect 5292 24998 5304 25050
rect 5366 24998 5368 25050
rect 5206 24996 5230 24998
rect 5286 24996 5310 24998
rect 5366 24996 5390 24998
rect 5150 24976 5446 24996
rect 6184 24274 6212 27520
rect 6172 24268 6224 24274
rect 6172 24210 6224 24216
rect 5150 23964 5446 23984
rect 5206 23962 5230 23964
rect 5286 23962 5310 23964
rect 5366 23962 5390 23964
rect 5228 23910 5230 23962
rect 5292 23910 5304 23962
rect 5366 23910 5368 23962
rect 5206 23908 5230 23910
rect 5286 23908 5310 23910
rect 5366 23908 5390 23910
rect 5150 23888 5446 23908
rect 6184 23866 6212 24210
rect 6264 24064 6316 24070
rect 6264 24006 6316 24012
rect 5068 23860 5120 23866
rect 5068 23802 5120 23808
rect 6172 23860 6224 23866
rect 6172 23802 6224 23808
rect 5080 23662 5108 23802
rect 5068 23656 5120 23662
rect 5068 23598 5120 23604
rect 4976 23520 5028 23526
rect 4976 23462 5028 23468
rect 4988 23089 5016 23462
rect 4974 23080 5030 23089
rect 4974 23015 5030 23024
rect 5150 22876 5446 22896
rect 5206 22874 5230 22876
rect 5286 22874 5310 22876
rect 5366 22874 5390 22876
rect 5228 22822 5230 22874
rect 5292 22822 5304 22874
rect 5366 22822 5368 22874
rect 5206 22820 5230 22822
rect 5286 22820 5310 22822
rect 5366 22820 5390 22822
rect 5150 22800 5446 22820
rect 6276 22001 6304 24006
rect 7196 23866 7224 27520
rect 8300 24274 8328 27520
rect 8378 24304 8434 24313
rect 8288 24268 8340 24274
rect 9312 24274 9340 27520
rect 9817 25596 10113 25616
rect 9873 25594 9897 25596
rect 9953 25594 9977 25596
rect 10033 25594 10057 25596
rect 9895 25542 9897 25594
rect 9959 25542 9971 25594
rect 10033 25542 10035 25594
rect 9873 25540 9897 25542
rect 9953 25540 9977 25542
rect 10033 25540 10057 25542
rect 9817 25520 10113 25540
rect 9817 24508 10113 24528
rect 9873 24506 9897 24508
rect 9953 24506 9977 24508
rect 10033 24506 10057 24508
rect 9895 24454 9897 24506
rect 9959 24454 9971 24506
rect 10033 24454 10035 24506
rect 9873 24452 9897 24454
rect 9953 24452 9977 24454
rect 10033 24452 10057 24454
rect 9817 24432 10113 24452
rect 8378 24239 8434 24248
rect 9300 24268 9352 24274
rect 8288 24210 8340 24216
rect 8196 24064 8248 24070
rect 8196 24006 8248 24012
rect 7184 23860 7236 23866
rect 7184 23802 7236 23808
rect 7196 23662 7224 23802
rect 7184 23656 7236 23662
rect 7184 23598 7236 23604
rect 7736 23520 7788 23526
rect 7736 23462 7788 23468
rect 7748 23225 7776 23462
rect 7734 23216 7790 23225
rect 7734 23151 7790 23160
rect 6262 21992 6318 22001
rect 6262 21927 6318 21936
rect 5150 21788 5446 21808
rect 5206 21786 5230 21788
rect 5286 21786 5310 21788
rect 5366 21786 5390 21788
rect 5228 21734 5230 21786
rect 5292 21734 5304 21786
rect 5366 21734 5368 21786
rect 5206 21732 5230 21734
rect 5286 21732 5310 21734
rect 5366 21732 5390 21734
rect 5150 21712 5446 21732
rect 4148 21684 4200 21690
rect 4148 21626 4200 21632
rect 2214 21584 2270 21593
rect 2214 21519 2270 21528
rect 4160 21486 4188 21626
rect 7458 21584 7514 21593
rect 7458 21519 7460 21528
rect 7512 21519 7514 21528
rect 7460 21490 7512 21496
rect 4148 21480 4200 21486
rect 4148 21422 4200 21428
rect 4976 21344 5028 21350
rect 4976 21286 5028 21292
rect 4988 19961 5016 21286
rect 7472 21146 7500 21490
rect 7644 21412 7696 21418
rect 7644 21354 7696 21360
rect 7460 21140 7512 21146
rect 7460 21082 7512 21088
rect 7656 21010 7684 21354
rect 7644 21004 7696 21010
rect 7644 20946 7696 20952
rect 5150 20700 5446 20720
rect 5206 20698 5230 20700
rect 5286 20698 5310 20700
rect 5366 20698 5390 20700
rect 5228 20646 5230 20698
rect 5292 20646 5304 20698
rect 5366 20646 5368 20698
rect 5206 20644 5230 20646
rect 5286 20644 5310 20646
rect 5366 20644 5390 20646
rect 5150 20624 5446 20644
rect 7656 20602 7684 20946
rect 7644 20596 7696 20602
rect 7644 20538 7696 20544
rect 4974 19952 5030 19961
rect 4974 19887 5030 19896
rect 5150 19612 5446 19632
rect 5206 19610 5230 19612
rect 5286 19610 5310 19612
rect 5366 19610 5390 19612
rect 5228 19558 5230 19610
rect 5292 19558 5304 19610
rect 5366 19558 5368 19610
rect 5206 19556 5230 19558
rect 5286 19556 5310 19558
rect 5366 19556 5390 19558
rect 5150 19536 5446 19556
rect 5150 18524 5446 18544
rect 5206 18522 5230 18524
rect 5286 18522 5310 18524
rect 5366 18522 5390 18524
rect 5228 18470 5230 18522
rect 5292 18470 5304 18522
rect 5366 18470 5368 18522
rect 5206 18468 5230 18470
rect 5286 18468 5310 18470
rect 5366 18468 5390 18470
rect 5150 18448 5446 18468
rect 5150 17436 5446 17456
rect 5206 17434 5230 17436
rect 5286 17434 5310 17436
rect 5366 17434 5390 17436
rect 5228 17382 5230 17434
rect 5292 17382 5304 17434
rect 5366 17382 5368 17434
rect 5206 17380 5230 17382
rect 5286 17380 5310 17382
rect 5366 17380 5390 17382
rect 5150 17360 5446 17380
rect 5150 16348 5446 16368
rect 5206 16346 5230 16348
rect 5286 16346 5310 16348
rect 5366 16346 5390 16348
rect 5228 16294 5230 16346
rect 5292 16294 5304 16346
rect 5366 16294 5368 16346
rect 5206 16292 5230 16294
rect 5286 16292 5310 16294
rect 5366 16292 5390 16294
rect 5150 16272 5446 16292
rect 5150 15260 5446 15280
rect 5206 15258 5230 15260
rect 5286 15258 5310 15260
rect 5366 15258 5390 15260
rect 5228 15206 5230 15258
rect 5292 15206 5304 15258
rect 5366 15206 5368 15258
rect 5206 15204 5230 15206
rect 5286 15204 5310 15206
rect 5366 15204 5390 15206
rect 5150 15184 5446 15204
rect 5150 14172 5446 14192
rect 5206 14170 5230 14172
rect 5286 14170 5310 14172
rect 5366 14170 5390 14172
rect 5228 14118 5230 14170
rect 5292 14118 5304 14170
rect 5366 14118 5368 14170
rect 5206 14116 5230 14118
rect 5286 14116 5310 14118
rect 5366 14116 5390 14118
rect 5150 14096 5446 14116
rect 5150 13084 5446 13104
rect 5206 13082 5230 13084
rect 5286 13082 5310 13084
rect 5366 13082 5390 13084
rect 5228 13030 5230 13082
rect 5292 13030 5304 13082
rect 5366 13030 5368 13082
rect 5206 13028 5230 13030
rect 5286 13028 5310 13030
rect 5366 13028 5390 13030
rect 5150 13008 5446 13028
rect 5150 11996 5446 12016
rect 5206 11994 5230 11996
rect 5286 11994 5310 11996
rect 5366 11994 5390 11996
rect 5228 11942 5230 11994
rect 5292 11942 5304 11994
rect 5366 11942 5368 11994
rect 5206 11940 5230 11942
rect 5286 11940 5310 11942
rect 5366 11940 5390 11942
rect 5150 11920 5446 11940
rect 5150 10908 5446 10928
rect 5206 10906 5230 10908
rect 5286 10906 5310 10908
rect 5366 10906 5390 10908
rect 5228 10854 5230 10906
rect 5292 10854 5304 10906
rect 5366 10854 5368 10906
rect 5206 10852 5230 10854
rect 5286 10852 5310 10854
rect 5366 10852 5390 10854
rect 5150 10832 5446 10852
rect 5150 9820 5446 9840
rect 5206 9818 5230 9820
rect 5286 9818 5310 9820
rect 5366 9818 5390 9820
rect 5228 9766 5230 9818
rect 5292 9766 5304 9818
rect 5366 9766 5368 9818
rect 5206 9764 5230 9766
rect 5286 9764 5310 9766
rect 5366 9764 5390 9766
rect 5150 9744 5446 9764
rect 5150 8732 5446 8752
rect 5206 8730 5230 8732
rect 5286 8730 5310 8732
rect 5366 8730 5390 8732
rect 5228 8678 5230 8730
rect 5292 8678 5304 8730
rect 5366 8678 5368 8730
rect 5206 8676 5230 8678
rect 5286 8676 5310 8678
rect 5366 8676 5390 8678
rect 5150 8656 5446 8676
rect 8208 7993 8236 24006
rect 8300 23798 8328 24210
rect 8392 23866 8420 24239
rect 9300 24210 9352 24216
rect 9312 23866 9340 24210
rect 9392 24064 9444 24070
rect 9392 24006 9444 24012
rect 8380 23860 8432 23866
rect 8380 23802 8432 23808
rect 9300 23860 9352 23866
rect 9300 23802 9352 23808
rect 8288 23792 8340 23798
rect 8288 23734 8340 23740
rect 8392 23662 8420 23802
rect 8380 23656 8432 23662
rect 8380 23598 8432 23604
rect 8932 23520 8984 23526
rect 8932 23462 8984 23468
rect 8748 21344 8800 21350
rect 8748 21286 8800 21292
rect 8760 21078 8788 21286
rect 8748 21072 8800 21078
rect 8748 21014 8800 21020
rect 8944 18986 8972 23462
rect 9208 23112 9260 23118
rect 9208 23054 9260 23060
rect 9220 22778 9248 23054
rect 9208 22772 9260 22778
rect 9208 22714 9260 22720
rect 9220 22438 9248 22714
rect 9208 22432 9260 22438
rect 9208 22374 9260 22380
rect 9024 21412 9076 21418
rect 9024 21354 9076 21360
rect 9036 20806 9064 21354
rect 9116 21004 9168 21010
rect 9116 20946 9168 20952
rect 9128 20890 9156 20946
rect 9300 20936 9352 20942
rect 9128 20862 9248 20890
rect 9300 20878 9352 20884
rect 9024 20800 9076 20806
rect 9024 20742 9076 20748
rect 9036 19825 9064 20742
rect 9220 20602 9248 20862
rect 9208 20596 9260 20602
rect 9208 20538 9260 20544
rect 9312 20466 9340 20878
rect 9300 20460 9352 20466
rect 9300 20402 9352 20408
rect 9116 20392 9168 20398
rect 9168 20352 9248 20380
rect 9116 20334 9168 20340
rect 9022 19816 9078 19825
rect 9022 19751 9078 19760
rect 9220 19174 9248 20352
rect 9312 20058 9340 20402
rect 9300 20052 9352 20058
rect 9300 19994 9352 20000
rect 9208 19168 9260 19174
rect 9208 19110 9260 19116
rect 8944 18958 9248 18986
rect 9220 18902 9248 18958
rect 9208 18896 9260 18902
rect 9208 18838 9260 18844
rect 9206 18728 9262 18737
rect 9206 18663 9262 18672
rect 9220 17218 9248 18663
rect 9036 17190 9248 17218
rect 9036 17134 9064 17190
rect 9024 17128 9076 17134
rect 9024 17070 9076 17076
rect 9036 16794 9064 17070
rect 9024 16788 9076 16794
rect 9024 16730 9076 16736
rect 9220 16250 9248 17190
rect 9208 16244 9260 16250
rect 9208 16186 9260 16192
rect 9404 11665 9432 24006
rect 10324 23866 10352 27520
rect 11336 24818 11364 27520
rect 11324 24812 11376 24818
rect 11324 24754 11376 24760
rect 11048 24608 11100 24614
rect 11048 24550 11100 24556
rect 10954 24304 11010 24313
rect 10954 24239 11010 24248
rect 10862 24168 10918 24177
rect 10862 24103 10918 24112
rect 10312 23860 10364 23866
rect 10312 23802 10364 23808
rect 10324 23662 10352 23802
rect 10312 23656 10364 23662
rect 10312 23598 10364 23604
rect 10312 23520 10364 23526
rect 10312 23462 10364 23468
rect 9817 23420 10113 23440
rect 9873 23418 9897 23420
rect 9953 23418 9977 23420
rect 10033 23418 10057 23420
rect 9895 23366 9897 23418
rect 9959 23366 9971 23418
rect 10033 23366 10035 23418
rect 9873 23364 9897 23366
rect 9953 23364 9977 23366
rect 10033 23364 10057 23366
rect 9817 23344 10113 23364
rect 9852 23180 9904 23186
rect 9852 23122 9904 23128
rect 9864 22778 9892 23122
rect 9576 22772 9628 22778
rect 9576 22714 9628 22720
rect 9852 22772 9904 22778
rect 9852 22714 9904 22720
rect 9588 22166 9616 22714
rect 10220 22500 10272 22506
rect 10220 22442 10272 22448
rect 9817 22332 10113 22352
rect 9873 22330 9897 22332
rect 9953 22330 9977 22332
rect 10033 22330 10057 22332
rect 9895 22278 9897 22330
rect 9959 22278 9971 22330
rect 10033 22278 10035 22330
rect 9873 22276 9897 22278
rect 9953 22276 9977 22278
rect 10033 22276 10057 22278
rect 9817 22256 10113 22276
rect 10232 22166 10260 22442
rect 9576 22160 9628 22166
rect 9576 22102 9628 22108
rect 10220 22160 10272 22166
rect 10220 22102 10272 22108
rect 9484 22024 9536 22030
rect 9484 21966 9536 21972
rect 9496 21554 9524 21966
rect 9588 21690 9616 22102
rect 9576 21684 9628 21690
rect 9576 21626 9628 21632
rect 10220 21684 10272 21690
rect 10220 21626 10272 21632
rect 9484 21548 9536 21554
rect 9484 21490 9536 21496
rect 9817 21244 10113 21264
rect 9873 21242 9897 21244
rect 9953 21242 9977 21244
rect 10033 21242 10057 21244
rect 9895 21190 9897 21242
rect 9959 21190 9971 21242
rect 10033 21190 10035 21242
rect 9873 21188 9897 21190
rect 9953 21188 9977 21190
rect 10033 21188 10057 21190
rect 9817 21168 10113 21188
rect 10232 21146 10260 21626
rect 10220 21140 10272 21146
rect 10220 21082 10272 21088
rect 9668 21072 9720 21078
rect 9668 21014 9720 21020
rect 9680 20330 9708 21014
rect 9668 20324 9720 20330
rect 9668 20266 9720 20272
rect 9576 19916 9628 19922
rect 9576 19858 9628 19864
rect 9588 19310 9616 19858
rect 9484 19304 9536 19310
rect 9484 19246 9536 19252
rect 9576 19304 9628 19310
rect 9576 19246 9628 19252
rect 9496 18737 9524 19246
rect 9482 18728 9538 18737
rect 9482 18663 9538 18672
rect 9588 18630 9616 19246
rect 9576 18624 9628 18630
rect 9574 18592 9576 18601
rect 9628 18592 9630 18601
rect 9574 18527 9630 18536
rect 9680 17814 9708 20266
rect 9817 20156 10113 20176
rect 9873 20154 9897 20156
rect 9953 20154 9977 20156
rect 10033 20154 10057 20156
rect 9895 20102 9897 20154
rect 9959 20102 9971 20154
rect 10033 20102 10035 20154
rect 9873 20100 9897 20102
rect 9953 20100 9977 20102
rect 10033 20100 10057 20102
rect 9817 20080 10113 20100
rect 10324 19938 10352 23462
rect 10876 23254 10904 24103
rect 10968 23866 10996 24239
rect 10956 23860 11008 23866
rect 10956 23802 11008 23808
rect 10956 23656 11008 23662
rect 10956 23598 11008 23604
rect 10864 23248 10916 23254
rect 10864 23190 10916 23196
rect 10876 22234 10904 23190
rect 10968 22778 10996 23598
rect 10956 22772 11008 22778
rect 10956 22714 11008 22720
rect 10864 22228 10916 22234
rect 10864 22170 10916 22176
rect 10324 19910 10444 19938
rect 10312 19848 10364 19854
rect 10312 19790 10364 19796
rect 10324 19174 10352 19790
rect 10312 19168 10364 19174
rect 10312 19110 10364 19116
rect 9817 19068 10113 19088
rect 9873 19066 9897 19068
rect 9953 19066 9977 19068
rect 10033 19066 10057 19068
rect 9895 19014 9897 19066
rect 9959 19014 9971 19066
rect 10033 19014 10035 19066
rect 9873 19012 9897 19014
rect 9953 19012 9977 19014
rect 10033 19012 10057 19014
rect 9817 18992 10113 19012
rect 9852 18896 9904 18902
rect 9852 18838 9904 18844
rect 10220 18896 10272 18902
rect 10220 18838 10272 18844
rect 9864 18426 9892 18838
rect 9852 18420 9904 18426
rect 9852 18362 9904 18368
rect 10232 18222 10260 18838
rect 10220 18216 10272 18222
rect 10220 18158 10272 18164
rect 9817 17980 10113 18000
rect 9873 17978 9897 17980
rect 9953 17978 9977 17980
rect 10033 17978 10057 17980
rect 9895 17926 9897 17978
rect 9959 17926 9971 17978
rect 10033 17926 10035 17978
rect 9873 17924 9897 17926
rect 9953 17924 9977 17926
rect 10033 17924 10057 17926
rect 9817 17904 10113 17924
rect 10232 17882 10260 18158
rect 10220 17876 10272 17882
rect 10220 17818 10272 17824
rect 9668 17808 9720 17814
rect 10324 17762 10352 19110
rect 9668 17750 9720 17756
rect 9484 17672 9536 17678
rect 9484 17614 9536 17620
rect 9496 17202 9524 17614
rect 9680 17338 9708 17750
rect 10232 17734 10352 17762
rect 9668 17332 9720 17338
rect 9668 17274 9720 17280
rect 9484 17196 9536 17202
rect 9484 17138 9536 17144
rect 9496 16794 9524 17138
rect 9817 16892 10113 16912
rect 9873 16890 9897 16892
rect 9953 16890 9977 16892
rect 10033 16890 10057 16892
rect 9895 16838 9897 16890
rect 9959 16838 9971 16890
rect 10033 16838 10035 16890
rect 9873 16836 9897 16838
rect 9953 16836 9977 16838
rect 10033 16836 10057 16838
rect 9817 16816 10113 16836
rect 9484 16788 9536 16794
rect 9484 16730 9536 16736
rect 10232 16658 10260 17734
rect 10416 17626 10444 19910
rect 10680 18760 10732 18766
rect 10680 18702 10732 18708
rect 10588 18624 10640 18630
rect 10588 18566 10640 18572
rect 10600 18358 10628 18566
rect 10588 18352 10640 18358
rect 10588 18294 10640 18300
rect 10324 17598 10444 17626
rect 10220 16652 10272 16658
rect 10220 16594 10272 16600
rect 10232 16250 10260 16594
rect 10220 16244 10272 16250
rect 10220 16186 10272 16192
rect 10220 15904 10272 15910
rect 10218 15872 10220 15881
rect 10272 15872 10274 15881
rect 9817 15804 10113 15824
rect 10218 15807 10274 15816
rect 9873 15802 9897 15804
rect 9953 15802 9977 15804
rect 10033 15802 10057 15804
rect 9895 15750 9897 15802
rect 9959 15750 9971 15802
rect 10033 15750 10035 15802
rect 9873 15748 9897 15750
rect 9953 15748 9977 15750
rect 10033 15748 10057 15750
rect 9817 15728 10113 15748
rect 9817 14716 10113 14736
rect 9873 14714 9897 14716
rect 9953 14714 9977 14716
rect 10033 14714 10057 14716
rect 9895 14662 9897 14714
rect 9959 14662 9971 14714
rect 10033 14662 10035 14714
rect 9873 14660 9897 14662
rect 9953 14660 9977 14662
rect 10033 14660 10057 14662
rect 9817 14640 10113 14660
rect 9817 13628 10113 13648
rect 9873 13626 9897 13628
rect 9953 13626 9977 13628
rect 10033 13626 10057 13628
rect 9895 13574 9897 13626
rect 9959 13574 9971 13626
rect 10033 13574 10035 13626
rect 9873 13572 9897 13574
rect 9953 13572 9977 13574
rect 10033 13572 10057 13574
rect 9817 13552 10113 13572
rect 9817 12540 10113 12560
rect 9873 12538 9897 12540
rect 9953 12538 9977 12540
rect 10033 12538 10057 12540
rect 9895 12486 9897 12538
rect 9959 12486 9971 12538
rect 10033 12486 10035 12538
rect 9873 12484 9897 12486
rect 9953 12484 9977 12486
rect 10033 12484 10057 12486
rect 9817 12464 10113 12484
rect 9390 11656 9446 11665
rect 9390 11591 9446 11600
rect 9817 11452 10113 11472
rect 9873 11450 9897 11452
rect 9953 11450 9977 11452
rect 10033 11450 10057 11452
rect 9895 11398 9897 11450
rect 9959 11398 9971 11450
rect 10033 11398 10035 11450
rect 9873 11396 9897 11398
rect 9953 11396 9977 11398
rect 10033 11396 10057 11398
rect 9817 11376 10113 11396
rect 9817 10364 10113 10384
rect 9873 10362 9897 10364
rect 9953 10362 9977 10364
rect 10033 10362 10057 10364
rect 9895 10310 9897 10362
rect 9959 10310 9971 10362
rect 10033 10310 10035 10362
rect 9873 10308 9897 10310
rect 9953 10308 9977 10310
rect 10033 10308 10057 10310
rect 9817 10288 10113 10308
rect 9817 9276 10113 9296
rect 9873 9274 9897 9276
rect 9953 9274 9977 9276
rect 10033 9274 10057 9276
rect 9895 9222 9897 9274
rect 9959 9222 9971 9274
rect 10033 9222 10035 9274
rect 9873 9220 9897 9222
rect 9953 9220 9977 9222
rect 10033 9220 10057 9222
rect 9817 9200 10113 9220
rect 9817 8188 10113 8208
rect 9873 8186 9897 8188
rect 9953 8186 9977 8188
rect 10033 8186 10057 8188
rect 9895 8134 9897 8186
rect 9959 8134 9971 8186
rect 10033 8134 10035 8186
rect 9873 8132 9897 8134
rect 9953 8132 9977 8134
rect 10033 8132 10057 8134
rect 9817 8112 10113 8132
rect 8194 7984 8250 7993
rect 8194 7919 8250 7928
rect 5150 7644 5446 7664
rect 5206 7642 5230 7644
rect 5286 7642 5310 7644
rect 5366 7642 5390 7644
rect 5228 7590 5230 7642
rect 5292 7590 5304 7642
rect 5366 7590 5368 7642
rect 5206 7588 5230 7590
rect 5286 7588 5310 7590
rect 5366 7588 5390 7590
rect 5150 7568 5446 7588
rect 9817 7100 10113 7120
rect 9873 7098 9897 7100
rect 9953 7098 9977 7100
rect 10033 7098 10057 7100
rect 9895 7046 9897 7098
rect 9959 7046 9971 7098
rect 10033 7046 10035 7098
rect 9873 7044 9897 7046
rect 9953 7044 9977 7046
rect 10033 7044 10057 7046
rect 9817 7024 10113 7044
rect 5150 6556 5446 6576
rect 5206 6554 5230 6556
rect 5286 6554 5310 6556
rect 5366 6554 5390 6556
rect 5228 6502 5230 6554
rect 5292 6502 5304 6554
rect 5366 6502 5368 6554
rect 5206 6500 5230 6502
rect 5286 6500 5310 6502
rect 5366 6500 5390 6502
rect 5150 6480 5446 6500
rect 9817 6012 10113 6032
rect 9873 6010 9897 6012
rect 9953 6010 9977 6012
rect 10033 6010 10057 6012
rect 9895 5958 9897 6010
rect 9959 5958 9971 6010
rect 10033 5958 10035 6010
rect 9873 5956 9897 5958
rect 9953 5956 9977 5958
rect 10033 5956 10057 5958
rect 9817 5936 10113 5956
rect 8286 5808 8342 5817
rect 8286 5743 8342 5752
rect 5150 5468 5446 5488
rect 5206 5466 5230 5468
rect 5286 5466 5310 5468
rect 5366 5466 5390 5468
rect 5228 5414 5230 5466
rect 5292 5414 5304 5466
rect 5366 5414 5368 5466
rect 5206 5412 5230 5414
rect 5286 5412 5310 5414
rect 5366 5412 5390 5414
rect 5150 5392 5446 5412
rect 5150 4380 5446 4400
rect 5206 4378 5230 4380
rect 5286 4378 5310 4380
rect 5366 4378 5390 4380
rect 5228 4326 5230 4378
rect 5292 4326 5304 4378
rect 5366 4326 5368 4378
rect 5206 4324 5230 4326
rect 5286 4324 5310 4326
rect 5366 4324 5390 4326
rect 5150 4304 5446 4324
rect 4790 4040 4846 4049
rect 4790 3975 4846 3984
rect 1294 3496 1350 3505
rect 1294 3431 1350 3440
rect 1308 480 1336 3431
rect 4804 480 4832 3975
rect 5150 3292 5446 3312
rect 5206 3290 5230 3292
rect 5286 3290 5310 3292
rect 5366 3290 5390 3292
rect 5228 3238 5230 3290
rect 5292 3238 5304 3290
rect 5366 3238 5368 3290
rect 5206 3236 5230 3238
rect 5286 3236 5310 3238
rect 5366 3236 5390 3238
rect 5150 3216 5446 3236
rect 5150 2204 5446 2224
rect 5206 2202 5230 2204
rect 5286 2202 5310 2204
rect 5366 2202 5390 2204
rect 5228 2150 5230 2202
rect 5292 2150 5304 2202
rect 5366 2150 5368 2202
rect 5206 2148 5230 2150
rect 5286 2148 5310 2150
rect 5366 2148 5390 2150
rect 5150 2128 5446 2148
rect 8300 480 8328 5743
rect 10324 5409 10352 17598
rect 10404 17196 10456 17202
rect 10404 17138 10456 17144
rect 10416 16697 10444 17138
rect 10402 16688 10458 16697
rect 10402 16623 10404 16632
rect 10456 16623 10458 16632
rect 10404 16594 10456 16600
rect 10600 16153 10628 18294
rect 10692 18290 10720 18702
rect 10680 18284 10732 18290
rect 10680 18226 10732 18232
rect 10680 17536 10732 17542
rect 10680 17478 10732 17484
rect 10692 17134 10720 17478
rect 10680 17128 10732 17134
rect 10680 17070 10732 17076
rect 10692 16726 10720 17070
rect 10680 16720 10732 16726
rect 10680 16662 10732 16668
rect 10770 16688 10826 16697
rect 10770 16623 10826 16632
rect 10784 16250 10812 16623
rect 10772 16244 10824 16250
rect 10772 16186 10824 16192
rect 10586 16144 10642 16153
rect 10586 16079 10642 16088
rect 10586 15872 10642 15881
rect 10586 15807 10642 15816
rect 10600 11529 10628 15807
rect 10586 11520 10642 11529
rect 10586 11455 10642 11464
rect 10600 11121 10628 11455
rect 10586 11112 10642 11121
rect 10586 11047 10642 11056
rect 10770 11112 10826 11121
rect 10770 11047 10826 11056
rect 10588 5636 10640 5642
rect 10588 5578 10640 5584
rect 10310 5400 10366 5409
rect 10310 5335 10366 5344
rect 9817 4924 10113 4944
rect 9873 4922 9897 4924
rect 9953 4922 9977 4924
rect 10033 4922 10057 4924
rect 9895 4870 9897 4922
rect 9959 4870 9971 4922
rect 10033 4870 10035 4922
rect 9873 4868 9897 4870
rect 9953 4868 9977 4870
rect 10033 4868 10057 4870
rect 9817 4848 10113 4868
rect 9817 3836 10113 3856
rect 9873 3834 9897 3836
rect 9953 3834 9977 3836
rect 10033 3834 10057 3836
rect 9895 3782 9897 3834
rect 9959 3782 9971 3834
rect 10033 3782 10035 3834
rect 9873 3780 9897 3782
rect 9953 3780 9977 3782
rect 10033 3780 10057 3782
rect 9817 3760 10113 3780
rect 10600 3505 10628 5578
rect 10784 4049 10812 11047
rect 11060 6905 11088 24550
rect 11692 24200 11744 24206
rect 11692 24142 11744 24148
rect 12152 24200 12204 24206
rect 12152 24142 12204 24148
rect 11704 23866 11732 24142
rect 12164 23866 12192 24142
rect 11692 23860 11744 23866
rect 11692 23802 11744 23808
rect 12152 23860 12204 23866
rect 12152 23802 12204 23808
rect 12164 23594 12192 23802
rect 12152 23588 12204 23594
rect 12152 23530 12204 23536
rect 11324 23248 11376 23254
rect 11324 23190 11376 23196
rect 12440 23202 12468 27520
rect 13452 27418 13480 27520
rect 13360 27390 13480 27418
rect 13360 26330 13388 27390
rect 13268 26302 13388 26330
rect 13268 25362 13296 26302
rect 13256 25356 13308 25362
rect 13256 25298 13308 25304
rect 13268 24954 13296 25298
rect 14464 25242 14492 27520
rect 14372 25214 14492 25242
rect 13256 24948 13308 24954
rect 13256 24890 13308 24896
rect 12612 24744 12664 24750
rect 12612 24686 12664 24692
rect 14084 24744 14136 24750
rect 14084 24686 14136 24692
rect 11336 22778 11364 23190
rect 12440 23174 12560 23202
rect 12428 23112 12480 23118
rect 12428 23054 12480 23060
rect 11324 22772 11376 22778
rect 11324 22714 11376 22720
rect 11336 22098 11364 22714
rect 12440 22642 12468 23054
rect 12428 22636 12480 22642
rect 12428 22578 12480 22584
rect 12060 22500 12112 22506
rect 12060 22442 12112 22448
rect 11876 22432 11928 22438
rect 11876 22374 11928 22380
rect 11888 22234 11916 22374
rect 11876 22228 11928 22234
rect 11876 22170 11928 22176
rect 11324 22092 11376 22098
rect 11324 22034 11376 22040
rect 11336 21690 11364 22034
rect 12072 21894 12100 22442
rect 12060 21888 12112 21894
rect 12060 21830 12112 21836
rect 12532 21690 12560 23174
rect 11324 21684 11376 21690
rect 11324 21626 11376 21632
rect 12520 21684 12572 21690
rect 12520 21626 12572 21632
rect 11336 21146 11364 21626
rect 12532 21486 12560 21626
rect 12520 21480 12572 21486
rect 12520 21422 12572 21428
rect 11692 21412 11744 21418
rect 11692 21354 11744 21360
rect 11324 21140 11376 21146
rect 11324 21082 11376 21088
rect 11704 21078 11732 21354
rect 12244 21344 12296 21350
rect 12244 21286 12296 21292
rect 11692 21072 11744 21078
rect 11692 21014 11744 21020
rect 11232 20936 11284 20942
rect 11232 20878 11284 20884
rect 11244 20330 11272 20878
rect 11232 20324 11284 20330
rect 11232 20266 11284 20272
rect 11704 20262 11732 21014
rect 12060 20392 12112 20398
rect 12060 20334 12112 20340
rect 11876 20324 11928 20330
rect 11876 20266 11928 20272
rect 11692 20256 11744 20262
rect 11692 20198 11744 20204
rect 11888 20210 11916 20266
rect 11888 20182 12008 20210
rect 11508 19916 11560 19922
rect 11508 19858 11560 19864
rect 11520 19310 11548 19858
rect 11508 19304 11560 19310
rect 11506 19272 11508 19281
rect 11560 19272 11562 19281
rect 11506 19207 11562 19216
rect 11980 19174 12008 20182
rect 12072 19854 12100 20334
rect 12152 19916 12204 19922
rect 12152 19858 12204 19864
rect 12060 19848 12112 19854
rect 12060 19790 12112 19796
rect 12060 19304 12112 19310
rect 12060 19246 12112 19252
rect 11968 19168 12020 19174
rect 11968 19110 12020 19116
rect 12072 18986 12100 19246
rect 12164 19242 12192 19858
rect 12152 19236 12204 19242
rect 12152 19178 12204 19184
rect 11980 18958 12100 18986
rect 11980 18766 12008 18958
rect 11324 18760 11376 18766
rect 11968 18760 12020 18766
rect 11324 18702 11376 18708
rect 11966 18728 11968 18737
rect 12020 18728 12022 18737
rect 11336 17678 11364 18702
rect 11966 18663 12022 18672
rect 12060 18624 12112 18630
rect 12060 18566 12112 18572
rect 12072 18290 12100 18566
rect 12060 18284 12112 18290
rect 12060 18226 12112 18232
rect 11784 18148 11836 18154
rect 11784 18090 11836 18096
rect 11600 17808 11652 17814
rect 11600 17750 11652 17756
rect 11324 17672 11376 17678
rect 11324 17614 11376 17620
rect 11336 16794 11364 17614
rect 11612 17338 11640 17750
rect 11600 17332 11652 17338
rect 11600 17274 11652 17280
rect 11612 16794 11640 17274
rect 11796 17134 11824 18090
rect 11784 17128 11836 17134
rect 11784 17070 11836 17076
rect 11324 16788 11376 16794
rect 11324 16730 11376 16736
rect 11600 16788 11652 16794
rect 11600 16730 11652 16736
rect 11796 16658 11824 17070
rect 11784 16652 11836 16658
rect 11784 16594 11836 16600
rect 11796 16250 11824 16594
rect 11784 16244 11836 16250
rect 11784 16186 11836 16192
rect 12152 13388 12204 13394
rect 12152 13330 12204 13336
rect 12164 12782 12192 13330
rect 12152 12776 12204 12782
rect 12152 12718 12204 12724
rect 12256 9081 12284 21286
rect 12624 18358 12652 24686
rect 12888 24268 12940 24274
rect 12888 24210 12940 24216
rect 13808 24268 13860 24274
rect 13808 24210 13860 24216
rect 12900 23254 12928 24210
rect 13820 23866 13848 24210
rect 14096 23866 14124 24686
rect 14176 24676 14228 24682
rect 14176 24618 14228 24624
rect 14188 24206 14216 24618
rect 14372 24274 14400 25214
rect 14484 25052 14780 25072
rect 14540 25050 14564 25052
rect 14620 25050 14644 25052
rect 14700 25050 14724 25052
rect 14562 24998 14564 25050
rect 14626 24998 14638 25050
rect 14700 24998 14702 25050
rect 14540 24996 14564 24998
rect 14620 24996 14644 24998
rect 14700 24996 14724 24998
rect 14484 24976 14780 24996
rect 15476 24750 15504 27520
rect 15464 24744 15516 24750
rect 14450 24712 14506 24721
rect 15464 24686 15516 24692
rect 14450 24647 14506 24656
rect 14464 24614 14492 24647
rect 14452 24608 14504 24614
rect 14452 24550 14504 24556
rect 16016 24608 16068 24614
rect 16016 24550 16068 24556
rect 15002 24440 15058 24449
rect 15002 24375 15004 24384
rect 15056 24375 15058 24384
rect 15004 24346 15056 24352
rect 14360 24268 14412 24274
rect 14360 24210 14412 24216
rect 14176 24200 14228 24206
rect 14176 24142 14228 24148
rect 14188 23866 14216 24142
rect 14268 24064 14320 24070
rect 14268 24006 14320 24012
rect 13808 23860 13860 23866
rect 13808 23802 13860 23808
rect 14084 23860 14136 23866
rect 14084 23802 14136 23808
rect 14176 23860 14228 23866
rect 14176 23802 14228 23808
rect 14082 23624 14138 23633
rect 13072 23588 13124 23594
rect 14082 23559 14138 23568
rect 13072 23530 13124 23536
rect 13084 23254 13112 23530
rect 12888 23248 12940 23254
rect 12888 23190 12940 23196
rect 13072 23248 13124 23254
rect 13072 23190 13124 23196
rect 12900 22438 12928 23190
rect 14096 22642 14124 23559
rect 14084 22636 14136 22642
rect 14084 22578 14136 22584
rect 12888 22432 12940 22438
rect 12888 22374 12940 22380
rect 13348 22432 13400 22438
rect 13348 22374 13400 22380
rect 12704 21888 12756 21894
rect 12704 21830 12756 21836
rect 12716 20369 12744 21830
rect 12900 20602 12928 22374
rect 13360 22114 13388 22374
rect 14096 22234 14124 22578
rect 14084 22228 14136 22234
rect 14084 22170 14136 22176
rect 13268 22098 13388 22114
rect 13256 22092 13388 22098
rect 13308 22086 13388 22092
rect 13808 22092 13860 22098
rect 13256 22034 13308 22040
rect 13808 22034 13860 22040
rect 13268 22003 13296 22034
rect 13820 21690 13848 22034
rect 13808 21684 13860 21690
rect 13808 21626 13860 21632
rect 13624 21480 13676 21486
rect 13624 21422 13676 21428
rect 13636 20806 13664 21422
rect 13624 20800 13676 20806
rect 13624 20742 13676 20748
rect 13900 20800 13952 20806
rect 13900 20742 13952 20748
rect 12888 20596 12940 20602
rect 12888 20538 12940 20544
rect 12702 20360 12758 20369
rect 12702 20295 12758 20304
rect 13348 19916 13400 19922
rect 13348 19858 13400 19864
rect 13360 19446 13388 19858
rect 13348 19440 13400 19446
rect 13176 19388 13348 19394
rect 13176 19382 13400 19388
rect 13176 19366 13388 19382
rect 13176 19281 13204 19366
rect 13360 19317 13388 19366
rect 13256 19304 13308 19310
rect 13162 19272 13218 19281
rect 13308 19252 13388 19258
rect 13256 19246 13388 19252
rect 13268 19230 13388 19246
rect 13162 19207 13164 19216
rect 13216 19207 13218 19216
rect 13164 19178 13216 19184
rect 12612 18352 12664 18358
rect 12612 18294 12664 18300
rect 12624 17814 12652 18294
rect 12612 17808 12664 17814
rect 12612 17750 12664 17756
rect 13256 17672 13308 17678
rect 13256 17614 13308 17620
rect 12704 17536 12756 17542
rect 12704 17478 12756 17484
rect 12980 17536 13032 17542
rect 12980 17478 13032 17484
rect 12520 17264 12572 17270
rect 12520 17206 12572 17212
rect 12532 15910 12560 17206
rect 12716 17066 12744 17478
rect 12992 17338 13020 17478
rect 12980 17332 13032 17338
rect 12980 17274 13032 17280
rect 12704 17060 12756 17066
rect 12704 17002 12756 17008
rect 12992 16794 13020 17274
rect 13268 17202 13296 17614
rect 13360 17338 13388 19230
rect 13636 19174 13664 20742
rect 13912 20398 13940 20742
rect 13900 20392 13952 20398
rect 13900 20334 13952 20340
rect 13912 19990 13940 20334
rect 13900 19984 13952 19990
rect 13900 19926 13952 19932
rect 13992 19916 14044 19922
rect 13992 19858 14044 19864
rect 14004 19310 14032 19858
rect 13716 19304 13768 19310
rect 13716 19246 13768 19252
rect 13992 19304 14044 19310
rect 13992 19246 14044 19252
rect 13624 19168 13676 19174
rect 13624 19110 13676 19116
rect 13728 18766 13756 19246
rect 14004 18970 14032 19246
rect 13992 18964 14044 18970
rect 13992 18906 14044 18912
rect 13716 18760 13768 18766
rect 13716 18702 13768 18708
rect 13624 18624 13676 18630
rect 13624 18566 13676 18572
rect 13806 18592 13862 18601
rect 13636 18426 13664 18566
rect 13806 18527 13862 18536
rect 13624 18420 13676 18426
rect 13624 18362 13676 18368
rect 13440 18284 13492 18290
rect 13440 18226 13492 18232
rect 13452 18086 13480 18226
rect 13440 18080 13492 18086
rect 13440 18022 13492 18028
rect 13452 17678 13480 18022
rect 13636 17814 13664 18362
rect 13716 18148 13768 18154
rect 13716 18090 13768 18096
rect 13624 17808 13676 17814
rect 13624 17750 13676 17756
rect 13728 17746 13756 18090
rect 13820 17882 13848 18527
rect 14004 18426 14032 18906
rect 13992 18420 14044 18426
rect 13992 18362 14044 18368
rect 13992 18284 14044 18290
rect 13992 18226 14044 18232
rect 14004 17882 14032 18226
rect 13808 17876 13860 17882
rect 13808 17818 13860 17824
rect 13992 17876 14044 17882
rect 13992 17818 14044 17824
rect 13716 17740 13768 17746
rect 13716 17682 13768 17688
rect 13440 17672 13492 17678
rect 13440 17614 13492 17620
rect 13440 17536 13492 17542
rect 13440 17478 13492 17484
rect 13348 17332 13400 17338
rect 13348 17274 13400 17280
rect 13256 17196 13308 17202
rect 13256 17138 13308 17144
rect 13164 17060 13216 17066
rect 13164 17002 13216 17008
rect 12980 16788 13032 16794
rect 12980 16730 13032 16736
rect 12612 16720 12664 16726
rect 12612 16662 12664 16668
rect 12520 15904 12572 15910
rect 12520 15846 12572 15852
rect 12336 13796 12388 13802
rect 12336 13738 12388 13744
rect 12348 13530 12376 13738
rect 12336 13524 12388 13530
rect 12336 13466 12388 13472
rect 12532 11830 12560 15846
rect 12520 11824 12572 11830
rect 12520 11766 12572 11772
rect 12532 11354 12560 11766
rect 12520 11348 12572 11354
rect 12520 11290 12572 11296
rect 12520 11212 12572 11218
rect 12520 11154 12572 11160
rect 12532 10810 12560 11154
rect 12520 10804 12572 10810
rect 12520 10746 12572 10752
rect 12624 9722 12652 16662
rect 12992 16454 13020 16730
rect 13176 16658 13204 17002
rect 13268 16998 13296 17138
rect 13452 17134 13480 17478
rect 14004 17270 14032 17818
rect 14280 17626 14308 24006
rect 14484 23964 14780 23984
rect 14540 23962 14564 23964
rect 14620 23962 14644 23964
rect 14700 23962 14724 23964
rect 14562 23910 14564 23962
rect 14626 23910 14638 23962
rect 14700 23910 14702 23962
rect 14540 23908 14564 23910
rect 14620 23908 14644 23910
rect 14700 23908 14724 23910
rect 14484 23888 14780 23908
rect 15832 23588 15884 23594
rect 15832 23530 15884 23536
rect 15188 23520 15240 23526
rect 15188 23462 15240 23468
rect 15200 23254 15228 23462
rect 15188 23248 15240 23254
rect 15188 23190 15240 23196
rect 15096 23112 15148 23118
rect 15096 23054 15148 23060
rect 14484 22876 14780 22896
rect 14540 22874 14564 22876
rect 14620 22874 14644 22876
rect 14700 22874 14724 22876
rect 14562 22822 14564 22874
rect 14626 22822 14638 22874
rect 14700 22822 14702 22874
rect 14540 22820 14564 22822
rect 14620 22820 14644 22822
rect 14700 22820 14724 22822
rect 14484 22800 14780 22820
rect 15108 22778 15136 23054
rect 15096 22772 15148 22778
rect 15096 22714 15148 22720
rect 14912 22160 14964 22166
rect 14912 22102 14964 22108
rect 14484 21788 14780 21808
rect 14540 21786 14564 21788
rect 14620 21786 14644 21788
rect 14700 21786 14724 21788
rect 14562 21734 14564 21786
rect 14626 21734 14638 21786
rect 14700 21734 14702 21786
rect 14540 21732 14564 21734
rect 14620 21732 14644 21734
rect 14700 21732 14724 21734
rect 14484 21712 14780 21732
rect 14924 21690 14952 22102
rect 14912 21684 14964 21690
rect 14912 21626 14964 21632
rect 15108 21554 15136 22714
rect 15200 22642 15228 23190
rect 15648 22976 15700 22982
rect 15648 22918 15700 22924
rect 15660 22642 15688 22918
rect 15188 22636 15240 22642
rect 15188 22578 15240 22584
rect 15648 22636 15700 22642
rect 15648 22578 15700 22584
rect 15660 22166 15688 22578
rect 15844 22506 15872 23530
rect 15924 23112 15976 23118
rect 15924 23054 15976 23060
rect 15936 22642 15964 23054
rect 15924 22636 15976 22642
rect 15924 22578 15976 22584
rect 15832 22500 15884 22506
rect 15832 22442 15884 22448
rect 15648 22160 15700 22166
rect 15648 22102 15700 22108
rect 15844 21894 15872 22442
rect 15924 22024 15976 22030
rect 15924 21966 15976 21972
rect 15832 21888 15884 21894
rect 15832 21830 15884 21836
rect 15096 21548 15148 21554
rect 15096 21490 15148 21496
rect 15372 21004 15424 21010
rect 15372 20946 15424 20952
rect 15280 20936 15332 20942
rect 15280 20878 15332 20884
rect 14484 20700 14780 20720
rect 14540 20698 14564 20700
rect 14620 20698 14644 20700
rect 14700 20698 14724 20700
rect 14562 20646 14564 20698
rect 14626 20646 14638 20698
rect 14700 20646 14702 20698
rect 14540 20644 14564 20646
rect 14620 20644 14644 20646
rect 14700 20644 14724 20646
rect 14484 20624 14780 20644
rect 15292 20262 15320 20878
rect 15280 20256 15332 20262
rect 15280 20198 15332 20204
rect 14912 19916 14964 19922
rect 14912 19858 14964 19864
rect 14820 19712 14872 19718
rect 14820 19654 14872 19660
rect 14484 19612 14780 19632
rect 14540 19610 14564 19612
rect 14620 19610 14644 19612
rect 14700 19610 14724 19612
rect 14562 19558 14564 19610
rect 14626 19558 14638 19610
rect 14700 19558 14702 19610
rect 14540 19556 14564 19558
rect 14620 19556 14644 19558
rect 14700 19556 14724 19558
rect 14484 19536 14780 19556
rect 14636 18760 14688 18766
rect 14832 18714 14860 19654
rect 14924 19446 14952 19858
rect 14912 19440 14964 19446
rect 14912 19382 14964 19388
rect 14924 18902 14952 19382
rect 15292 19310 15320 20198
rect 15384 19922 15412 20946
rect 15740 20936 15792 20942
rect 15740 20878 15792 20884
rect 15752 20466 15780 20878
rect 15844 20602 15872 21830
rect 15936 21622 15964 21966
rect 15924 21616 15976 21622
rect 15922 21584 15924 21593
rect 15976 21584 15978 21593
rect 15922 21519 15978 21528
rect 15832 20596 15884 20602
rect 15832 20538 15884 20544
rect 15740 20460 15792 20466
rect 15740 20402 15792 20408
rect 15372 19916 15424 19922
rect 15372 19858 15424 19864
rect 15280 19304 15332 19310
rect 15280 19246 15332 19252
rect 15556 19304 15608 19310
rect 15556 19246 15608 19252
rect 14912 18896 14964 18902
rect 14912 18838 14964 18844
rect 15292 18834 15320 19246
rect 15280 18828 15332 18834
rect 15280 18770 15332 18776
rect 14688 18708 14860 18714
rect 14636 18702 14860 18708
rect 14648 18686 14860 18702
rect 14484 18524 14780 18544
rect 14540 18522 14564 18524
rect 14620 18522 14644 18524
rect 14700 18522 14724 18524
rect 14562 18470 14564 18522
rect 14626 18470 14638 18522
rect 14700 18470 14702 18522
rect 14540 18468 14564 18470
rect 14620 18468 14644 18470
rect 14700 18468 14724 18470
rect 14484 18448 14780 18468
rect 14544 18080 14596 18086
rect 14544 18022 14596 18028
rect 14556 17882 14584 18022
rect 14544 17876 14596 17882
rect 14544 17818 14596 17824
rect 14096 17598 14308 17626
rect 13992 17264 14044 17270
rect 13992 17206 14044 17212
rect 13440 17128 13492 17134
rect 13440 17070 13492 17076
rect 13256 16992 13308 16998
rect 13256 16934 13308 16940
rect 13164 16652 13216 16658
rect 13164 16594 13216 16600
rect 13176 16561 13204 16594
rect 13268 16590 13296 16934
rect 13808 16788 13860 16794
rect 13808 16730 13860 16736
rect 13820 16697 13848 16730
rect 13806 16688 13862 16697
rect 13806 16623 13862 16632
rect 13256 16584 13308 16590
rect 13162 16552 13218 16561
rect 13256 16526 13308 16532
rect 14096 16538 14124 17598
rect 14176 17536 14228 17542
rect 14360 17536 14412 17542
rect 14228 17484 14308 17490
rect 14176 17478 14308 17484
rect 14360 17478 14412 17484
rect 14188 17462 14308 17478
rect 14280 17338 14308 17462
rect 14268 17332 14320 17338
rect 14268 17274 14320 17280
rect 14176 16992 14228 16998
rect 14176 16934 14228 16940
rect 14188 16726 14216 16934
rect 14176 16720 14228 16726
rect 14176 16662 14228 16668
rect 13162 16487 13218 16496
rect 12980 16448 13032 16454
rect 12980 16390 13032 16396
rect 12992 16250 13020 16390
rect 12980 16244 13032 16250
rect 12980 16186 13032 16192
rect 13176 15366 13204 16487
rect 13268 15910 13296 16526
rect 14096 16510 14216 16538
rect 14280 16522 14308 17274
rect 14372 17066 14400 17478
rect 14484 17436 14780 17456
rect 14540 17434 14564 17436
rect 14620 17434 14644 17436
rect 14700 17434 14724 17436
rect 14562 17382 14564 17434
rect 14626 17382 14638 17434
rect 14700 17382 14702 17434
rect 14540 17380 14564 17382
rect 14620 17380 14644 17382
rect 14700 17380 14724 17382
rect 14484 17360 14780 17380
rect 14636 17264 14688 17270
rect 14634 17232 14636 17241
rect 14688 17232 14690 17241
rect 14634 17167 14690 17176
rect 14360 17060 14412 17066
rect 14360 17002 14412 17008
rect 14084 16244 14136 16250
rect 14084 16186 14136 16192
rect 13440 16108 13492 16114
rect 13440 16050 13492 16056
rect 13256 15904 13308 15910
rect 13256 15846 13308 15852
rect 13164 15360 13216 15366
rect 13164 15302 13216 15308
rect 13164 13864 13216 13870
rect 13164 13806 13216 13812
rect 13176 13394 13204 13806
rect 13164 13388 13216 13394
rect 13164 13330 13216 13336
rect 13072 12980 13124 12986
rect 13072 12922 13124 12928
rect 12704 12300 12756 12306
rect 12704 12242 12756 12248
rect 12716 11762 12744 12242
rect 13084 11898 13112 12922
rect 13176 12170 13204 13330
rect 13268 12646 13296 15846
rect 13348 15360 13400 15366
rect 13348 15302 13400 15308
rect 13360 14006 13388 15302
rect 13348 14000 13400 14006
rect 13348 13942 13400 13948
rect 13452 13190 13480 16050
rect 14096 15706 14124 16186
rect 14188 15745 14216 16510
rect 14268 16516 14320 16522
rect 14268 16458 14320 16464
rect 14280 16114 14308 16458
rect 14372 16454 14400 17002
rect 14360 16448 14412 16454
rect 14360 16390 14412 16396
rect 14268 16108 14320 16114
rect 14268 16050 14320 16056
rect 14372 15978 14400 16390
rect 14484 16348 14780 16368
rect 14540 16346 14564 16348
rect 14620 16346 14644 16348
rect 14700 16346 14724 16348
rect 14562 16294 14564 16346
rect 14626 16294 14638 16346
rect 14700 16294 14702 16346
rect 14540 16292 14564 16294
rect 14620 16292 14644 16294
rect 14700 16292 14724 16294
rect 14484 16272 14780 16292
rect 14832 16250 14860 18686
rect 15568 18630 15596 19246
rect 15832 18828 15884 18834
rect 15832 18770 15884 18776
rect 15556 18624 15608 18630
rect 15556 18566 15608 18572
rect 15188 18080 15240 18086
rect 15188 18022 15240 18028
rect 15004 17740 15056 17746
rect 15004 17682 15056 17688
rect 14912 17604 14964 17610
rect 14912 17546 14964 17552
rect 14924 16726 14952 17546
rect 15016 16794 15044 17682
rect 15200 17678 15228 18022
rect 15568 17814 15596 18566
rect 15844 18426 15872 18770
rect 15832 18420 15884 18426
rect 15832 18362 15884 18368
rect 15556 17808 15608 17814
rect 15556 17750 15608 17756
rect 15188 17672 15240 17678
rect 15188 17614 15240 17620
rect 15200 17202 15228 17614
rect 15372 17536 15424 17542
rect 15372 17478 15424 17484
rect 15922 17504 15978 17513
rect 15384 17270 15412 17478
rect 15922 17439 15978 17448
rect 15936 17338 15964 17439
rect 15924 17332 15976 17338
rect 15924 17274 15976 17280
rect 15372 17264 15424 17270
rect 15372 17206 15424 17212
rect 15188 17196 15240 17202
rect 15188 17138 15240 17144
rect 15004 16788 15056 16794
rect 15004 16730 15056 16736
rect 14912 16720 14964 16726
rect 14912 16662 14964 16668
rect 14924 16561 14952 16662
rect 15004 16652 15056 16658
rect 15004 16594 15056 16600
rect 14910 16552 14966 16561
rect 14910 16487 14966 16496
rect 15016 16250 15044 16594
rect 14820 16244 14872 16250
rect 14820 16186 14872 16192
rect 15004 16244 15056 16250
rect 15004 16186 15056 16192
rect 15200 16114 15228 17138
rect 15648 17060 15700 17066
rect 15648 17002 15700 17008
rect 15660 16726 15688 17002
rect 16028 16726 16056 24550
rect 16580 24177 16608 27520
rect 17120 25152 17172 25158
rect 17120 25094 17172 25100
rect 16752 24268 16804 24274
rect 16752 24210 16804 24216
rect 16566 24168 16622 24177
rect 16566 24103 16622 24112
rect 16764 23526 16792 24210
rect 16292 23520 16344 23526
rect 16292 23462 16344 23468
rect 16752 23520 16804 23526
rect 16752 23462 16804 23468
rect 16304 23118 16332 23462
rect 16764 23254 16792 23462
rect 16752 23248 16804 23254
rect 16752 23190 16804 23196
rect 16292 23112 16344 23118
rect 16660 23112 16712 23118
rect 16292 23054 16344 23060
rect 16658 23080 16660 23089
rect 16712 23080 16714 23089
rect 16658 23015 16714 23024
rect 16672 22778 16700 23015
rect 16660 22772 16712 22778
rect 16660 22714 16712 22720
rect 16764 22658 16792 23190
rect 16672 22630 16792 22658
rect 16672 22438 16700 22630
rect 16660 22432 16712 22438
rect 16660 22374 16712 22380
rect 16384 20936 16436 20942
rect 16384 20878 16436 20884
rect 16396 20330 16424 20878
rect 16672 20602 16700 22374
rect 16752 21072 16804 21078
rect 16752 21014 16804 21020
rect 16660 20596 16712 20602
rect 16660 20538 16712 20544
rect 16764 20398 16792 21014
rect 16752 20392 16804 20398
rect 16752 20334 16804 20340
rect 16200 20324 16252 20330
rect 16200 20266 16252 20272
rect 16384 20324 16436 20330
rect 16384 20266 16436 20272
rect 16212 19514 16240 20266
rect 16396 19990 16424 20266
rect 16764 19990 16792 20334
rect 16384 19984 16436 19990
rect 16384 19926 16436 19932
rect 16752 19984 16804 19990
rect 16752 19926 16804 19932
rect 16476 19848 16528 19854
rect 16476 19790 16528 19796
rect 16200 19508 16252 19514
rect 16200 19450 16252 19456
rect 16488 19310 16516 19790
rect 16752 19508 16804 19514
rect 16752 19450 16804 19456
rect 16764 19378 16792 19450
rect 16752 19372 16804 19378
rect 16752 19314 16804 19320
rect 16476 19304 16528 19310
rect 16476 19246 16528 19252
rect 16568 18760 16620 18766
rect 16568 18702 16620 18708
rect 16580 18426 16608 18702
rect 16108 18420 16160 18426
rect 16108 18362 16160 18368
rect 16568 18420 16620 18426
rect 16568 18362 16620 18368
rect 16120 17882 16148 18362
rect 16200 18080 16252 18086
rect 16200 18022 16252 18028
rect 16108 17876 16160 17882
rect 16108 17818 16160 17824
rect 16212 17270 16240 18022
rect 16384 17740 16436 17746
rect 16384 17682 16436 17688
rect 16396 17270 16424 17682
rect 16200 17264 16252 17270
rect 16198 17232 16200 17241
rect 16384 17264 16436 17270
rect 16252 17232 16254 17241
rect 16384 17206 16436 17212
rect 16198 17167 16254 17176
rect 15648 16720 15700 16726
rect 15648 16662 15700 16668
rect 16016 16720 16068 16726
rect 16016 16662 16068 16668
rect 16200 16720 16252 16726
rect 16200 16662 16252 16668
rect 15188 16108 15240 16114
rect 15188 16050 15240 16056
rect 14360 15972 14412 15978
rect 14360 15914 14412 15920
rect 14174 15736 14230 15745
rect 14084 15700 14136 15706
rect 14174 15671 14230 15680
rect 14084 15642 14136 15648
rect 14372 15366 14400 15914
rect 15200 15910 15228 16050
rect 15188 15904 15240 15910
rect 15108 15852 15188 15858
rect 15108 15846 15240 15852
rect 15108 15830 15228 15846
rect 14912 15496 14964 15502
rect 14912 15438 14964 15444
rect 14360 15360 14412 15366
rect 14360 15302 14412 15308
rect 14372 14958 14400 15302
rect 14484 15260 14780 15280
rect 14540 15258 14564 15260
rect 14620 15258 14644 15260
rect 14700 15258 14724 15260
rect 14562 15206 14564 15258
rect 14626 15206 14638 15258
rect 14700 15206 14702 15258
rect 14540 15204 14564 15206
rect 14620 15204 14644 15206
rect 14700 15204 14724 15206
rect 14484 15184 14780 15204
rect 14360 14952 14412 14958
rect 14360 14894 14412 14900
rect 14636 14952 14688 14958
rect 14636 14894 14688 14900
rect 13900 14816 13952 14822
rect 13900 14758 13952 14764
rect 13912 14618 13940 14758
rect 13900 14612 13952 14618
rect 13900 14554 13952 14560
rect 14372 14074 14400 14894
rect 14648 14482 14676 14894
rect 14924 14890 14952 15438
rect 15004 14952 15056 14958
rect 15004 14894 15056 14900
rect 14912 14884 14964 14890
rect 14912 14826 14964 14832
rect 14924 14618 14952 14826
rect 14912 14612 14964 14618
rect 14912 14554 14964 14560
rect 15016 14482 15044 14894
rect 14636 14476 14688 14482
rect 14636 14418 14688 14424
rect 15004 14476 15056 14482
rect 15004 14418 15056 14424
rect 14484 14172 14780 14192
rect 14540 14170 14564 14172
rect 14620 14170 14644 14172
rect 14700 14170 14724 14172
rect 14562 14118 14564 14170
rect 14626 14118 14638 14170
rect 14700 14118 14702 14170
rect 14540 14116 14564 14118
rect 14620 14116 14644 14118
rect 14700 14116 14724 14118
rect 14484 14096 14780 14116
rect 14360 14068 14412 14074
rect 14360 14010 14412 14016
rect 14268 14000 14320 14006
rect 14268 13942 14320 13948
rect 14280 13870 14308 13942
rect 15016 13870 15044 14418
rect 14084 13864 14136 13870
rect 14084 13806 14136 13812
rect 14268 13864 14320 13870
rect 14268 13806 14320 13812
rect 14728 13864 14780 13870
rect 14728 13806 14780 13812
rect 15004 13864 15056 13870
rect 15004 13806 15056 13812
rect 13900 13456 13952 13462
rect 13898 13424 13900 13433
rect 13952 13424 13954 13433
rect 13898 13359 13954 13368
rect 13532 13320 13584 13326
rect 13532 13262 13584 13268
rect 13440 13184 13492 13190
rect 13440 13126 13492 13132
rect 13452 12986 13480 13126
rect 13440 12980 13492 12986
rect 13440 12922 13492 12928
rect 13544 12646 13572 13262
rect 13808 13184 13860 13190
rect 13808 13126 13860 13132
rect 13820 12782 13848 13126
rect 13900 12980 13952 12986
rect 13900 12922 13952 12928
rect 13808 12776 13860 12782
rect 13808 12718 13860 12724
rect 13256 12640 13308 12646
rect 13256 12582 13308 12588
rect 13532 12640 13584 12646
rect 13532 12582 13584 12588
rect 13268 12442 13296 12582
rect 13256 12436 13308 12442
rect 13256 12378 13308 12384
rect 13716 12300 13768 12306
rect 13716 12242 13768 12248
rect 13164 12164 13216 12170
rect 13164 12106 13216 12112
rect 13072 11892 13124 11898
rect 13072 11834 13124 11840
rect 12704 11756 12756 11762
rect 12704 11698 12756 11704
rect 13624 11620 13676 11626
rect 13624 11562 13676 11568
rect 13532 11076 13584 11082
rect 13532 11018 13584 11024
rect 13348 10804 13400 10810
rect 13348 10746 13400 10752
rect 13360 9926 13388 10746
rect 13544 10130 13572 11018
rect 13636 10470 13664 11562
rect 13728 11558 13756 12242
rect 13820 11626 13848 12718
rect 13912 12322 13940 12922
rect 13912 12294 14032 12322
rect 14004 12238 14032 12294
rect 13992 12232 14044 12238
rect 13992 12174 14044 12180
rect 14004 11694 14032 12174
rect 14096 12102 14124 13806
rect 14740 13394 14768 13806
rect 14728 13388 14780 13394
rect 14780 13348 14860 13376
rect 14728 13330 14780 13336
rect 14358 13288 14414 13297
rect 14358 13223 14414 13232
rect 14268 13184 14320 13190
rect 14268 13126 14320 13132
rect 14280 12986 14308 13126
rect 14372 12986 14400 13223
rect 14484 13084 14780 13104
rect 14540 13082 14564 13084
rect 14620 13082 14644 13084
rect 14700 13082 14724 13084
rect 14562 13030 14564 13082
rect 14626 13030 14638 13082
rect 14700 13030 14702 13082
rect 14540 13028 14564 13030
rect 14620 13028 14644 13030
rect 14700 13028 14724 13030
rect 14484 13008 14780 13028
rect 14832 12986 14860 13348
rect 15016 13326 15044 13806
rect 15004 13320 15056 13326
rect 14924 13268 15004 13274
rect 14924 13262 15056 13268
rect 14924 13246 15044 13262
rect 14268 12980 14320 12986
rect 14268 12922 14320 12928
rect 14360 12980 14412 12986
rect 14360 12922 14412 12928
rect 14820 12980 14872 12986
rect 14820 12922 14872 12928
rect 14176 12912 14228 12918
rect 14176 12854 14228 12860
rect 14188 12442 14216 12854
rect 14924 12442 14952 13246
rect 15108 13138 15136 15830
rect 15740 15632 15792 15638
rect 16028 15620 16056 16662
rect 16212 16046 16240 16662
rect 16200 16040 16252 16046
rect 16200 15982 16252 15988
rect 16212 15706 16240 15982
rect 16200 15700 16252 15706
rect 16200 15642 16252 15648
rect 16108 15632 16160 15638
rect 16028 15592 16108 15620
rect 15740 15574 15792 15580
rect 16108 15574 16160 15580
rect 15752 15162 15780 15574
rect 16764 15570 16792 19314
rect 16844 17536 16896 17542
rect 16844 17478 16896 17484
rect 16856 17202 16884 17478
rect 16844 17196 16896 17202
rect 16844 17138 16896 17144
rect 16752 15564 16804 15570
rect 16752 15506 16804 15512
rect 16660 15496 16712 15502
rect 16660 15438 16712 15444
rect 15740 15156 15792 15162
rect 15568 15116 15740 15144
rect 15188 14952 15240 14958
rect 15188 14894 15240 14900
rect 15200 14550 15228 14894
rect 15464 14816 15516 14822
rect 15464 14758 15516 14764
rect 15476 14618 15504 14758
rect 15464 14612 15516 14618
rect 15464 14554 15516 14560
rect 15188 14544 15240 14550
rect 15188 14486 15240 14492
rect 15200 13394 15228 14486
rect 15464 13728 15516 13734
rect 15464 13670 15516 13676
rect 15476 13530 15504 13670
rect 15464 13524 15516 13530
rect 15464 13466 15516 13472
rect 15188 13388 15240 13394
rect 15188 13330 15240 13336
rect 15016 13110 15136 13138
rect 14176 12436 14228 12442
rect 14176 12378 14228 12384
rect 14912 12436 14964 12442
rect 14912 12378 14964 12384
rect 14176 12300 14228 12306
rect 14176 12242 14228 12248
rect 14820 12300 14872 12306
rect 14820 12242 14872 12248
rect 14084 12096 14136 12102
rect 14084 12038 14136 12044
rect 13992 11688 14044 11694
rect 13992 11630 14044 11636
rect 13808 11620 13860 11626
rect 13808 11562 13860 11568
rect 13716 11552 13768 11558
rect 13714 11520 13716 11529
rect 13768 11520 13770 11529
rect 13714 11455 13770 11464
rect 13820 11150 13848 11562
rect 14004 11286 14032 11630
rect 14096 11354 14124 12038
rect 14084 11348 14136 11354
rect 14084 11290 14136 11296
rect 13992 11280 14044 11286
rect 13992 11222 14044 11228
rect 13808 11144 13860 11150
rect 13808 11086 13860 11092
rect 13624 10464 13676 10470
rect 13624 10406 13676 10412
rect 13532 10124 13584 10130
rect 13532 10066 13584 10072
rect 13348 9920 13400 9926
rect 13348 9862 13400 9868
rect 12612 9716 12664 9722
rect 12612 9658 12664 9664
rect 12336 9444 12388 9450
rect 12336 9386 12388 9392
rect 12348 9110 12376 9386
rect 13544 9382 13572 10066
rect 13532 9376 13584 9382
rect 13532 9318 13584 9324
rect 12336 9104 12388 9110
rect 12242 9072 12298 9081
rect 12336 9046 12388 9052
rect 12242 9007 12298 9016
rect 13256 9036 13308 9042
rect 13256 8978 13308 8984
rect 12888 8900 12940 8906
rect 12888 8842 12940 8848
rect 12900 8634 12928 8842
rect 12888 8628 12940 8634
rect 12888 8570 12940 8576
rect 13268 8362 13296 8978
rect 13544 8974 13572 9318
rect 13532 8968 13584 8974
rect 13532 8910 13584 8916
rect 13544 8634 13572 8910
rect 13636 8838 13664 10406
rect 13716 9512 13768 9518
rect 13716 9454 13768 9460
rect 13728 9042 13756 9454
rect 13716 9036 13768 9042
rect 13716 8978 13768 8984
rect 13624 8832 13676 8838
rect 13624 8774 13676 8780
rect 13532 8628 13584 8634
rect 13532 8570 13584 8576
rect 13636 8498 13664 8774
rect 13624 8492 13676 8498
rect 13624 8434 13676 8440
rect 13256 8356 13308 8362
rect 13256 8298 13308 8304
rect 13268 8090 13296 8298
rect 13438 8256 13494 8265
rect 13438 8191 13494 8200
rect 13256 8084 13308 8090
rect 13256 8026 13308 8032
rect 12244 7336 12296 7342
rect 12244 7278 12296 7284
rect 12060 7268 12112 7274
rect 12060 7210 12112 7216
rect 11782 7168 11838 7177
rect 11782 7103 11838 7112
rect 11046 6896 11102 6905
rect 11046 6831 11102 6840
rect 11600 6792 11652 6798
rect 11600 6734 11652 6740
rect 11612 6118 11640 6734
rect 11600 6112 11652 6118
rect 11600 6054 11652 6060
rect 11612 5817 11640 6054
rect 11598 5808 11654 5817
rect 11598 5743 11654 5752
rect 10770 4040 10826 4049
rect 10770 3975 10826 3984
rect 10586 3496 10642 3505
rect 10586 3431 10642 3440
rect 9817 2748 10113 2768
rect 9873 2746 9897 2748
rect 9953 2746 9977 2748
rect 10033 2746 10057 2748
rect 9895 2694 9897 2746
rect 9959 2694 9971 2746
rect 10033 2694 10035 2746
rect 9873 2692 9897 2694
rect 9953 2692 9977 2694
rect 10033 2692 10057 2694
rect 9817 2672 10113 2692
rect 11796 480 11824 7103
rect 11876 6860 11928 6866
rect 11876 6802 11928 6808
rect 11888 6254 11916 6802
rect 12072 6458 12100 7210
rect 12256 6866 12284 7278
rect 13452 6866 13480 8191
rect 13636 7478 13664 8434
rect 13820 8294 13848 11086
rect 13900 10600 13952 10606
rect 13900 10542 13952 10548
rect 13912 10198 13940 10542
rect 13900 10192 13952 10198
rect 13900 10134 13952 10140
rect 14004 9466 14032 11222
rect 14084 11212 14136 11218
rect 14084 11154 14136 11160
rect 14096 10810 14124 11154
rect 14084 10804 14136 10810
rect 14084 10746 14136 10752
rect 14096 10266 14124 10746
rect 14084 10260 14136 10266
rect 14084 10202 14136 10208
rect 14096 9586 14124 10202
rect 14084 9580 14136 9586
rect 14084 9522 14136 9528
rect 14004 9438 14124 9466
rect 13808 8288 13860 8294
rect 13808 8230 13860 8236
rect 13624 7472 13676 7478
rect 13624 7414 13676 7420
rect 13636 7206 13664 7414
rect 13820 7274 13848 8230
rect 14096 7342 14124 9438
rect 14188 9178 14216 12242
rect 14360 12096 14412 12102
rect 14360 12038 14412 12044
rect 14372 11830 14400 12038
rect 14484 11996 14780 12016
rect 14540 11994 14564 11996
rect 14620 11994 14644 11996
rect 14700 11994 14724 11996
rect 14562 11942 14564 11994
rect 14626 11942 14638 11994
rect 14700 11942 14702 11994
rect 14540 11940 14564 11942
rect 14620 11940 14644 11942
rect 14700 11940 14724 11942
rect 14484 11920 14780 11940
rect 14832 11898 14860 12242
rect 14820 11892 14872 11898
rect 14820 11834 14872 11840
rect 14360 11824 14412 11830
rect 14360 11766 14412 11772
rect 14268 11756 14320 11762
rect 14268 11698 14320 11704
rect 14280 11082 14308 11698
rect 14360 11552 14412 11558
rect 14360 11494 14412 11500
rect 14268 11076 14320 11082
rect 14268 11018 14320 11024
rect 14372 10713 14400 11494
rect 14820 11348 14872 11354
rect 14820 11290 14872 11296
rect 14832 11218 14860 11290
rect 14820 11212 14872 11218
rect 14820 11154 14872 11160
rect 14484 10908 14780 10928
rect 14540 10906 14564 10908
rect 14620 10906 14644 10908
rect 14700 10906 14724 10908
rect 14562 10854 14564 10906
rect 14626 10854 14638 10906
rect 14700 10854 14702 10906
rect 14540 10852 14564 10854
rect 14620 10852 14644 10854
rect 14700 10852 14724 10854
rect 14484 10832 14780 10852
rect 14358 10704 14414 10713
rect 14358 10639 14414 10648
rect 14636 10464 14688 10470
rect 14832 10418 14860 11154
rect 15016 10810 15044 13110
rect 15476 12850 15504 13466
rect 15568 12986 15596 15116
rect 15740 15098 15792 15104
rect 16672 14618 16700 15438
rect 16764 15162 16792 15506
rect 16752 15156 16804 15162
rect 16752 15098 16804 15104
rect 16660 14612 16712 14618
rect 16660 14554 16712 14560
rect 16764 14550 16792 15098
rect 17132 14770 17160 25094
rect 17592 24449 17620 27520
rect 18498 24848 18554 24857
rect 18498 24783 18554 24792
rect 18040 24608 18092 24614
rect 18040 24550 18092 24556
rect 17578 24440 17634 24449
rect 17578 24375 17634 24384
rect 17212 24064 17264 24070
rect 17212 24006 17264 24012
rect 17764 24064 17816 24070
rect 17764 24006 17816 24012
rect 17224 22778 17252 24006
rect 17776 23594 17804 24006
rect 17764 23588 17816 23594
rect 17764 23530 17816 23536
rect 17396 23520 17448 23526
rect 17396 23462 17448 23468
rect 17304 23112 17356 23118
rect 17304 23054 17356 23060
rect 17212 22772 17264 22778
rect 17212 22714 17264 22720
rect 17224 22438 17252 22714
rect 17316 22642 17344 23054
rect 17304 22636 17356 22642
rect 17304 22578 17356 22584
rect 17212 22432 17264 22438
rect 17212 22374 17264 22380
rect 17408 22098 17436 23462
rect 17776 23118 17804 23530
rect 18052 23118 18080 24550
rect 18512 24410 18540 24783
rect 18500 24404 18552 24410
rect 18500 24346 18552 24352
rect 18604 24313 18632 27520
rect 19150 25596 19446 25616
rect 19206 25594 19230 25596
rect 19286 25594 19310 25596
rect 19366 25594 19390 25596
rect 19228 25542 19230 25594
rect 19292 25542 19304 25594
rect 19366 25542 19368 25594
rect 19206 25540 19230 25542
rect 19286 25540 19310 25542
rect 19366 25540 19390 25542
rect 19150 25520 19446 25540
rect 19616 24721 19644 27520
rect 20720 24857 20748 27520
rect 20800 25356 20852 25362
rect 20800 25298 20852 25304
rect 20812 24954 20840 25298
rect 20800 24948 20852 24954
rect 20800 24890 20852 24896
rect 20706 24848 20762 24857
rect 20706 24783 20762 24792
rect 20156 24744 20208 24750
rect 19602 24712 19658 24721
rect 20156 24686 20208 24692
rect 19602 24647 19658 24656
rect 19150 24508 19446 24528
rect 19206 24506 19230 24508
rect 19286 24506 19310 24508
rect 19366 24506 19390 24508
rect 19228 24454 19230 24506
rect 19292 24454 19304 24506
rect 19366 24454 19368 24506
rect 19206 24452 19230 24454
rect 19286 24452 19310 24454
rect 19366 24452 19390 24454
rect 19150 24432 19446 24452
rect 18590 24304 18646 24313
rect 18316 24268 18368 24274
rect 18590 24239 18646 24248
rect 18316 24210 18368 24216
rect 18328 23798 18356 24210
rect 19694 23896 19750 23905
rect 19694 23831 19696 23840
rect 19748 23831 19750 23840
rect 19696 23802 19748 23808
rect 18316 23792 18368 23798
rect 18316 23734 18368 23740
rect 20168 23610 20196 24686
rect 20524 24676 20576 24682
rect 20524 24618 20576 24624
rect 20536 24342 20564 24618
rect 20524 24336 20576 24342
rect 20524 24278 20576 24284
rect 20614 24304 20670 24313
rect 20536 23866 20564 24278
rect 20614 24239 20670 24248
rect 20628 24206 20656 24239
rect 20616 24200 20668 24206
rect 20812 24177 20840 24890
rect 21352 24744 21404 24750
rect 21352 24686 21404 24692
rect 20616 24142 20668 24148
rect 20798 24168 20854 24177
rect 20524 23860 20576 23866
rect 20524 23802 20576 23808
rect 18500 23588 18552 23594
rect 20168 23582 20288 23610
rect 18500 23530 18552 23536
rect 18224 23248 18276 23254
rect 18144 23196 18224 23202
rect 18144 23190 18276 23196
rect 18144 23174 18264 23190
rect 17764 23112 17816 23118
rect 17670 23080 17726 23089
rect 17764 23054 17816 23060
rect 18040 23112 18092 23118
rect 18040 23054 18092 23060
rect 17670 23015 17672 23024
rect 17724 23015 17726 23024
rect 17672 22986 17724 22992
rect 17684 22506 17712 22986
rect 18052 22778 18080 23054
rect 18040 22772 18092 22778
rect 18040 22714 18092 22720
rect 17672 22500 17724 22506
rect 17672 22442 17724 22448
rect 18144 22438 18172 23174
rect 18512 23118 18540 23530
rect 19512 23520 19564 23526
rect 19512 23462 19564 23468
rect 20156 23520 20208 23526
rect 20156 23462 20208 23468
rect 19150 23420 19446 23440
rect 19206 23418 19230 23420
rect 19286 23418 19310 23420
rect 19366 23418 19390 23420
rect 19228 23366 19230 23418
rect 19292 23366 19304 23418
rect 19366 23366 19368 23418
rect 19206 23364 19230 23366
rect 19286 23364 19310 23366
rect 19366 23364 19390 23366
rect 19150 23344 19446 23364
rect 18500 23112 18552 23118
rect 18500 23054 18552 23060
rect 18512 22574 18540 23054
rect 19524 22778 19552 23462
rect 19512 22772 19564 22778
rect 19512 22714 19564 22720
rect 18500 22568 18552 22574
rect 18500 22510 18552 22516
rect 18132 22432 18184 22438
rect 18132 22374 18184 22380
rect 18144 22166 18172 22374
rect 19150 22332 19446 22352
rect 19206 22330 19230 22332
rect 19286 22330 19310 22332
rect 19366 22330 19390 22332
rect 19228 22278 19230 22330
rect 19292 22278 19304 22330
rect 19366 22278 19368 22330
rect 19206 22276 19230 22278
rect 19286 22276 19310 22278
rect 19366 22276 19390 22278
rect 19150 22256 19446 22276
rect 18132 22160 18184 22166
rect 18132 22102 18184 22108
rect 17396 22092 17448 22098
rect 17396 22034 17448 22040
rect 17764 22092 17816 22098
rect 17764 22034 17816 22040
rect 17776 21690 17804 22034
rect 18500 21888 18552 21894
rect 18500 21830 18552 21836
rect 17764 21684 17816 21690
rect 17764 21626 17816 21632
rect 17776 21146 17804 21626
rect 18512 21418 18540 21830
rect 18960 21548 19012 21554
rect 18960 21490 19012 21496
rect 18590 21448 18646 21457
rect 18500 21412 18552 21418
rect 18590 21383 18592 21392
rect 18500 21354 18552 21360
rect 18644 21383 18646 21392
rect 18592 21354 18644 21360
rect 17764 21140 17816 21146
rect 17764 21082 17816 21088
rect 18512 21049 18540 21354
rect 18868 21072 18920 21078
rect 18498 21040 18554 21049
rect 18868 21014 18920 21020
rect 18498 20975 18554 20984
rect 17672 20800 17724 20806
rect 17672 20742 17724 20748
rect 17684 20641 17712 20742
rect 17670 20632 17726 20641
rect 17670 20567 17726 20576
rect 17684 20312 17712 20567
rect 18592 20460 18644 20466
rect 18592 20402 18644 20408
rect 17764 20324 17816 20330
rect 17684 20284 17764 20312
rect 17580 20256 17632 20262
rect 17580 20198 17632 20204
rect 17592 19938 17620 20198
rect 17684 20058 17712 20284
rect 17764 20266 17816 20272
rect 18500 20256 18552 20262
rect 18500 20198 18552 20204
rect 17672 20052 17724 20058
rect 17672 19994 17724 20000
rect 17670 19952 17726 19961
rect 17592 19910 17670 19938
rect 17670 19887 17672 19896
rect 17724 19887 17726 19896
rect 17672 19858 17724 19864
rect 17580 19304 17632 19310
rect 17580 19246 17632 19252
rect 17592 18902 17620 19246
rect 18512 18970 18540 20198
rect 18604 20058 18632 20402
rect 18592 20052 18644 20058
rect 18592 19994 18644 20000
rect 18880 19922 18908 21014
rect 18972 20942 19000 21490
rect 20168 21486 20196 23462
rect 20260 22166 20288 23582
rect 20628 23322 20656 24142
rect 20798 24103 20854 24112
rect 20800 24064 20852 24070
rect 20800 24006 20852 24012
rect 20812 23730 20840 24006
rect 20800 23724 20852 23730
rect 20800 23666 20852 23672
rect 20616 23316 20668 23322
rect 20616 23258 20668 23264
rect 20708 22976 20760 22982
rect 20708 22918 20760 22924
rect 20720 22506 20748 22918
rect 20708 22500 20760 22506
rect 20708 22442 20760 22448
rect 20616 22432 20668 22438
rect 20616 22374 20668 22380
rect 20248 22160 20300 22166
rect 20248 22102 20300 22108
rect 20156 21480 20208 21486
rect 20156 21422 20208 21428
rect 20260 21350 20288 22102
rect 20524 22024 20576 22030
rect 20522 21992 20524 22001
rect 20576 21992 20578 22001
rect 20522 21927 20578 21936
rect 20536 21622 20564 21927
rect 20628 21690 20656 22374
rect 20720 22234 20748 22442
rect 20708 22228 20760 22234
rect 20708 22170 20760 22176
rect 20812 22030 20840 23666
rect 21364 23594 21392 24686
rect 21352 23588 21404 23594
rect 21352 23530 21404 23536
rect 21364 22642 21392 23530
rect 21444 23248 21496 23254
rect 21442 23216 21444 23225
rect 21628 23248 21680 23254
rect 21496 23216 21498 23225
rect 21628 23190 21680 23196
rect 21442 23151 21498 23160
rect 21456 22710 21484 23151
rect 21640 22778 21668 23190
rect 21628 22772 21680 22778
rect 21628 22714 21680 22720
rect 21444 22704 21496 22710
rect 21444 22646 21496 22652
rect 21352 22636 21404 22642
rect 21352 22578 21404 22584
rect 20800 22024 20852 22030
rect 20800 21966 20852 21972
rect 20616 21684 20668 21690
rect 20616 21626 20668 21632
rect 20524 21616 20576 21622
rect 20524 21558 20576 21564
rect 20708 21480 20760 21486
rect 20430 21448 20486 21457
rect 20708 21422 20760 21428
rect 21640 21434 21668 22714
rect 21732 21690 21760 27520
rect 21996 25152 22048 25158
rect 21996 25094 22048 25100
rect 21812 24608 21864 24614
rect 21812 24550 21864 24556
rect 21824 24274 21852 24550
rect 21812 24268 21864 24274
rect 21812 24210 21864 24216
rect 21824 23866 21852 24210
rect 21812 23860 21864 23866
rect 21812 23802 21864 23808
rect 21720 21684 21772 21690
rect 21720 21626 21772 21632
rect 20430 21383 20486 21392
rect 20248 21344 20300 21350
rect 20168 21304 20248 21332
rect 19150 21244 19446 21264
rect 19206 21242 19230 21244
rect 19286 21242 19310 21244
rect 19366 21242 19390 21244
rect 19228 21190 19230 21242
rect 19292 21190 19304 21242
rect 19366 21190 19368 21242
rect 19206 21188 19230 21190
rect 19286 21188 19310 21190
rect 19366 21188 19390 21190
rect 19150 21168 19446 21188
rect 18960 20936 19012 20942
rect 18960 20878 19012 20884
rect 19512 20936 19564 20942
rect 19512 20878 19564 20884
rect 18972 20466 19000 20878
rect 19524 20466 19552 20878
rect 18960 20460 19012 20466
rect 18960 20402 19012 20408
rect 19512 20460 19564 20466
rect 19512 20402 19564 20408
rect 18960 20256 19012 20262
rect 18960 20198 19012 20204
rect 18972 20058 19000 20198
rect 19150 20156 19446 20176
rect 19206 20154 19230 20156
rect 19286 20154 19310 20156
rect 19366 20154 19390 20156
rect 19228 20102 19230 20154
rect 19292 20102 19304 20154
rect 19366 20102 19368 20154
rect 19206 20100 19230 20102
rect 19286 20100 19310 20102
rect 19366 20100 19390 20102
rect 19150 20080 19446 20100
rect 18960 20052 19012 20058
rect 18960 19994 19012 20000
rect 19524 19922 19552 20402
rect 18868 19916 18920 19922
rect 18868 19858 18920 19864
rect 19512 19916 19564 19922
rect 19512 19858 19564 19864
rect 18880 19514 18908 19858
rect 18868 19508 18920 19514
rect 18868 19450 18920 19456
rect 18880 19310 18908 19450
rect 18868 19304 18920 19310
rect 18868 19246 18920 19252
rect 19788 19304 19840 19310
rect 19788 19246 19840 19252
rect 18960 19236 19012 19242
rect 18960 19178 19012 19184
rect 18500 18964 18552 18970
rect 18500 18906 18552 18912
rect 17580 18896 17632 18902
rect 17580 18838 17632 18844
rect 18868 18828 18920 18834
rect 18868 18770 18920 18776
rect 18224 18216 18276 18222
rect 18224 18158 18276 18164
rect 17856 17536 17908 17542
rect 17856 17478 17908 17484
rect 17212 17264 17264 17270
rect 17212 17206 17264 17212
rect 17224 15162 17252 17206
rect 17868 17202 17896 17478
rect 18236 17270 18264 18158
rect 18880 18086 18908 18770
rect 18972 18426 19000 19178
rect 19150 19068 19446 19088
rect 19206 19066 19230 19068
rect 19286 19066 19310 19068
rect 19366 19066 19390 19068
rect 19228 19014 19230 19066
rect 19292 19014 19304 19066
rect 19366 19014 19368 19066
rect 19206 19012 19230 19014
rect 19286 19012 19310 19014
rect 19366 19012 19390 19014
rect 19150 18992 19446 19012
rect 19800 18902 19828 19246
rect 19788 18896 19840 18902
rect 19788 18838 19840 18844
rect 19052 18828 19104 18834
rect 19052 18770 19104 18776
rect 18960 18420 19012 18426
rect 18960 18362 19012 18368
rect 18972 18154 19000 18362
rect 18960 18148 19012 18154
rect 18960 18090 19012 18096
rect 19064 18086 19092 18770
rect 20168 18426 20196 21304
rect 20248 21286 20300 21292
rect 20444 21078 20472 21383
rect 20432 21072 20484 21078
rect 20432 21014 20484 21020
rect 20524 21004 20576 21010
rect 20524 20946 20576 20952
rect 20536 20641 20564 20946
rect 20522 20632 20578 20641
rect 20522 20567 20524 20576
rect 20576 20567 20578 20576
rect 20524 20538 20576 20544
rect 20536 20507 20564 20538
rect 20720 19310 20748 21422
rect 21640 21406 21760 21434
rect 21628 21344 21680 21350
rect 21548 21292 21628 21298
rect 21548 21286 21680 21292
rect 21548 21270 21668 21286
rect 21168 20392 21220 20398
rect 21168 20334 21220 20340
rect 21076 20256 21128 20262
rect 21076 20198 21128 20204
rect 21088 19990 21116 20198
rect 21076 19984 21128 19990
rect 21076 19926 21128 19932
rect 20984 19916 21036 19922
rect 20984 19858 21036 19864
rect 20996 19514 21024 19858
rect 20984 19508 21036 19514
rect 20984 19450 21036 19456
rect 20708 19304 20760 19310
rect 20708 19246 20760 19252
rect 21088 19242 21116 19926
rect 21180 19718 21208 20334
rect 21548 20058 21576 21270
rect 21732 20602 21760 21406
rect 22008 20890 22036 25094
rect 22270 24440 22326 24449
rect 22270 24375 22272 24384
rect 22324 24375 22326 24384
rect 22272 24346 22324 24352
rect 22640 24268 22692 24274
rect 22640 24210 22692 24216
rect 22652 23866 22680 24210
rect 22744 23905 22772 27520
rect 23756 24449 23784 27520
rect 24294 26344 24350 26353
rect 24294 26279 24350 26288
rect 23817 25052 24113 25072
rect 23873 25050 23897 25052
rect 23953 25050 23977 25052
rect 24033 25050 24057 25052
rect 23895 24998 23897 25050
rect 23959 24998 23971 25050
rect 24033 24998 24035 25050
rect 23873 24996 23897 24998
rect 23953 24996 23977 24998
rect 24033 24996 24057 24998
rect 23817 24976 24113 24996
rect 24308 24818 24336 26279
rect 24570 25392 24626 25401
rect 24570 25327 24626 25336
rect 24296 24812 24348 24818
rect 24296 24754 24348 24760
rect 24204 24608 24256 24614
rect 24204 24550 24256 24556
rect 23742 24440 23798 24449
rect 23742 24375 23798 24384
rect 23817 23964 24113 23984
rect 23873 23962 23897 23964
rect 23953 23962 23977 23964
rect 24033 23962 24057 23964
rect 23895 23910 23897 23962
rect 23959 23910 23971 23962
rect 24033 23910 24035 23962
rect 23873 23908 23897 23910
rect 23953 23908 23977 23910
rect 24033 23908 24057 23910
rect 22730 23896 22786 23905
rect 22640 23860 22692 23866
rect 23817 23888 24113 23908
rect 22730 23831 22786 23840
rect 22640 23802 22692 23808
rect 23008 23656 23060 23662
rect 23008 23598 23060 23604
rect 23020 23338 23048 23598
rect 23192 23588 23244 23594
rect 23192 23530 23244 23536
rect 22928 23322 23048 23338
rect 22916 23316 23048 23322
rect 22968 23310 23048 23316
rect 22916 23258 22968 23264
rect 23204 23254 23232 23530
rect 24216 23322 24244 24550
rect 24478 24304 24534 24313
rect 24296 24268 24348 24274
rect 24584 24274 24612 25327
rect 24860 24410 24888 27520
rect 25398 27432 25454 27441
rect 25398 27367 25454 27376
rect 25412 24818 25440 27367
rect 25400 24812 25452 24818
rect 25400 24754 25452 24760
rect 25032 24608 25084 24614
rect 25032 24550 25084 24556
rect 24848 24404 24900 24410
rect 24848 24346 24900 24352
rect 24478 24239 24534 24248
rect 24572 24268 24624 24274
rect 24296 24210 24348 24216
rect 24308 24154 24336 24210
rect 24308 24126 24428 24154
rect 24492 24138 24520 24239
rect 24572 24210 24624 24216
rect 24294 23488 24350 23497
rect 24294 23423 24350 23432
rect 24204 23316 24256 23322
rect 24204 23258 24256 23264
rect 23192 23248 23244 23254
rect 23192 23190 23244 23196
rect 23204 22778 23232 23190
rect 23284 23112 23336 23118
rect 23284 23054 23336 23060
rect 23192 22772 23244 22778
rect 23192 22714 23244 22720
rect 23296 22642 23324 23054
rect 23817 22876 24113 22896
rect 23873 22874 23897 22876
rect 23953 22874 23977 22876
rect 24033 22874 24057 22876
rect 23895 22822 23897 22874
rect 23959 22822 23971 22874
rect 24033 22822 24035 22874
rect 23873 22820 23897 22822
rect 23953 22820 23977 22822
rect 24033 22820 24057 22822
rect 23817 22800 24113 22820
rect 24216 22778 24244 23258
rect 24204 22772 24256 22778
rect 24204 22714 24256 22720
rect 23284 22636 23336 22642
rect 23284 22578 23336 22584
rect 23560 22636 23612 22642
rect 23560 22578 23612 22584
rect 23192 22432 23244 22438
rect 23192 22374 23244 22380
rect 23008 22160 23060 22166
rect 23008 22102 23060 22108
rect 23204 22114 23232 22374
rect 23296 22234 23324 22578
rect 23284 22228 23336 22234
rect 23284 22170 23336 22176
rect 23572 22166 23600 22578
rect 23560 22160 23612 22166
rect 22548 22024 22600 22030
rect 22548 21966 22600 21972
rect 22560 21690 22588 21966
rect 22548 21684 22600 21690
rect 22548 21626 22600 21632
rect 22560 21146 22588 21626
rect 23020 21554 23048 22102
rect 23204 22086 23324 22114
rect 23560 22102 23612 22108
rect 23008 21548 23060 21554
rect 23008 21490 23060 21496
rect 23296 21486 23324 22086
rect 23817 21788 24113 21808
rect 23873 21786 23897 21788
rect 23953 21786 23977 21788
rect 24033 21786 24057 21788
rect 23895 21734 23897 21786
rect 23959 21734 23971 21786
rect 24033 21734 24035 21786
rect 23873 21732 23897 21734
rect 23953 21732 23977 21734
rect 24033 21732 24057 21734
rect 23817 21712 24113 21732
rect 23284 21480 23336 21486
rect 23284 21422 23336 21428
rect 22548 21140 22600 21146
rect 22548 21082 22600 21088
rect 21824 20862 22036 20890
rect 21720 20596 21772 20602
rect 21720 20538 21772 20544
rect 21536 20052 21588 20058
rect 21536 19994 21588 20000
rect 21536 19848 21588 19854
rect 21536 19790 21588 19796
rect 21168 19712 21220 19718
rect 21168 19654 21220 19660
rect 21076 19236 21128 19242
rect 21076 19178 21128 19184
rect 20708 18828 20760 18834
rect 20708 18770 20760 18776
rect 20984 18828 21036 18834
rect 20984 18770 21036 18776
rect 20156 18420 20208 18426
rect 20156 18362 20208 18368
rect 19512 18284 19564 18290
rect 19512 18226 19564 18232
rect 18868 18080 18920 18086
rect 18868 18022 18920 18028
rect 19052 18080 19104 18086
rect 19052 18022 19104 18028
rect 18880 17814 18908 18022
rect 18868 17808 18920 17814
rect 18868 17750 18920 17756
rect 19064 17762 19092 18022
rect 19150 17980 19446 18000
rect 19206 17978 19230 17980
rect 19286 17978 19310 17980
rect 19366 17978 19390 17980
rect 19228 17926 19230 17978
rect 19292 17926 19304 17978
rect 19366 17926 19368 17978
rect 19206 17924 19230 17926
rect 19286 17924 19310 17926
rect 19366 17924 19390 17926
rect 19150 17904 19446 17924
rect 19524 17814 19552 18226
rect 20720 18086 20748 18770
rect 20708 18080 20760 18086
rect 20708 18022 20760 18028
rect 19512 17808 19564 17814
rect 19064 17746 19184 17762
rect 19512 17750 19564 17756
rect 18684 17740 18736 17746
rect 19064 17740 19196 17746
rect 19064 17734 19144 17740
rect 18684 17682 18736 17688
rect 19144 17682 19196 17688
rect 18224 17264 18276 17270
rect 18224 17206 18276 17212
rect 17856 17196 17908 17202
rect 17856 17138 17908 17144
rect 17948 17196 18000 17202
rect 17948 17138 18000 17144
rect 17304 16992 17356 16998
rect 17304 16934 17356 16940
rect 17316 16114 17344 16934
rect 17580 16652 17632 16658
rect 17580 16594 17632 16600
rect 17304 16108 17356 16114
rect 17304 16050 17356 16056
rect 17592 15994 17620 16594
rect 17316 15966 17620 15994
rect 17316 15910 17344 15966
rect 17304 15904 17356 15910
rect 17302 15872 17304 15881
rect 17356 15872 17358 15881
rect 17302 15807 17358 15816
rect 17670 15736 17726 15745
rect 17670 15671 17726 15680
rect 17212 15156 17264 15162
rect 17212 15098 17264 15104
rect 17224 14958 17252 15098
rect 17684 15026 17712 15671
rect 17672 15020 17724 15026
rect 17672 14962 17724 14968
rect 17212 14952 17264 14958
rect 17212 14894 17264 14900
rect 17764 14884 17816 14890
rect 17764 14826 17816 14832
rect 17132 14742 17436 14770
rect 16752 14544 16804 14550
rect 16752 14486 16804 14492
rect 15648 14476 15700 14482
rect 15648 14418 15700 14424
rect 15660 13870 15688 14418
rect 15740 14408 15792 14414
rect 15740 14350 15792 14356
rect 15752 14074 15780 14350
rect 15740 14068 15792 14074
rect 15740 14010 15792 14016
rect 15648 13864 15700 13870
rect 15648 13806 15700 13812
rect 15922 13832 15978 13841
rect 15922 13767 15978 13776
rect 15936 13462 15964 13767
rect 15924 13456 15976 13462
rect 15924 13398 15976 13404
rect 15740 13388 15792 13394
rect 15740 13330 15792 13336
rect 15556 12980 15608 12986
rect 15556 12922 15608 12928
rect 15464 12844 15516 12850
rect 15464 12786 15516 12792
rect 15568 12714 15596 12922
rect 15556 12708 15608 12714
rect 15556 12650 15608 12656
rect 15752 12374 15780 13330
rect 16108 12708 16160 12714
rect 16108 12650 16160 12656
rect 15740 12368 15792 12374
rect 15740 12310 15792 12316
rect 15372 12096 15424 12102
rect 15372 12038 15424 12044
rect 15384 11626 15412 12038
rect 15648 11688 15700 11694
rect 15648 11630 15700 11636
rect 15372 11620 15424 11626
rect 15372 11562 15424 11568
rect 15188 11552 15240 11558
rect 15188 11494 15240 11500
rect 15200 11082 15228 11494
rect 15280 11212 15332 11218
rect 15280 11154 15332 11160
rect 15188 11076 15240 11082
rect 15188 11018 15240 11024
rect 15004 10804 15056 10810
rect 15004 10746 15056 10752
rect 14688 10412 14952 10418
rect 14636 10406 14952 10412
rect 14648 10390 14952 10406
rect 14820 10124 14872 10130
rect 14820 10066 14872 10072
rect 14484 9820 14780 9840
rect 14540 9818 14564 9820
rect 14620 9818 14644 9820
rect 14700 9818 14724 9820
rect 14562 9766 14564 9818
rect 14626 9766 14638 9818
rect 14700 9766 14702 9818
rect 14540 9764 14564 9766
rect 14620 9764 14644 9766
rect 14700 9764 14724 9766
rect 14484 9744 14780 9764
rect 14832 9518 14860 10066
rect 14268 9512 14320 9518
rect 14268 9454 14320 9460
rect 14820 9512 14872 9518
rect 14820 9454 14872 9460
rect 14176 9172 14228 9178
rect 14176 9114 14228 9120
rect 14280 8906 14308 9454
rect 14360 9104 14412 9110
rect 14360 9046 14412 9052
rect 14268 8900 14320 8906
rect 14268 8842 14320 8848
rect 14084 7336 14136 7342
rect 14084 7278 14136 7284
rect 13808 7268 13860 7274
rect 13808 7210 13860 7216
rect 13624 7200 13676 7206
rect 13622 7168 13624 7177
rect 13676 7168 13678 7177
rect 13622 7103 13678 7112
rect 14096 6934 14124 7278
rect 14084 6928 14136 6934
rect 14084 6870 14136 6876
rect 12244 6860 12296 6866
rect 12244 6802 12296 6808
rect 13440 6860 13492 6866
rect 13440 6802 13492 6808
rect 13452 6458 13480 6802
rect 13900 6792 13952 6798
rect 13900 6734 13952 6740
rect 12060 6452 12112 6458
rect 12060 6394 12112 6400
rect 13440 6452 13492 6458
rect 13440 6394 13492 6400
rect 11876 6248 11928 6254
rect 11876 6190 11928 6196
rect 11888 5642 11916 6190
rect 13912 5778 13940 6734
rect 13900 5772 13952 5778
rect 13900 5714 13952 5720
rect 11876 5636 11928 5642
rect 11876 5578 11928 5584
rect 13990 5400 14046 5409
rect 13990 5335 13992 5344
rect 14044 5335 14046 5344
rect 13992 5306 14044 5312
rect 14280 4049 14308 8842
rect 14372 8430 14400 9046
rect 14924 9042 14952 10390
rect 14912 9036 14964 9042
rect 14912 8978 14964 8984
rect 14484 8732 14780 8752
rect 14540 8730 14564 8732
rect 14620 8730 14644 8732
rect 14700 8730 14724 8732
rect 14562 8678 14564 8730
rect 14626 8678 14638 8730
rect 14700 8678 14702 8730
rect 14540 8676 14564 8678
rect 14620 8676 14644 8678
rect 14700 8676 14724 8678
rect 14484 8656 14780 8676
rect 14924 8430 14952 8978
rect 14360 8424 14412 8430
rect 14360 8366 14412 8372
rect 14912 8424 14964 8430
rect 14912 8366 14964 8372
rect 14372 8090 14400 8366
rect 14924 8265 14952 8366
rect 14910 8256 14966 8265
rect 14910 8191 14966 8200
rect 14360 8084 14412 8090
rect 14360 8026 14412 8032
rect 14372 7857 14400 8026
rect 15016 8022 15044 10746
rect 15188 10600 15240 10606
rect 15188 10542 15240 10548
rect 15200 10062 15228 10542
rect 15188 10056 15240 10062
rect 15188 9998 15240 10004
rect 15200 9722 15228 9998
rect 15292 9994 15320 11154
rect 15280 9988 15332 9994
rect 15280 9930 15332 9936
rect 15188 9716 15240 9722
rect 15188 9658 15240 9664
rect 15096 9376 15148 9382
rect 15096 9318 15148 9324
rect 15108 8362 15136 9318
rect 15200 9178 15228 9658
rect 15384 9450 15412 11562
rect 15660 11286 15688 11630
rect 15648 11280 15700 11286
rect 15648 11222 15700 11228
rect 15752 10810 15780 12310
rect 16120 11830 16148 12650
rect 17408 12238 17436 14742
rect 17776 14618 17804 14826
rect 17764 14612 17816 14618
rect 17764 14554 17816 14560
rect 17776 13394 17804 14554
rect 17764 13388 17816 13394
rect 17764 13330 17816 13336
rect 17776 12986 17804 13330
rect 17764 12980 17816 12986
rect 17764 12922 17816 12928
rect 17488 12776 17540 12782
rect 17488 12718 17540 12724
rect 17500 12374 17528 12718
rect 17488 12368 17540 12374
rect 17488 12310 17540 12316
rect 17396 12232 17448 12238
rect 17396 12174 17448 12180
rect 16108 11824 16160 11830
rect 16108 11766 16160 11772
rect 16752 11824 16804 11830
rect 16752 11766 16804 11772
rect 16200 11620 16252 11626
rect 16200 11562 16252 11568
rect 16212 11257 16240 11562
rect 16764 11286 16792 11766
rect 17408 11286 17436 12174
rect 17500 11898 17528 12310
rect 17488 11892 17540 11898
rect 17488 11834 17540 11840
rect 17500 11354 17528 11834
rect 17580 11688 17632 11694
rect 17580 11630 17632 11636
rect 17488 11348 17540 11354
rect 17488 11290 17540 11296
rect 16752 11280 16804 11286
rect 16198 11248 16254 11257
rect 16752 11222 16804 11228
rect 17396 11280 17448 11286
rect 17396 11222 17448 11228
rect 16198 11183 16254 11192
rect 16384 11144 16436 11150
rect 16384 11086 16436 11092
rect 16396 10810 16424 11086
rect 16568 11008 16620 11014
rect 16568 10950 16620 10956
rect 15740 10804 15792 10810
rect 15740 10746 15792 10752
rect 16384 10804 16436 10810
rect 16384 10746 16436 10752
rect 15752 10606 15780 10746
rect 16580 10674 16608 10950
rect 16764 10742 16792 11222
rect 17592 11082 17620 11630
rect 17580 11076 17632 11082
rect 17580 11018 17632 11024
rect 16752 10736 16804 10742
rect 16752 10678 16804 10684
rect 16568 10668 16620 10674
rect 16568 10610 16620 10616
rect 15740 10600 15792 10606
rect 15740 10542 15792 10548
rect 16292 10600 16344 10606
rect 16292 10542 16344 10548
rect 15556 9920 15608 9926
rect 15556 9862 15608 9868
rect 15568 9654 15596 9862
rect 15556 9648 15608 9654
rect 15556 9590 15608 9596
rect 15372 9444 15424 9450
rect 15372 9386 15424 9392
rect 15188 9172 15240 9178
rect 15188 9114 15240 9120
rect 15280 8628 15332 8634
rect 15280 8570 15332 8576
rect 15096 8356 15148 8362
rect 15096 8298 15148 8304
rect 15004 8016 15056 8022
rect 15004 7958 15056 7964
rect 14358 7848 14414 7857
rect 14358 7783 14414 7792
rect 14484 7644 14780 7664
rect 14540 7642 14564 7644
rect 14620 7642 14644 7644
rect 14700 7642 14724 7644
rect 14562 7590 14564 7642
rect 14626 7590 14638 7642
rect 14700 7590 14702 7642
rect 14540 7588 14564 7590
rect 14620 7588 14644 7590
rect 14700 7588 14724 7590
rect 14484 7568 14780 7588
rect 15016 7478 15044 7958
rect 15004 7472 15056 7478
rect 15004 7414 15056 7420
rect 14360 7200 14412 7206
rect 14360 7142 14412 7148
rect 14372 6866 14400 7142
rect 14360 6860 14412 6866
rect 14360 6802 14412 6808
rect 15096 6860 15148 6866
rect 15096 6802 15148 6808
rect 15188 6860 15240 6866
rect 15188 6802 15240 6808
rect 14372 6390 14400 6802
rect 14484 6556 14780 6576
rect 14540 6554 14564 6556
rect 14620 6554 14644 6556
rect 14700 6554 14724 6556
rect 14562 6502 14564 6554
rect 14626 6502 14638 6554
rect 14700 6502 14702 6554
rect 14540 6500 14564 6502
rect 14620 6500 14644 6502
rect 14700 6500 14724 6502
rect 14484 6480 14780 6500
rect 15108 6458 15136 6802
rect 15096 6452 15148 6458
rect 15096 6394 15148 6400
rect 15200 6390 15228 6802
rect 14360 6384 14412 6390
rect 14360 6326 14412 6332
rect 15188 6384 15240 6390
rect 15188 6326 15240 6332
rect 15096 6112 15148 6118
rect 15096 6054 15148 6060
rect 15108 5846 15136 6054
rect 15096 5840 15148 5846
rect 15096 5782 15148 5788
rect 15004 5772 15056 5778
rect 15004 5714 15056 5720
rect 14484 5468 14780 5488
rect 14540 5466 14564 5468
rect 14620 5466 14644 5468
rect 14700 5466 14724 5468
rect 14562 5414 14564 5466
rect 14626 5414 14638 5466
rect 14700 5414 14702 5466
rect 14540 5412 14564 5414
rect 14620 5412 14644 5414
rect 14700 5412 14724 5414
rect 14484 5392 14780 5412
rect 14912 5024 14964 5030
rect 14912 4966 14964 4972
rect 14484 4380 14780 4400
rect 14540 4378 14564 4380
rect 14620 4378 14644 4380
rect 14700 4378 14724 4380
rect 14562 4326 14564 4378
rect 14626 4326 14638 4378
rect 14700 4326 14702 4378
rect 14540 4324 14564 4326
rect 14620 4324 14644 4326
rect 14700 4324 14724 4326
rect 14484 4304 14780 4324
rect 14924 4282 14952 4966
rect 15016 4826 15044 5714
rect 15108 5370 15136 5782
rect 15096 5364 15148 5370
rect 15096 5306 15148 5312
rect 15004 4820 15056 4826
rect 15004 4762 15056 4768
rect 14912 4276 14964 4282
rect 14912 4218 14964 4224
rect 14924 4078 14952 4218
rect 14912 4072 14964 4078
rect 14266 4040 14322 4049
rect 14912 4014 14964 4020
rect 14266 3975 14322 3984
rect 14484 3292 14780 3312
rect 14540 3290 14564 3292
rect 14620 3290 14644 3292
rect 14700 3290 14724 3292
rect 14562 3238 14564 3290
rect 14626 3238 14638 3290
rect 14700 3238 14702 3290
rect 14540 3236 14564 3238
rect 14620 3236 14644 3238
rect 14700 3236 14724 3238
rect 14484 3216 14780 3236
rect 14484 2204 14780 2224
rect 14540 2202 14564 2204
rect 14620 2202 14644 2204
rect 14700 2202 14724 2204
rect 14562 2150 14564 2202
rect 14626 2150 14638 2202
rect 14700 2150 14702 2202
rect 14540 2148 14564 2150
rect 14620 2148 14644 2150
rect 14700 2148 14724 2150
rect 14484 2128 14780 2148
rect 15292 480 15320 8570
rect 15384 7750 15412 9386
rect 15464 9036 15516 9042
rect 15464 8978 15516 8984
rect 15476 8634 15504 8978
rect 15752 8634 15780 10542
rect 16304 10266 16332 10542
rect 16292 10260 16344 10266
rect 16292 10202 16344 10208
rect 16304 9994 16332 10202
rect 16292 9988 16344 9994
rect 16292 9930 16344 9936
rect 15832 9920 15884 9926
rect 15832 9862 15884 9868
rect 15844 9654 15872 9862
rect 15832 9648 15884 9654
rect 15832 9590 15884 9596
rect 15924 9376 15976 9382
rect 15924 9318 15976 9324
rect 15936 9042 15964 9318
rect 16764 9110 16792 10678
rect 17868 9602 17896 17138
rect 17960 16726 17988 17138
rect 18040 17060 18092 17066
rect 18040 17002 18092 17008
rect 17948 16720 18000 16726
rect 17948 16662 18000 16668
rect 18052 16658 18080 17002
rect 18236 16658 18264 17206
rect 18696 16998 18724 17682
rect 19156 17338 19184 17682
rect 20156 17536 20208 17542
rect 20154 17504 20156 17513
rect 20208 17504 20210 17513
rect 20154 17439 20210 17448
rect 19144 17332 19196 17338
rect 19144 17274 19196 17280
rect 20720 16998 20748 18022
rect 20996 17746 21024 18770
rect 21088 18426 21116 19178
rect 21180 18902 21208 19654
rect 21548 19122 21576 19790
rect 21628 19168 21680 19174
rect 21548 19116 21628 19122
rect 21548 19110 21680 19116
rect 21548 19094 21668 19110
rect 21168 18896 21220 18902
rect 21168 18838 21220 18844
rect 21352 18624 21404 18630
rect 21352 18566 21404 18572
rect 21076 18420 21128 18426
rect 21076 18362 21128 18368
rect 21364 18222 21392 18566
rect 21352 18216 21404 18222
rect 21352 18158 21404 18164
rect 20800 17740 20852 17746
rect 20800 17682 20852 17688
rect 20984 17740 21036 17746
rect 20984 17682 21036 17688
rect 20812 17134 20840 17682
rect 21364 17202 21392 18158
rect 21548 17814 21576 19094
rect 21628 18420 21680 18426
rect 21628 18362 21680 18368
rect 21640 18154 21668 18362
rect 21628 18148 21680 18154
rect 21628 18090 21680 18096
rect 21640 17814 21668 18090
rect 21536 17808 21588 17814
rect 21536 17750 21588 17756
rect 21628 17808 21680 17814
rect 21628 17750 21680 17756
rect 21536 17604 21588 17610
rect 21536 17546 21588 17552
rect 21444 17536 21496 17542
rect 21444 17478 21496 17484
rect 21352 17196 21404 17202
rect 21352 17138 21404 17144
rect 21456 17134 21484 17478
rect 21548 17338 21576 17546
rect 21536 17332 21588 17338
rect 21536 17274 21588 17280
rect 21640 17134 21668 17750
rect 20800 17128 20852 17134
rect 20800 17070 20852 17076
rect 20892 17128 20944 17134
rect 20892 17070 20944 17076
rect 21444 17128 21496 17134
rect 21444 17070 21496 17076
rect 21628 17128 21680 17134
rect 21628 17070 21680 17076
rect 18684 16992 18736 16998
rect 18684 16934 18736 16940
rect 20708 16992 20760 16998
rect 20708 16934 20760 16940
rect 18696 16794 18724 16934
rect 19150 16892 19446 16912
rect 19206 16890 19230 16892
rect 19286 16890 19310 16892
rect 19366 16890 19390 16892
rect 19228 16838 19230 16890
rect 19292 16838 19304 16890
rect 19366 16838 19368 16890
rect 19206 16836 19230 16838
rect 19286 16836 19310 16838
rect 19366 16836 19390 16838
rect 19150 16816 19446 16836
rect 18684 16788 18736 16794
rect 18684 16730 18736 16736
rect 18776 16720 18828 16726
rect 18776 16662 18828 16668
rect 20154 16688 20210 16697
rect 18040 16652 18092 16658
rect 18040 16594 18092 16600
rect 18224 16652 18276 16658
rect 18224 16594 18276 16600
rect 18788 16232 18816 16662
rect 19052 16652 19104 16658
rect 20720 16658 20748 16934
rect 20154 16623 20210 16632
rect 20708 16652 20760 16658
rect 19052 16594 19104 16600
rect 18868 16244 18920 16250
rect 18788 16204 18868 16232
rect 18868 16186 18920 16192
rect 17948 16040 18000 16046
rect 17948 15982 18000 15988
rect 17960 15706 17988 15982
rect 18592 15972 18644 15978
rect 18592 15914 18644 15920
rect 18222 15736 18278 15745
rect 17948 15700 18000 15706
rect 18222 15671 18224 15680
rect 17948 15642 18000 15648
rect 18276 15671 18278 15680
rect 18224 15642 18276 15648
rect 18604 15638 18632 15914
rect 18592 15632 18644 15638
rect 18592 15574 18644 15580
rect 18604 15162 18632 15574
rect 18776 15496 18828 15502
rect 19064 15484 19092 16594
rect 20168 16114 20196 16623
rect 20708 16594 20760 16600
rect 20156 16108 20208 16114
rect 20156 16050 20208 16056
rect 19150 15804 19446 15824
rect 19206 15802 19230 15804
rect 19286 15802 19310 15804
rect 19366 15802 19390 15804
rect 19228 15750 19230 15802
rect 19292 15750 19304 15802
rect 19366 15750 19368 15802
rect 19206 15748 19230 15750
rect 19286 15748 19310 15750
rect 19366 15748 19390 15750
rect 19150 15728 19446 15748
rect 20168 15638 20196 16050
rect 20720 15978 20748 16594
rect 20708 15972 20760 15978
rect 20708 15914 20760 15920
rect 20156 15632 20208 15638
rect 20156 15574 20208 15580
rect 18828 15456 19092 15484
rect 18776 15438 18828 15444
rect 18960 15360 19012 15366
rect 18960 15302 19012 15308
rect 18592 15156 18644 15162
rect 18592 15098 18644 15104
rect 18972 14890 19000 15302
rect 19064 15162 19092 15456
rect 20524 15496 20576 15502
rect 20524 15438 20576 15444
rect 19052 15156 19104 15162
rect 19052 15098 19104 15104
rect 18960 14884 19012 14890
rect 18960 14826 19012 14832
rect 17948 14544 18000 14550
rect 17948 14486 18000 14492
rect 17960 14074 17988 14486
rect 18132 14408 18184 14414
rect 18132 14350 18184 14356
rect 17948 14068 18000 14074
rect 17948 14010 18000 14016
rect 18144 13870 18172 14350
rect 18132 13864 18184 13870
rect 18130 13832 18132 13841
rect 18184 13832 18186 13841
rect 18130 13767 18186 13776
rect 18776 13456 18828 13462
rect 18776 13398 18828 13404
rect 18684 13252 18736 13258
rect 18684 13194 18736 13200
rect 18316 12708 18368 12714
rect 18316 12650 18368 12656
rect 18328 11286 18356 12650
rect 18500 12232 18552 12238
rect 18500 12174 18552 12180
rect 18512 11762 18540 12174
rect 18696 12084 18724 13194
rect 18788 12986 18816 13398
rect 18972 13326 19000 14826
rect 19052 14816 19104 14822
rect 19052 14758 19104 14764
rect 19064 14498 19092 14758
rect 19150 14716 19446 14736
rect 19206 14714 19230 14716
rect 19286 14714 19310 14716
rect 19366 14714 19390 14716
rect 19228 14662 19230 14714
rect 19292 14662 19304 14714
rect 19366 14662 19368 14714
rect 19206 14660 19230 14662
rect 19286 14660 19310 14662
rect 19366 14660 19390 14662
rect 19150 14640 19446 14660
rect 19064 14470 19184 14498
rect 19156 14278 19184 14470
rect 20536 14414 20564 15438
rect 20708 14884 20760 14890
rect 20708 14826 20760 14832
rect 20720 14793 20748 14826
rect 20706 14784 20762 14793
rect 20706 14719 20762 14728
rect 20616 14544 20668 14550
rect 20616 14486 20668 14492
rect 20524 14408 20576 14414
rect 20524 14350 20576 14356
rect 19144 14272 19196 14278
rect 19144 14214 19196 14220
rect 19156 13870 19184 14214
rect 20536 14074 20564 14350
rect 20524 14068 20576 14074
rect 20524 14010 20576 14016
rect 20628 13938 20656 14486
rect 20720 14414 20748 14719
rect 20708 14408 20760 14414
rect 20708 14350 20760 14356
rect 20616 13932 20668 13938
rect 20616 13874 20668 13880
rect 19144 13864 19196 13870
rect 19144 13806 19196 13812
rect 19150 13628 19446 13648
rect 19206 13626 19230 13628
rect 19286 13626 19310 13628
rect 19366 13626 19390 13628
rect 19228 13574 19230 13626
rect 19292 13574 19304 13626
rect 19366 13574 19368 13626
rect 19206 13572 19230 13574
rect 19286 13572 19310 13574
rect 19366 13572 19390 13574
rect 19150 13552 19446 13572
rect 20812 13394 20840 17070
rect 20904 16658 20932 17070
rect 20892 16652 20944 16658
rect 20892 16594 20944 16600
rect 20904 15910 20932 16594
rect 21444 15972 21496 15978
rect 21444 15914 21496 15920
rect 20892 15904 20944 15910
rect 20892 15846 20944 15852
rect 20800 13388 20852 13394
rect 20800 13330 20852 13336
rect 18960 13320 19012 13326
rect 18960 13262 19012 13268
rect 18776 12980 18828 12986
rect 18776 12922 18828 12928
rect 19512 12844 19564 12850
rect 19512 12786 19564 12792
rect 18960 12640 19012 12646
rect 18960 12582 19012 12588
rect 18776 12096 18828 12102
rect 18696 12064 18776 12084
rect 18828 12064 18830 12073
rect 18696 12056 18774 12064
rect 18774 11999 18830 12008
rect 18500 11756 18552 11762
rect 18500 11698 18552 11704
rect 18316 11280 18368 11286
rect 18316 11222 18368 11228
rect 17948 11144 18000 11150
rect 17948 11086 18000 11092
rect 17960 10470 17988 11086
rect 18328 10810 18356 11222
rect 18512 11150 18540 11698
rect 18592 11552 18644 11558
rect 18592 11494 18644 11500
rect 18500 11144 18552 11150
rect 18500 11086 18552 11092
rect 18604 10810 18632 11494
rect 18972 10810 19000 12582
rect 19150 12540 19446 12560
rect 19206 12538 19230 12540
rect 19286 12538 19310 12540
rect 19366 12538 19390 12540
rect 19228 12486 19230 12538
rect 19292 12486 19304 12538
rect 19366 12486 19368 12538
rect 19206 12484 19230 12486
rect 19286 12484 19310 12486
rect 19366 12484 19390 12486
rect 19150 12464 19446 12484
rect 19524 12374 19552 12786
rect 20524 12776 20576 12782
rect 20524 12718 20576 12724
rect 19972 12708 20024 12714
rect 19972 12650 20024 12656
rect 19512 12368 19564 12374
rect 19512 12310 19564 12316
rect 19984 11830 20012 12650
rect 20536 12646 20564 12718
rect 20812 12646 20840 13330
rect 20904 13297 20932 15846
rect 20984 15360 21036 15366
rect 20984 15302 21036 15308
rect 20996 14958 21024 15302
rect 20984 14952 21036 14958
rect 20984 14894 21036 14900
rect 21456 14482 21484 15914
rect 21640 15178 21668 17070
rect 21824 15502 21852 20862
rect 23296 20806 23324 21422
rect 24308 21298 24336 23423
rect 24400 23322 24428 24126
rect 24480 24132 24532 24138
rect 24480 24074 24532 24080
rect 24584 23866 24612 24210
rect 24572 23860 24624 23866
rect 24572 23802 24624 23808
rect 24480 23520 24532 23526
rect 24480 23462 24532 23468
rect 24388 23316 24440 23322
rect 24388 23258 24440 23264
rect 24492 23089 24520 23462
rect 24572 23180 24624 23186
rect 24572 23122 24624 23128
rect 24478 23080 24534 23089
rect 24478 23015 24534 23024
rect 24584 22642 24612 23122
rect 24572 22636 24624 22642
rect 24572 22578 24624 22584
rect 24478 22264 24534 22273
rect 24478 22199 24534 22208
rect 24492 22098 24520 22199
rect 24480 22092 24532 22098
rect 24480 22034 24532 22040
rect 24388 21888 24440 21894
rect 24388 21830 24440 21836
rect 24400 21593 24428 21830
rect 24492 21690 24520 22034
rect 24480 21684 24532 21690
rect 24480 21626 24532 21632
rect 24386 21584 24442 21593
rect 24386 21519 24442 21528
rect 24216 21270 24336 21298
rect 24480 21344 24532 21350
rect 24480 21286 24532 21292
rect 24216 21146 24244 21270
rect 24294 21176 24350 21185
rect 24204 21140 24256 21146
rect 24294 21111 24350 21120
rect 24204 21082 24256 21088
rect 23008 20800 23060 20806
rect 22928 20748 23008 20754
rect 22928 20742 23060 20748
rect 23284 20800 23336 20806
rect 23284 20742 23336 20748
rect 22928 20726 23048 20742
rect 22928 20058 22956 20726
rect 23817 20700 24113 20720
rect 23873 20698 23897 20700
rect 23953 20698 23977 20700
rect 24033 20698 24057 20700
rect 23895 20646 23897 20698
rect 23959 20646 23971 20698
rect 24033 20646 24035 20698
rect 23873 20644 23897 20646
rect 23953 20644 23977 20646
rect 24033 20644 24057 20646
rect 23817 20624 24113 20644
rect 24308 20534 24336 21111
rect 24492 21049 24520 21286
rect 24478 21040 24534 21049
rect 24388 21004 24440 21010
rect 24478 20975 24534 20984
rect 24388 20946 24440 20952
rect 24400 20602 24428 20946
rect 24388 20596 24440 20602
rect 24388 20538 24440 20544
rect 24296 20528 24348 20534
rect 24296 20470 24348 20476
rect 24480 20392 24532 20398
rect 23006 20360 23062 20369
rect 24480 20334 24532 20340
rect 23006 20295 23062 20304
rect 23020 20262 23048 20295
rect 23008 20256 23060 20262
rect 23008 20198 23060 20204
rect 22916 20052 22968 20058
rect 22916 19994 22968 20000
rect 23652 19916 23704 19922
rect 23652 19858 23704 19864
rect 23560 19712 23612 19718
rect 23560 19654 23612 19660
rect 22272 19304 22324 19310
rect 22272 19246 22324 19252
rect 22284 18426 22312 19246
rect 23572 19242 23600 19654
rect 23664 19378 23692 19858
rect 24386 19816 24442 19825
rect 24386 19751 24388 19760
rect 24440 19751 24442 19760
rect 24388 19722 24440 19728
rect 23817 19612 24113 19632
rect 23873 19610 23897 19612
rect 23953 19610 23977 19612
rect 24033 19610 24057 19612
rect 23895 19558 23897 19610
rect 23959 19558 23971 19610
rect 24033 19558 24035 19610
rect 23873 19556 23897 19558
rect 23953 19556 23977 19558
rect 24033 19556 24057 19558
rect 23817 19536 24113 19556
rect 24492 19378 24520 20334
rect 23652 19372 23704 19378
rect 23652 19314 23704 19320
rect 24204 19372 24256 19378
rect 24204 19314 24256 19320
rect 24480 19372 24532 19378
rect 24480 19314 24532 19320
rect 23376 19236 23428 19242
rect 23376 19178 23428 19184
rect 23560 19236 23612 19242
rect 23560 19178 23612 19184
rect 23388 18970 23416 19178
rect 23376 18964 23428 18970
rect 23376 18906 23428 18912
rect 23664 18902 23692 19314
rect 23742 19136 23798 19145
rect 23742 19071 23798 19080
rect 23652 18896 23704 18902
rect 23652 18838 23704 18844
rect 23560 18760 23612 18766
rect 23560 18702 23612 18708
rect 23572 18426 23600 18702
rect 22272 18420 22324 18426
rect 22272 18362 22324 18368
rect 23560 18420 23612 18426
rect 23560 18362 23612 18368
rect 23664 18306 23692 18838
rect 23572 18278 23692 18306
rect 23572 17882 23600 18278
rect 23652 18080 23704 18086
rect 23652 18022 23704 18028
rect 23560 17876 23612 17882
rect 23560 17818 23612 17824
rect 22364 17672 22416 17678
rect 22364 17614 22416 17620
rect 22376 16998 22404 17614
rect 23664 17338 23692 18022
rect 23652 17332 23704 17338
rect 23652 17274 23704 17280
rect 22364 16992 22416 16998
rect 22364 16934 22416 16940
rect 22376 16726 22404 16934
rect 22364 16720 22416 16726
rect 22364 16662 22416 16668
rect 23190 16688 23246 16697
rect 23756 16658 23784 19071
rect 24216 18902 24244 19314
rect 24296 19168 24348 19174
rect 24296 19110 24348 19116
rect 24204 18896 24256 18902
rect 24204 18838 24256 18844
rect 23817 18524 24113 18544
rect 23873 18522 23897 18524
rect 23953 18522 23977 18524
rect 24033 18522 24057 18524
rect 23895 18470 23897 18522
rect 23959 18470 23971 18522
rect 24033 18470 24035 18522
rect 23873 18468 23897 18470
rect 23953 18468 23977 18470
rect 24033 18468 24057 18470
rect 23817 18448 24113 18468
rect 23928 18148 23980 18154
rect 23928 18090 23980 18096
rect 23940 18057 23968 18090
rect 23926 18048 23982 18057
rect 23926 17983 23982 17992
rect 24204 17808 24256 17814
rect 24204 17750 24256 17756
rect 23817 17436 24113 17456
rect 23873 17434 23897 17436
rect 23953 17434 23977 17436
rect 24033 17434 24057 17436
rect 23895 17382 23897 17434
rect 23959 17382 23971 17434
rect 24033 17382 24035 17434
rect 23873 17380 23897 17382
rect 23953 17380 23977 17382
rect 24033 17380 24057 17382
rect 23817 17360 24113 17380
rect 24216 17134 24244 17750
rect 24308 17678 24336 19110
rect 24388 18284 24440 18290
rect 24388 18226 24440 18232
rect 24296 17672 24348 17678
rect 24296 17614 24348 17620
rect 24204 17128 24256 17134
rect 24204 17070 24256 17076
rect 24308 16794 24336 17614
rect 24400 17610 24428 18226
rect 24478 18048 24534 18057
rect 24478 17983 24534 17992
rect 24388 17604 24440 17610
rect 24388 17546 24440 17552
rect 24492 17338 24520 17983
rect 24480 17332 24532 17338
rect 24480 17274 24532 17280
rect 24938 17096 24994 17105
rect 24938 17031 24994 17040
rect 24296 16788 24348 16794
rect 24296 16730 24348 16736
rect 24388 16720 24440 16726
rect 24388 16662 24440 16668
rect 23190 16623 23192 16632
rect 23244 16623 23246 16632
rect 23744 16652 23796 16658
rect 23192 16594 23244 16600
rect 23744 16594 23796 16600
rect 24296 16652 24348 16658
rect 24296 16594 24348 16600
rect 23008 16448 23060 16454
rect 23008 16390 23060 16396
rect 23020 16153 23048 16390
rect 23817 16348 24113 16368
rect 23873 16346 23897 16348
rect 23953 16346 23977 16348
rect 24033 16346 24057 16348
rect 23895 16294 23897 16346
rect 23959 16294 23971 16346
rect 24033 16294 24035 16346
rect 23873 16292 23897 16294
rect 23953 16292 23977 16294
rect 24033 16292 24057 16294
rect 23817 16272 24113 16292
rect 24308 16250 24336 16594
rect 24296 16244 24348 16250
rect 24296 16186 24348 16192
rect 23006 16144 23062 16153
rect 23006 16079 23062 16088
rect 24400 16046 24428 16662
rect 24952 16250 24980 17031
rect 24940 16244 24992 16250
rect 24940 16186 24992 16192
rect 25044 16114 25072 24550
rect 25306 24304 25362 24313
rect 25306 24239 25362 24248
rect 25320 23866 25348 24239
rect 25308 23860 25360 23866
rect 25308 23802 25360 23808
rect 25320 23662 25348 23802
rect 25308 23656 25360 23662
rect 25308 23598 25360 23604
rect 25872 23497 25900 27520
rect 25858 23488 25914 23497
rect 25858 23423 25914 23432
rect 25306 23216 25362 23225
rect 25306 23151 25362 23160
rect 25320 21690 25348 23151
rect 25308 21684 25360 21690
rect 25308 21626 25360 21632
rect 25320 21486 25348 21626
rect 25308 21480 25360 21486
rect 25308 21422 25360 21428
rect 25398 20088 25454 20097
rect 25398 20023 25454 20032
rect 25412 19922 25440 20023
rect 25400 19916 25452 19922
rect 25400 19858 25452 19864
rect 25412 19514 25440 19858
rect 25400 19508 25452 19514
rect 25400 19450 25452 19456
rect 26884 19310 26912 27520
rect 26872 19304 26924 19310
rect 26872 19246 26924 19252
rect 25490 18048 25546 18057
rect 25490 17983 25546 17992
rect 25504 17338 25532 17983
rect 25492 17332 25544 17338
rect 25492 17274 25544 17280
rect 25504 17134 25532 17274
rect 25492 17128 25544 17134
rect 25492 17070 25544 17076
rect 25032 16108 25084 16114
rect 25032 16050 25084 16056
rect 24388 16040 24440 16046
rect 24202 16008 24258 16017
rect 23376 15972 23428 15978
rect 23376 15914 23428 15920
rect 23928 15972 23980 15978
rect 24388 15982 24440 15988
rect 24202 15943 24258 15952
rect 23928 15914 23980 15920
rect 23388 15706 23416 15914
rect 23376 15700 23428 15706
rect 23376 15642 23428 15648
rect 23940 15638 23968 15914
rect 21904 15632 21956 15638
rect 21904 15574 21956 15580
rect 23192 15632 23244 15638
rect 23192 15574 23244 15580
rect 23928 15632 23980 15638
rect 23928 15574 23980 15580
rect 21812 15496 21864 15502
rect 21812 15438 21864 15444
rect 21548 15150 21668 15178
rect 21548 14890 21576 15150
rect 21824 15094 21852 15438
rect 21916 15162 21944 15574
rect 21904 15156 21956 15162
rect 21904 15098 21956 15104
rect 21812 15088 21864 15094
rect 21812 15030 21864 15036
rect 22088 14952 22140 14958
rect 22088 14894 22140 14900
rect 21536 14884 21588 14890
rect 21536 14826 21588 14832
rect 21444 14476 21496 14482
rect 21444 14418 21496 14424
rect 21352 14272 21404 14278
rect 21352 14214 21404 14220
rect 21364 13870 21392 14214
rect 21352 13864 21404 13870
rect 21352 13806 21404 13812
rect 21364 13462 21392 13806
rect 21352 13456 21404 13462
rect 21074 13424 21130 13433
rect 21352 13398 21404 13404
rect 21074 13359 21076 13368
rect 21128 13359 21130 13368
rect 21076 13330 21128 13336
rect 20890 13288 20946 13297
rect 20890 13223 20946 13232
rect 21456 12918 21484 14418
rect 21548 13802 21576 14826
rect 22100 14618 22128 14894
rect 23204 14618 23232 15574
rect 23376 15564 23428 15570
rect 23376 15506 23428 15512
rect 23388 15162 23416 15506
rect 23817 15260 24113 15280
rect 23873 15258 23897 15260
rect 23953 15258 23977 15260
rect 24033 15258 24057 15260
rect 23895 15206 23897 15258
rect 23959 15206 23971 15258
rect 24033 15206 24035 15258
rect 23873 15204 23897 15206
rect 23953 15204 23977 15206
rect 24033 15204 24057 15206
rect 23817 15184 24113 15204
rect 23376 15156 23428 15162
rect 23376 15098 23428 15104
rect 24216 14822 24244 15943
rect 24848 15564 24900 15570
rect 24848 15506 24900 15512
rect 24296 15360 24348 15366
rect 24296 15302 24348 15308
rect 24308 15162 24336 15302
rect 24296 15156 24348 15162
rect 24296 15098 24348 15104
rect 24860 14822 24888 15506
rect 24938 14920 24994 14929
rect 24938 14855 24994 14864
rect 24204 14816 24256 14822
rect 24848 14816 24900 14822
rect 24204 14758 24256 14764
rect 24846 14784 24848 14793
rect 24900 14784 24902 14793
rect 24846 14719 24902 14728
rect 22088 14612 22140 14618
rect 22088 14554 22140 14560
rect 23192 14612 23244 14618
rect 23192 14554 23244 14560
rect 22364 14476 22416 14482
rect 22364 14418 22416 14424
rect 21812 14408 21864 14414
rect 21812 14350 21864 14356
rect 21536 13796 21588 13802
rect 21536 13738 21588 13744
rect 21444 12912 21496 12918
rect 21444 12854 21496 12860
rect 21352 12844 21404 12850
rect 21352 12786 21404 12792
rect 21168 12776 21220 12782
rect 21168 12718 21220 12724
rect 20524 12640 20576 12646
rect 20524 12582 20576 12588
rect 20800 12640 20852 12646
rect 20800 12582 20852 12588
rect 19972 11824 20024 11830
rect 19972 11766 20024 11772
rect 19150 11452 19446 11472
rect 19206 11450 19230 11452
rect 19286 11450 19310 11452
rect 19366 11450 19390 11452
rect 19228 11398 19230 11450
rect 19292 11398 19304 11450
rect 19366 11398 19368 11450
rect 19206 11396 19230 11398
rect 19286 11396 19310 11398
rect 19366 11396 19390 11398
rect 19150 11376 19446 11396
rect 18316 10804 18368 10810
rect 18316 10746 18368 10752
rect 18592 10804 18644 10810
rect 18592 10746 18644 10752
rect 18960 10804 19012 10810
rect 18960 10746 19012 10752
rect 18604 10606 18632 10746
rect 19694 10704 19750 10713
rect 19694 10639 19696 10648
rect 19748 10639 19750 10648
rect 19696 10610 19748 10616
rect 18592 10600 18644 10606
rect 18592 10542 18644 10548
rect 17948 10464 18000 10470
rect 17948 10406 18000 10412
rect 17960 9761 17988 10406
rect 19150 10364 19446 10384
rect 19206 10362 19230 10364
rect 19286 10362 19310 10364
rect 19366 10362 19390 10364
rect 19228 10310 19230 10362
rect 19292 10310 19304 10362
rect 19366 10310 19368 10362
rect 19206 10308 19230 10310
rect 19286 10308 19310 10310
rect 19366 10308 19390 10310
rect 19150 10288 19446 10308
rect 20536 10130 20564 12582
rect 20812 12306 20840 12582
rect 21180 12306 21208 12718
rect 20800 12300 20852 12306
rect 20800 12242 20852 12248
rect 21168 12300 21220 12306
rect 21168 12242 21220 12248
rect 20616 12232 20668 12238
rect 20616 12174 20668 12180
rect 20628 11286 20656 12174
rect 20812 11898 20840 12242
rect 21260 12232 21312 12238
rect 21260 12174 21312 12180
rect 20800 11892 20852 11898
rect 20800 11834 20852 11840
rect 20616 11280 20668 11286
rect 20614 11248 20616 11257
rect 20668 11248 20670 11257
rect 20614 11183 20670 11192
rect 20812 10674 20840 11834
rect 21272 11218 21300 12174
rect 21364 11762 21392 12786
rect 21548 11898 21576 13738
rect 21824 13394 21852 14350
rect 22376 14006 22404 14418
rect 23204 14006 23232 14554
rect 24204 14476 24256 14482
rect 24204 14418 24256 14424
rect 23560 14408 23612 14414
rect 23560 14350 23612 14356
rect 23376 14068 23428 14074
rect 23376 14010 23428 14016
rect 22364 14000 22416 14006
rect 22364 13942 22416 13948
rect 23192 14000 23244 14006
rect 23192 13942 23244 13948
rect 23388 13802 23416 14010
rect 23376 13796 23428 13802
rect 23376 13738 23428 13744
rect 23468 13728 23520 13734
rect 23468 13670 23520 13676
rect 21812 13388 21864 13394
rect 21812 13330 21864 13336
rect 22180 13388 22232 13394
rect 22180 13330 22232 13336
rect 21824 12986 21852 13330
rect 21812 12980 21864 12986
rect 21812 12922 21864 12928
rect 22192 12714 22220 13330
rect 23480 13326 23508 13670
rect 23572 13462 23600 14350
rect 23817 14172 24113 14192
rect 23873 14170 23897 14172
rect 23953 14170 23977 14172
rect 24033 14170 24057 14172
rect 23895 14118 23897 14170
rect 23959 14118 23971 14170
rect 24033 14118 24035 14170
rect 23873 14116 23897 14118
rect 23953 14116 23977 14118
rect 24033 14116 24057 14118
rect 23817 14096 24113 14116
rect 24216 14074 24244 14418
rect 24204 14068 24256 14074
rect 24204 14010 24256 14016
rect 23928 13796 23980 13802
rect 23928 13738 23980 13744
rect 23940 13462 23968 13738
rect 24952 13530 24980 14855
rect 24940 13524 24992 13530
rect 24940 13466 24992 13472
rect 23560 13456 23612 13462
rect 23560 13398 23612 13404
rect 23928 13456 23980 13462
rect 23928 13398 23980 13404
rect 24204 13456 24256 13462
rect 24204 13398 24256 13404
rect 23468 13320 23520 13326
rect 23468 13262 23520 13268
rect 23480 12850 23508 13262
rect 23572 12986 23600 13398
rect 23817 13084 24113 13104
rect 23873 13082 23897 13084
rect 23953 13082 23977 13084
rect 24033 13082 24057 13084
rect 23895 13030 23897 13082
rect 23959 13030 23971 13082
rect 24033 13030 24035 13082
rect 23873 13028 23897 13030
rect 23953 13028 23977 13030
rect 24033 13028 24057 13030
rect 23817 13008 24113 13028
rect 24216 12986 24244 13398
rect 24756 13388 24808 13394
rect 24756 13330 24808 13336
rect 24768 12986 24796 13330
rect 23560 12980 23612 12986
rect 23560 12922 23612 12928
rect 24204 12980 24256 12986
rect 24204 12922 24256 12928
rect 24756 12980 24808 12986
rect 24756 12922 24808 12928
rect 23468 12844 23520 12850
rect 23468 12786 23520 12792
rect 24216 12782 24244 12922
rect 24846 12880 24902 12889
rect 24846 12815 24902 12824
rect 24204 12776 24256 12782
rect 24204 12718 24256 12724
rect 22180 12708 22232 12714
rect 22180 12650 22232 12656
rect 23376 12640 23428 12646
rect 23376 12582 23428 12588
rect 22916 12300 22968 12306
rect 22916 12242 22968 12248
rect 22928 11898 22956 12242
rect 23190 12064 23246 12073
rect 23190 11999 23246 12008
rect 21536 11892 21588 11898
rect 21536 11834 21588 11840
rect 22916 11892 22968 11898
rect 22916 11834 22968 11840
rect 21352 11756 21404 11762
rect 21352 11698 21404 11704
rect 21364 11354 21392 11698
rect 21548 11626 21576 11834
rect 21536 11620 21588 11626
rect 21536 11562 21588 11568
rect 21352 11348 21404 11354
rect 21352 11290 21404 11296
rect 21548 11286 21576 11562
rect 22928 11558 22956 11834
rect 22916 11552 22968 11558
rect 22916 11494 22968 11500
rect 21536 11280 21588 11286
rect 21536 11222 21588 11228
rect 21812 11280 21864 11286
rect 21812 11222 21864 11228
rect 21260 11212 21312 11218
rect 21260 11154 21312 11160
rect 20800 10668 20852 10674
rect 20800 10610 20852 10616
rect 20892 10532 20944 10538
rect 20892 10474 20944 10480
rect 21536 10532 21588 10538
rect 21536 10474 21588 10480
rect 20708 10260 20760 10266
rect 20708 10202 20760 10208
rect 18868 10124 18920 10130
rect 18868 10066 18920 10072
rect 20524 10124 20576 10130
rect 20524 10066 20576 10072
rect 17946 9752 18002 9761
rect 17946 9687 18002 9696
rect 18880 9654 18908 10066
rect 18960 9920 19012 9926
rect 18960 9862 19012 9868
rect 18868 9648 18920 9654
rect 17868 9574 17988 9602
rect 18868 9590 18920 9596
rect 16752 9104 16804 9110
rect 16752 9046 16804 9052
rect 17672 9104 17724 9110
rect 17672 9046 17724 9052
rect 15924 9036 15976 9042
rect 15924 8978 15976 8984
rect 16384 9036 16436 9042
rect 16384 8978 16436 8984
rect 16396 8838 16424 8978
rect 16568 8968 16620 8974
rect 16568 8910 16620 8916
rect 16384 8832 16436 8838
rect 16384 8774 16436 8780
rect 15464 8628 15516 8634
rect 15464 8570 15516 8576
rect 15740 8628 15792 8634
rect 15740 8570 15792 8576
rect 15752 8430 15780 8570
rect 16396 8430 16424 8774
rect 15740 8424 15792 8430
rect 15740 8366 15792 8372
rect 16200 8424 16252 8430
rect 16200 8366 16252 8372
rect 16384 8424 16436 8430
rect 16384 8366 16436 8372
rect 16106 8256 16162 8265
rect 16106 8191 16162 8200
rect 16120 7954 16148 8191
rect 16108 7948 16160 7954
rect 16108 7890 16160 7896
rect 15372 7744 15424 7750
rect 15372 7686 15424 7692
rect 15556 7744 15608 7750
rect 15556 7686 15608 7692
rect 15384 7274 15412 7686
rect 15568 7478 15596 7686
rect 16120 7546 16148 7890
rect 16108 7540 16160 7546
rect 16108 7482 16160 7488
rect 15556 7472 15608 7478
rect 15556 7414 15608 7420
rect 15568 7342 15596 7414
rect 15556 7336 15608 7342
rect 15556 7278 15608 7284
rect 15372 7268 15424 7274
rect 15372 7210 15424 7216
rect 15384 7002 15412 7210
rect 15372 6996 15424 7002
rect 15372 6938 15424 6944
rect 16212 6866 16240 8366
rect 16580 8090 16608 8910
rect 16764 8634 16792 9046
rect 17684 8838 17712 9046
rect 17672 8832 17724 8838
rect 17672 8774 17724 8780
rect 16752 8628 16804 8634
rect 16752 8570 16804 8576
rect 17580 8424 17632 8430
rect 17580 8366 17632 8372
rect 17592 8090 17620 8366
rect 17684 8294 17712 8774
rect 17764 8356 17816 8362
rect 17764 8298 17816 8304
rect 17672 8288 17724 8294
rect 17672 8230 17724 8236
rect 16568 8084 16620 8090
rect 16568 8026 16620 8032
rect 17580 8084 17632 8090
rect 17580 8026 17632 8032
rect 16476 7948 16528 7954
rect 16476 7890 16528 7896
rect 16488 7206 16516 7890
rect 17488 7880 17540 7886
rect 17488 7822 17540 7828
rect 16476 7200 16528 7206
rect 16476 7142 16528 7148
rect 16936 7200 16988 7206
rect 16936 7142 16988 7148
rect 16948 6866 16976 7142
rect 17118 7032 17174 7041
rect 17118 6967 17174 6976
rect 17132 6934 17160 6967
rect 17120 6928 17172 6934
rect 17120 6870 17172 6876
rect 16200 6860 16252 6866
rect 16200 6802 16252 6808
rect 16568 6860 16620 6866
rect 16568 6802 16620 6808
rect 16936 6860 16988 6866
rect 16936 6802 16988 6808
rect 15372 6792 15424 6798
rect 15372 6734 15424 6740
rect 15384 6322 15412 6734
rect 16580 6458 16608 6802
rect 16948 6458 16976 6802
rect 16568 6452 16620 6458
rect 16568 6394 16620 6400
rect 16936 6452 16988 6458
rect 16936 6394 16988 6400
rect 17500 6322 17528 7822
rect 17684 7342 17712 8230
rect 17672 7336 17724 7342
rect 17672 7278 17724 7284
rect 15372 6316 15424 6322
rect 15372 6258 15424 6264
rect 17488 6316 17540 6322
rect 17488 6258 17540 6264
rect 16292 6112 16344 6118
rect 16292 6054 16344 6060
rect 16304 5846 16332 6054
rect 17500 5914 17528 6258
rect 17776 6186 17804 8298
rect 17960 6361 17988 9574
rect 18776 9444 18828 9450
rect 18776 9386 18828 9392
rect 18406 9072 18462 9081
rect 18406 9007 18462 9016
rect 18420 8974 18448 9007
rect 18788 8974 18816 9386
rect 18880 9382 18908 9590
rect 18868 9376 18920 9382
rect 18868 9318 18920 9324
rect 18408 8968 18460 8974
rect 18408 8910 18460 8916
rect 18776 8968 18828 8974
rect 18776 8910 18828 8916
rect 18420 8090 18448 8910
rect 18788 8514 18816 8910
rect 18880 8634 18908 9318
rect 18972 8634 19000 9862
rect 20536 9586 20564 10066
rect 20524 9580 20576 9586
rect 20524 9522 20576 9528
rect 19694 9480 19750 9489
rect 19694 9415 19696 9424
rect 19748 9415 19750 9424
rect 19696 9386 19748 9392
rect 19150 9276 19446 9296
rect 19206 9274 19230 9276
rect 19286 9274 19310 9276
rect 19366 9274 19390 9276
rect 19228 9222 19230 9274
rect 19292 9222 19304 9274
rect 19366 9222 19368 9274
rect 19206 9220 19230 9222
rect 19286 9220 19310 9222
rect 19366 9220 19390 9222
rect 19150 9200 19446 9220
rect 19512 9172 19564 9178
rect 19512 9114 19564 9120
rect 18868 8628 18920 8634
rect 18868 8570 18920 8576
rect 18960 8628 19012 8634
rect 18960 8570 19012 8576
rect 18788 8486 18908 8514
rect 19524 8498 19552 9114
rect 19708 8498 19736 9386
rect 20432 9376 20484 9382
rect 20432 9318 20484 9324
rect 20444 9178 20472 9318
rect 20432 9172 20484 9178
rect 20432 9114 20484 9120
rect 20720 9042 20748 10202
rect 20904 10130 20932 10474
rect 20892 10124 20944 10130
rect 20892 10066 20944 10072
rect 20904 9722 20932 10066
rect 20892 9716 20944 9722
rect 20892 9658 20944 9664
rect 21548 9178 21576 10474
rect 21824 10470 21852 11222
rect 22548 11212 22600 11218
rect 22548 11154 22600 11160
rect 22560 10810 22588 11154
rect 23008 11008 23060 11014
rect 23008 10950 23060 10956
rect 22548 10804 22600 10810
rect 22548 10746 22600 10752
rect 22914 10568 22970 10577
rect 22914 10503 22970 10512
rect 21812 10464 21864 10470
rect 21812 10406 21864 10412
rect 22088 10464 22140 10470
rect 22088 10406 22140 10412
rect 21536 9172 21588 9178
rect 21536 9114 21588 9120
rect 21260 9104 21312 9110
rect 21260 9046 21312 9052
rect 20708 9036 20760 9042
rect 20708 8978 20760 8984
rect 20720 8634 20748 8978
rect 21272 8634 21300 9046
rect 20708 8628 20760 8634
rect 20708 8570 20760 8576
rect 21260 8628 21312 8634
rect 21260 8570 21312 8576
rect 18408 8084 18460 8090
rect 18408 8026 18460 8032
rect 18592 8016 18644 8022
rect 18592 7958 18644 7964
rect 18500 7880 18552 7886
rect 18500 7822 18552 7828
rect 18512 7206 18540 7822
rect 18604 7410 18632 7958
rect 18880 7886 18908 8486
rect 19512 8492 19564 8498
rect 19512 8434 19564 8440
rect 19696 8492 19748 8498
rect 19696 8434 19748 8440
rect 21272 8362 21300 8570
rect 21548 8498 21576 9114
rect 21824 9110 21852 10406
rect 22100 9722 22128 10406
rect 22928 10266 22956 10503
rect 23020 10470 23048 10950
rect 23008 10464 23060 10470
rect 23008 10406 23060 10412
rect 22916 10260 22968 10266
rect 22916 10202 22968 10208
rect 22640 10124 22692 10130
rect 22640 10066 22692 10072
rect 22652 9994 22680 10066
rect 22916 10056 22968 10062
rect 22916 9998 22968 10004
rect 22640 9988 22692 9994
rect 22640 9930 22692 9936
rect 22088 9716 22140 9722
rect 22088 9658 22140 9664
rect 22088 9512 22140 9518
rect 22086 9480 22088 9489
rect 22140 9480 22142 9489
rect 22086 9415 22142 9424
rect 22652 9178 22680 9930
rect 22928 9722 22956 9998
rect 22916 9716 22968 9722
rect 22916 9658 22968 9664
rect 22640 9172 22692 9178
rect 22640 9114 22692 9120
rect 21812 9104 21864 9110
rect 21812 9046 21864 9052
rect 23100 9104 23152 9110
rect 23100 9046 23152 9052
rect 23008 8968 23060 8974
rect 23008 8910 23060 8916
rect 21628 8832 21680 8838
rect 21628 8774 21680 8780
rect 21536 8492 21588 8498
rect 21536 8434 21588 8440
rect 21260 8356 21312 8362
rect 21260 8298 21312 8304
rect 19150 8188 19446 8208
rect 19206 8186 19230 8188
rect 19286 8186 19310 8188
rect 19366 8186 19390 8188
rect 19228 8134 19230 8186
rect 19292 8134 19304 8186
rect 19366 8134 19368 8186
rect 19206 8132 19230 8134
rect 19286 8132 19310 8134
rect 19366 8132 19390 8134
rect 19150 8112 19446 8132
rect 21640 8022 21668 8774
rect 23020 8634 23048 8910
rect 22824 8628 22876 8634
rect 22824 8570 22876 8576
rect 23008 8628 23060 8634
rect 23008 8570 23060 8576
rect 21628 8016 21680 8022
rect 20982 7984 21038 7993
rect 21628 7958 21680 7964
rect 20982 7919 21038 7928
rect 20996 7886 21024 7919
rect 18868 7880 18920 7886
rect 18868 7822 18920 7828
rect 20984 7880 21036 7886
rect 20984 7822 21036 7828
rect 20996 7546 21024 7822
rect 21640 7546 21668 7958
rect 22270 7848 22326 7857
rect 22270 7783 22326 7792
rect 20984 7540 21036 7546
rect 20984 7482 21036 7488
rect 21628 7540 21680 7546
rect 21628 7482 21680 7488
rect 18592 7404 18644 7410
rect 18592 7346 18644 7352
rect 21640 7342 21668 7482
rect 21628 7336 21680 7342
rect 21628 7278 21680 7284
rect 18500 7200 18552 7206
rect 19604 7200 19656 7206
rect 18500 7142 18552 7148
rect 19602 7168 19604 7177
rect 20248 7200 20300 7206
rect 19656 7168 19658 7177
rect 19150 7100 19446 7120
rect 20248 7142 20300 7148
rect 19602 7103 19658 7112
rect 19206 7098 19230 7100
rect 19286 7098 19310 7100
rect 19366 7098 19390 7100
rect 19228 7046 19230 7098
rect 19292 7046 19304 7098
rect 19366 7046 19368 7098
rect 19206 7044 19230 7046
rect 19286 7044 19310 7046
rect 19366 7044 19390 7046
rect 18958 7032 19014 7041
rect 19150 7024 19446 7044
rect 19014 6990 19092 7018
rect 18958 6967 19014 6976
rect 18868 6928 18920 6934
rect 18498 6896 18554 6905
rect 18868 6870 18920 6876
rect 18498 6831 18500 6840
rect 18552 6831 18554 6840
rect 18500 6802 18552 6808
rect 18880 6458 18908 6870
rect 18868 6452 18920 6458
rect 18868 6394 18920 6400
rect 17946 6352 18002 6361
rect 17946 6287 18002 6296
rect 17764 6180 17816 6186
rect 17764 6122 17816 6128
rect 17488 5908 17540 5914
rect 17488 5850 17540 5856
rect 16292 5840 16344 5846
rect 16292 5782 16344 5788
rect 16936 5840 16988 5846
rect 16936 5782 16988 5788
rect 16660 5704 16712 5710
rect 16660 5646 16712 5652
rect 15740 5568 15792 5574
rect 15740 5510 15792 5516
rect 15752 5098 15780 5510
rect 16672 5370 16700 5646
rect 16948 5370 16976 5782
rect 18592 5772 18644 5778
rect 18592 5714 18644 5720
rect 17396 5704 17448 5710
rect 17396 5646 17448 5652
rect 18132 5704 18184 5710
rect 18132 5646 18184 5652
rect 17408 5545 17436 5646
rect 17394 5536 17450 5545
rect 17394 5471 17450 5480
rect 16660 5364 16712 5370
rect 16660 5306 16712 5312
rect 16936 5364 16988 5370
rect 16936 5306 16988 5312
rect 15740 5092 15792 5098
rect 15740 5034 15792 5040
rect 16672 4758 16700 5306
rect 17408 5250 17436 5471
rect 17408 5234 17528 5250
rect 17408 5228 17540 5234
rect 17408 5222 17488 5228
rect 17488 5170 17540 5176
rect 18144 5098 18172 5646
rect 18604 5370 18632 5714
rect 18592 5364 18644 5370
rect 18592 5306 18644 5312
rect 17672 5092 17724 5098
rect 17672 5034 17724 5040
rect 18132 5092 18184 5098
rect 18132 5034 18184 5040
rect 17684 4826 17712 5034
rect 17672 4820 17724 4826
rect 17672 4762 17724 4768
rect 15924 4752 15976 4758
rect 15924 4694 15976 4700
rect 16660 4752 16712 4758
rect 16660 4694 16712 4700
rect 15936 4146 15964 4694
rect 18880 4690 18908 6394
rect 19064 6322 19092 6990
rect 19880 6792 19932 6798
rect 19880 6734 19932 6740
rect 19052 6316 19104 6322
rect 19052 6258 19104 6264
rect 19064 5914 19092 6258
rect 19696 6180 19748 6186
rect 19696 6122 19748 6128
rect 19708 6089 19736 6122
rect 19694 6080 19750 6089
rect 19150 6012 19446 6032
rect 19694 6015 19750 6024
rect 19206 6010 19230 6012
rect 19286 6010 19310 6012
rect 19366 6010 19390 6012
rect 19228 5958 19230 6010
rect 19292 5958 19304 6010
rect 19366 5958 19368 6010
rect 19206 5956 19230 5958
rect 19286 5956 19310 5958
rect 19366 5956 19390 5958
rect 19150 5936 19446 5956
rect 19052 5908 19104 5914
rect 19052 5850 19104 5856
rect 19892 5710 19920 6734
rect 20260 6458 20288 7142
rect 21640 7002 21668 7278
rect 21628 6996 21680 7002
rect 21628 6938 21680 6944
rect 21076 6860 21128 6866
rect 21076 6802 21128 6808
rect 20892 6656 20944 6662
rect 20892 6598 20944 6604
rect 20904 6458 20932 6598
rect 21088 6458 21116 6802
rect 20248 6452 20300 6458
rect 20248 6394 20300 6400
rect 20892 6452 20944 6458
rect 20892 6394 20944 6400
rect 21076 6452 21128 6458
rect 21076 6394 21128 6400
rect 20800 6384 20852 6390
rect 20852 6332 21024 6338
rect 20800 6326 21024 6332
rect 20812 6322 21024 6326
rect 20812 6316 21036 6322
rect 20812 6310 20984 6316
rect 20984 6258 21036 6264
rect 20248 6112 20300 6118
rect 20248 6054 20300 6060
rect 20260 5914 20288 6054
rect 21088 5914 21116 6394
rect 21444 6316 21496 6322
rect 21444 6258 21496 6264
rect 20248 5908 20300 5914
rect 20248 5850 20300 5856
rect 21076 5908 21128 5914
rect 21076 5850 21128 5856
rect 19880 5704 19932 5710
rect 19880 5646 19932 5652
rect 19892 5234 19920 5646
rect 20260 5370 20288 5850
rect 21456 5846 21484 6258
rect 21444 5840 21496 5846
rect 21444 5782 21496 5788
rect 20248 5364 20300 5370
rect 20248 5306 20300 5312
rect 19880 5228 19932 5234
rect 19880 5170 19932 5176
rect 19604 5092 19656 5098
rect 19604 5034 19656 5040
rect 19512 5024 19564 5030
rect 19512 4966 19564 4972
rect 19150 4924 19446 4944
rect 19206 4922 19230 4924
rect 19286 4922 19310 4924
rect 19366 4922 19390 4924
rect 19228 4870 19230 4922
rect 19292 4870 19304 4922
rect 19366 4870 19368 4922
rect 19206 4868 19230 4870
rect 19286 4868 19310 4870
rect 19366 4868 19390 4870
rect 19150 4848 19446 4868
rect 19524 4758 19552 4966
rect 19512 4752 19564 4758
rect 19512 4694 19564 4700
rect 18868 4684 18920 4690
rect 18868 4626 18920 4632
rect 16200 4616 16252 4622
rect 16200 4558 16252 4564
rect 16212 4146 16240 4558
rect 18880 4282 18908 4626
rect 18868 4276 18920 4282
rect 18868 4218 18920 4224
rect 15924 4140 15976 4146
rect 15924 4082 15976 4088
rect 16200 4140 16252 4146
rect 16200 4082 16252 4088
rect 16212 3738 16240 4082
rect 19616 4049 19644 5034
rect 18774 4040 18830 4049
rect 18774 3975 18830 3984
rect 19602 4040 19658 4049
rect 19602 3975 19658 3984
rect 16200 3732 16252 3738
rect 16200 3674 16252 3680
rect 16292 3596 16344 3602
rect 16292 3538 16344 3544
rect 16304 2990 16332 3538
rect 16292 2984 16344 2990
rect 16290 2952 16292 2961
rect 16344 2952 16346 2961
rect 16290 2887 16346 2896
rect 18788 480 18816 3975
rect 19150 3836 19446 3856
rect 19206 3834 19230 3836
rect 19286 3834 19310 3836
rect 19366 3834 19390 3836
rect 19228 3782 19230 3834
rect 19292 3782 19304 3834
rect 19366 3782 19368 3834
rect 19206 3780 19230 3782
rect 19286 3780 19310 3782
rect 19366 3780 19390 3782
rect 19150 3760 19446 3780
rect 19150 2748 19446 2768
rect 19206 2746 19230 2748
rect 19286 2746 19310 2748
rect 19366 2746 19390 2748
rect 19228 2694 19230 2746
rect 19292 2694 19304 2746
rect 19366 2694 19368 2746
rect 19206 2692 19230 2694
rect 19286 2692 19310 2694
rect 19366 2692 19390 2694
rect 19150 2672 19446 2692
rect 22284 480 22312 7783
rect 22836 6866 22864 8570
rect 23112 8294 23140 9046
rect 23100 8288 23152 8294
rect 23020 8236 23100 8242
rect 23020 8230 23152 8236
rect 23020 8214 23140 8230
rect 23020 7410 23048 8214
rect 23204 8129 23232 11999
rect 23282 11656 23338 11665
rect 23282 11591 23284 11600
rect 23336 11591 23338 11600
rect 23284 11562 23336 11568
rect 23296 11354 23324 11562
rect 23284 11348 23336 11354
rect 23284 11290 23336 11296
rect 23284 10464 23336 10470
rect 23284 10406 23336 10412
rect 23296 9926 23324 10406
rect 23284 9920 23336 9926
rect 23284 9862 23336 9868
rect 23296 9518 23324 9862
rect 23284 9512 23336 9518
rect 23284 9454 23336 9460
rect 23284 8832 23336 8838
rect 23284 8774 23336 8780
rect 23296 8498 23324 8774
rect 23388 8537 23416 12582
rect 23468 12232 23520 12238
rect 23468 12174 23520 12180
rect 23480 11286 23508 12174
rect 23817 11996 24113 12016
rect 23873 11994 23897 11996
rect 23953 11994 23977 11996
rect 24033 11994 24057 11996
rect 23895 11942 23897 11994
rect 23959 11942 23971 11994
rect 24033 11942 24035 11994
rect 23873 11940 23897 11942
rect 23953 11940 23977 11942
rect 24033 11940 24057 11942
rect 23817 11920 24113 11940
rect 24204 11620 24256 11626
rect 24204 11562 24256 11568
rect 23468 11280 23520 11286
rect 23468 11222 23520 11228
rect 23468 11144 23520 11150
rect 23468 11086 23520 11092
rect 23374 8528 23430 8537
rect 23284 8492 23336 8498
rect 23374 8463 23430 8472
rect 23284 8434 23336 8440
rect 23190 8120 23246 8129
rect 23190 8055 23246 8064
rect 23192 8016 23244 8022
rect 23192 7958 23244 7964
rect 23100 7880 23152 7886
rect 23100 7822 23152 7828
rect 23008 7404 23060 7410
rect 23008 7346 23060 7352
rect 23112 7274 23140 7822
rect 23204 7546 23232 7958
rect 23296 7886 23324 8434
rect 23376 8356 23428 8362
rect 23376 8298 23428 8304
rect 23284 7880 23336 7886
rect 23284 7822 23336 7828
rect 23192 7540 23244 7546
rect 23192 7482 23244 7488
rect 23388 7342 23416 8298
rect 23376 7336 23428 7342
rect 23376 7278 23428 7284
rect 23100 7268 23152 7274
rect 23100 7210 23152 7216
rect 23190 7168 23246 7177
rect 23190 7103 23246 7112
rect 22824 6860 22876 6866
rect 22824 6802 22876 6808
rect 23006 6352 23062 6361
rect 23006 6287 23008 6296
rect 23060 6287 23062 6296
rect 23008 6258 23060 6264
rect 23100 5772 23152 5778
rect 23100 5714 23152 5720
rect 23112 5545 23140 5714
rect 23098 5536 23154 5545
rect 23098 5471 23154 5480
rect 23112 5370 23140 5471
rect 23100 5364 23152 5370
rect 23100 5306 23152 5312
rect 23204 4826 23232 7103
rect 23388 7002 23416 7278
rect 23376 6996 23428 7002
rect 23376 6938 23428 6944
rect 23192 4820 23244 4826
rect 23192 4762 23244 4768
rect 23006 4040 23062 4049
rect 23006 3975 23008 3984
rect 23060 3975 23062 3984
rect 23008 3946 23060 3952
rect 23480 2650 23508 11086
rect 24216 11082 24244 11562
rect 24388 11280 24440 11286
rect 24388 11222 24440 11228
rect 24204 11076 24256 11082
rect 24204 11018 24256 11024
rect 23817 10908 24113 10928
rect 23873 10906 23897 10908
rect 23953 10906 23977 10908
rect 24033 10906 24057 10908
rect 23895 10854 23897 10906
rect 23959 10854 23971 10906
rect 24033 10854 24035 10906
rect 23873 10852 23897 10854
rect 23953 10852 23977 10854
rect 24033 10852 24057 10854
rect 23817 10832 24113 10852
rect 24216 10674 24244 11018
rect 24400 10810 24428 11222
rect 24756 11008 24808 11014
rect 24756 10950 24808 10956
rect 24768 10810 24796 10950
rect 24388 10804 24440 10810
rect 24388 10746 24440 10752
rect 24756 10804 24808 10810
rect 24756 10746 24808 10752
rect 24204 10668 24256 10674
rect 24204 10610 24256 10616
rect 23928 10532 23980 10538
rect 23928 10474 23980 10480
rect 23652 10192 23704 10198
rect 23652 10134 23704 10140
rect 23664 9704 23692 10134
rect 23940 10062 23968 10474
rect 24216 10266 24244 10610
rect 24204 10260 24256 10266
rect 24204 10202 24256 10208
rect 23928 10056 23980 10062
rect 23928 9998 23980 10004
rect 23817 9820 24113 9840
rect 23873 9818 23897 9820
rect 23953 9818 23977 9820
rect 24033 9818 24057 9820
rect 23895 9766 23897 9818
rect 23959 9766 23971 9818
rect 24033 9766 24035 9818
rect 23873 9764 23897 9766
rect 23953 9764 23977 9766
rect 24033 9764 24057 9766
rect 23817 9744 24113 9764
rect 24294 9752 24350 9761
rect 24204 9716 24256 9722
rect 23664 9676 23784 9704
rect 23650 9616 23706 9625
rect 23756 9586 23784 9676
rect 24294 9687 24350 9696
rect 24662 9752 24718 9761
rect 24662 9687 24718 9696
rect 24204 9658 24256 9664
rect 23650 9551 23706 9560
rect 23744 9580 23796 9586
rect 23664 9466 23692 9551
rect 23744 9522 23796 9528
rect 23664 9438 23784 9466
rect 23560 8900 23612 8906
rect 23560 8842 23612 8848
rect 23572 8498 23600 8842
rect 23560 8492 23612 8498
rect 23560 8434 23612 8440
rect 23572 6866 23600 8434
rect 23650 7984 23706 7993
rect 23650 7919 23706 7928
rect 23560 6860 23612 6866
rect 23560 6802 23612 6808
rect 23572 6458 23600 6802
rect 23560 6452 23612 6458
rect 23560 6394 23612 6400
rect 23664 5642 23692 7919
rect 23652 5636 23704 5642
rect 23652 5578 23704 5584
rect 23756 5370 23784 9438
rect 23817 8732 24113 8752
rect 23873 8730 23897 8732
rect 23953 8730 23977 8732
rect 24033 8730 24057 8732
rect 23895 8678 23897 8730
rect 23959 8678 23971 8730
rect 24033 8678 24035 8730
rect 23873 8676 23897 8678
rect 23953 8676 23977 8678
rect 24033 8676 24057 8678
rect 23817 8656 24113 8676
rect 23817 7644 24113 7664
rect 23873 7642 23897 7644
rect 23953 7642 23977 7644
rect 24033 7642 24057 7644
rect 23895 7590 23897 7642
rect 23959 7590 23971 7642
rect 24033 7590 24035 7642
rect 23873 7588 23897 7590
rect 23953 7588 23977 7590
rect 24033 7588 24057 7590
rect 23817 7568 24113 7588
rect 24216 7546 24244 9658
rect 24308 9602 24336 9687
rect 24388 9648 24440 9654
rect 24308 9596 24388 9602
rect 24308 9590 24440 9596
rect 24308 9574 24428 9590
rect 24676 9178 24704 9687
rect 24664 9172 24716 9178
rect 24664 9114 24716 9120
rect 24388 9036 24440 9042
rect 24860 9024 24888 12815
rect 25766 11792 25822 11801
rect 25766 11727 25822 11736
rect 25122 10840 25178 10849
rect 25122 10775 25124 10784
rect 25176 10775 25178 10784
rect 25124 10746 25176 10752
rect 24940 10600 24992 10606
rect 24938 10568 24940 10577
rect 24992 10568 24994 10577
rect 24938 10503 24994 10512
rect 25780 9722 25808 11727
rect 25768 9716 25820 9722
rect 25768 9658 25820 9664
rect 24388 8978 24440 8984
rect 24676 8996 24888 9024
rect 24400 8362 24428 8978
rect 24388 8356 24440 8362
rect 24308 8316 24388 8344
rect 24204 7540 24256 7546
rect 24204 7482 24256 7488
rect 24204 7200 24256 7206
rect 24204 7142 24256 7148
rect 23817 6556 24113 6576
rect 23873 6554 23897 6556
rect 23953 6554 23977 6556
rect 24033 6554 24057 6556
rect 23895 6502 23897 6554
rect 23959 6502 23971 6554
rect 24033 6502 24035 6554
rect 23873 6500 23897 6502
rect 23953 6500 23977 6502
rect 24033 6500 24057 6502
rect 23817 6480 24113 6500
rect 24216 6390 24244 7142
rect 24308 6866 24336 8316
rect 24388 8298 24440 8304
rect 24676 8090 24704 8996
rect 24938 8800 24994 8809
rect 24938 8735 24994 8744
rect 24952 8634 24980 8735
rect 24940 8628 24992 8634
rect 24940 8570 24992 8576
rect 24754 8528 24810 8537
rect 24754 8463 24810 8472
rect 24768 8430 24796 8463
rect 24756 8424 24808 8430
rect 24756 8366 24808 8372
rect 24664 8084 24716 8090
rect 24664 8026 24716 8032
rect 24572 7948 24624 7954
rect 24572 7890 24624 7896
rect 24480 7336 24532 7342
rect 24480 7278 24532 7284
rect 24388 7268 24440 7274
rect 24388 7210 24440 7216
rect 24296 6860 24348 6866
rect 24296 6802 24348 6808
rect 24400 6730 24428 7210
rect 24388 6724 24440 6730
rect 24388 6666 24440 6672
rect 24492 6610 24520 7278
rect 24584 7206 24612 7890
rect 24754 7712 24810 7721
rect 24754 7647 24810 7656
rect 24572 7200 24624 7206
rect 24572 7142 24624 7148
rect 24308 6582 24520 6610
rect 24204 6384 24256 6390
rect 24204 6326 24256 6332
rect 24308 5914 24336 6582
rect 24768 6458 24796 7647
rect 25124 6860 25176 6866
rect 25124 6802 25176 6808
rect 25030 6624 25086 6633
rect 25030 6559 25086 6568
rect 24756 6452 24808 6458
rect 24756 6394 24808 6400
rect 24768 6254 24796 6394
rect 24756 6248 24808 6254
rect 24756 6190 24808 6196
rect 24296 5908 24348 5914
rect 24296 5850 24348 5856
rect 25044 5778 25072 6559
rect 25136 6118 25164 6802
rect 25124 6112 25176 6118
rect 25124 6054 25176 6060
rect 25766 6080 25822 6089
rect 25032 5772 25084 5778
rect 25032 5714 25084 5720
rect 24662 5536 24718 5545
rect 23817 5468 24113 5488
rect 24662 5471 24718 5480
rect 23873 5466 23897 5468
rect 23953 5466 23977 5468
rect 24033 5466 24057 5468
rect 23895 5414 23897 5466
rect 23959 5414 23971 5466
rect 24033 5414 24035 5466
rect 23873 5412 23897 5414
rect 23953 5412 23977 5414
rect 24033 5412 24057 5414
rect 23817 5392 24113 5412
rect 24676 5370 24704 5471
rect 25044 5370 25072 5714
rect 23744 5364 23796 5370
rect 23744 5306 23796 5312
rect 24664 5364 24716 5370
rect 24664 5306 24716 5312
rect 25032 5364 25084 5370
rect 25032 5306 25084 5312
rect 24676 5166 24704 5306
rect 24664 5160 24716 5166
rect 24664 5102 24716 5108
rect 24204 4684 24256 4690
rect 24204 4626 24256 4632
rect 24216 4593 24244 4626
rect 24202 4584 24258 4593
rect 24202 4519 24258 4528
rect 25030 4584 25086 4593
rect 25030 4519 25086 4528
rect 23817 4380 24113 4400
rect 23873 4378 23897 4380
rect 23953 4378 23977 4380
rect 24033 4378 24057 4380
rect 23895 4326 23897 4378
rect 23959 4326 23971 4378
rect 24033 4326 24035 4378
rect 23873 4324 23897 4326
rect 23953 4324 23977 4326
rect 24033 4324 24057 4326
rect 23817 4304 24113 4324
rect 25044 4146 25072 4519
rect 25032 4140 25084 4146
rect 25032 4082 25084 4088
rect 24664 3936 24716 3942
rect 24664 3878 24716 3884
rect 24676 3505 24704 3878
rect 24662 3496 24718 3505
rect 24662 3431 24718 3440
rect 23817 3292 24113 3312
rect 23873 3290 23897 3292
rect 23953 3290 23977 3292
rect 24033 3290 24057 3292
rect 23895 3238 23897 3290
rect 23959 3238 23971 3290
rect 24033 3238 24035 3290
rect 23873 3236 23897 3238
rect 23953 3236 23977 3238
rect 24033 3236 24057 3238
rect 23817 3216 24113 3236
rect 23468 2644 23520 2650
rect 23468 2586 23520 2592
rect 24664 2508 24716 2514
rect 24664 2450 24716 2456
rect 24676 2310 24704 2450
rect 24664 2304 24716 2310
rect 24664 2246 24716 2252
rect 23817 2204 24113 2224
rect 23873 2202 23897 2204
rect 23953 2202 23977 2204
rect 24033 2202 24057 2204
rect 23895 2150 23897 2202
rect 23959 2150 23971 2202
rect 24033 2150 24035 2202
rect 23873 2148 23897 2150
rect 23953 2148 23977 2150
rect 24033 2148 24057 2150
rect 23817 2128 24113 2148
rect 24676 1465 24704 2246
rect 24662 1456 24718 1465
rect 24662 1391 24718 1400
rect 25136 513 25164 6054
rect 25766 6015 25822 6024
rect 25122 504 25178 513
rect 1294 0 1350 480
rect 4790 0 4846 480
rect 8286 0 8342 480
rect 11782 0 11838 480
rect 15278 0 15334 480
rect 18774 0 18830 480
rect 22270 0 22326 480
rect 25780 480 25808 6015
rect 25122 439 25178 448
rect 25766 0 25822 480
<< via2 >>
rect 6 24248 62 24304
rect 1938 24112 1994 24168
rect 3594 23568 3650 23624
rect 5150 25050 5206 25052
rect 5230 25050 5286 25052
rect 5310 25050 5366 25052
rect 5390 25050 5446 25052
rect 5150 24998 5176 25050
rect 5176 24998 5206 25050
rect 5230 24998 5240 25050
rect 5240 24998 5286 25050
rect 5310 24998 5356 25050
rect 5356 24998 5366 25050
rect 5390 24998 5420 25050
rect 5420 24998 5446 25050
rect 5150 24996 5206 24998
rect 5230 24996 5286 24998
rect 5310 24996 5366 24998
rect 5390 24996 5446 24998
rect 5150 23962 5206 23964
rect 5230 23962 5286 23964
rect 5310 23962 5366 23964
rect 5390 23962 5446 23964
rect 5150 23910 5176 23962
rect 5176 23910 5206 23962
rect 5230 23910 5240 23962
rect 5240 23910 5286 23962
rect 5310 23910 5356 23962
rect 5356 23910 5366 23962
rect 5390 23910 5420 23962
rect 5420 23910 5446 23962
rect 5150 23908 5206 23910
rect 5230 23908 5286 23910
rect 5310 23908 5366 23910
rect 5390 23908 5446 23910
rect 4974 23024 5030 23080
rect 5150 22874 5206 22876
rect 5230 22874 5286 22876
rect 5310 22874 5366 22876
rect 5390 22874 5446 22876
rect 5150 22822 5176 22874
rect 5176 22822 5206 22874
rect 5230 22822 5240 22874
rect 5240 22822 5286 22874
rect 5310 22822 5356 22874
rect 5356 22822 5366 22874
rect 5390 22822 5420 22874
rect 5420 22822 5446 22874
rect 5150 22820 5206 22822
rect 5230 22820 5286 22822
rect 5310 22820 5366 22822
rect 5390 22820 5446 22822
rect 8378 24248 8434 24304
rect 9817 25594 9873 25596
rect 9897 25594 9953 25596
rect 9977 25594 10033 25596
rect 10057 25594 10113 25596
rect 9817 25542 9843 25594
rect 9843 25542 9873 25594
rect 9897 25542 9907 25594
rect 9907 25542 9953 25594
rect 9977 25542 10023 25594
rect 10023 25542 10033 25594
rect 10057 25542 10087 25594
rect 10087 25542 10113 25594
rect 9817 25540 9873 25542
rect 9897 25540 9953 25542
rect 9977 25540 10033 25542
rect 10057 25540 10113 25542
rect 9817 24506 9873 24508
rect 9897 24506 9953 24508
rect 9977 24506 10033 24508
rect 10057 24506 10113 24508
rect 9817 24454 9843 24506
rect 9843 24454 9873 24506
rect 9897 24454 9907 24506
rect 9907 24454 9953 24506
rect 9977 24454 10023 24506
rect 10023 24454 10033 24506
rect 10057 24454 10087 24506
rect 10087 24454 10113 24506
rect 9817 24452 9873 24454
rect 9897 24452 9953 24454
rect 9977 24452 10033 24454
rect 10057 24452 10113 24454
rect 7734 23160 7790 23216
rect 6262 21936 6318 21992
rect 5150 21786 5206 21788
rect 5230 21786 5286 21788
rect 5310 21786 5366 21788
rect 5390 21786 5446 21788
rect 5150 21734 5176 21786
rect 5176 21734 5206 21786
rect 5230 21734 5240 21786
rect 5240 21734 5286 21786
rect 5310 21734 5356 21786
rect 5356 21734 5366 21786
rect 5390 21734 5420 21786
rect 5420 21734 5446 21786
rect 5150 21732 5206 21734
rect 5230 21732 5286 21734
rect 5310 21732 5366 21734
rect 5390 21732 5446 21734
rect 2214 21528 2270 21584
rect 7458 21548 7514 21584
rect 7458 21528 7460 21548
rect 7460 21528 7512 21548
rect 7512 21528 7514 21548
rect 5150 20698 5206 20700
rect 5230 20698 5286 20700
rect 5310 20698 5366 20700
rect 5390 20698 5446 20700
rect 5150 20646 5176 20698
rect 5176 20646 5206 20698
rect 5230 20646 5240 20698
rect 5240 20646 5286 20698
rect 5310 20646 5356 20698
rect 5356 20646 5366 20698
rect 5390 20646 5420 20698
rect 5420 20646 5446 20698
rect 5150 20644 5206 20646
rect 5230 20644 5286 20646
rect 5310 20644 5366 20646
rect 5390 20644 5446 20646
rect 4974 19896 5030 19952
rect 5150 19610 5206 19612
rect 5230 19610 5286 19612
rect 5310 19610 5366 19612
rect 5390 19610 5446 19612
rect 5150 19558 5176 19610
rect 5176 19558 5206 19610
rect 5230 19558 5240 19610
rect 5240 19558 5286 19610
rect 5310 19558 5356 19610
rect 5356 19558 5366 19610
rect 5390 19558 5420 19610
rect 5420 19558 5446 19610
rect 5150 19556 5206 19558
rect 5230 19556 5286 19558
rect 5310 19556 5366 19558
rect 5390 19556 5446 19558
rect 5150 18522 5206 18524
rect 5230 18522 5286 18524
rect 5310 18522 5366 18524
rect 5390 18522 5446 18524
rect 5150 18470 5176 18522
rect 5176 18470 5206 18522
rect 5230 18470 5240 18522
rect 5240 18470 5286 18522
rect 5310 18470 5356 18522
rect 5356 18470 5366 18522
rect 5390 18470 5420 18522
rect 5420 18470 5446 18522
rect 5150 18468 5206 18470
rect 5230 18468 5286 18470
rect 5310 18468 5366 18470
rect 5390 18468 5446 18470
rect 5150 17434 5206 17436
rect 5230 17434 5286 17436
rect 5310 17434 5366 17436
rect 5390 17434 5446 17436
rect 5150 17382 5176 17434
rect 5176 17382 5206 17434
rect 5230 17382 5240 17434
rect 5240 17382 5286 17434
rect 5310 17382 5356 17434
rect 5356 17382 5366 17434
rect 5390 17382 5420 17434
rect 5420 17382 5446 17434
rect 5150 17380 5206 17382
rect 5230 17380 5286 17382
rect 5310 17380 5366 17382
rect 5390 17380 5446 17382
rect 5150 16346 5206 16348
rect 5230 16346 5286 16348
rect 5310 16346 5366 16348
rect 5390 16346 5446 16348
rect 5150 16294 5176 16346
rect 5176 16294 5206 16346
rect 5230 16294 5240 16346
rect 5240 16294 5286 16346
rect 5310 16294 5356 16346
rect 5356 16294 5366 16346
rect 5390 16294 5420 16346
rect 5420 16294 5446 16346
rect 5150 16292 5206 16294
rect 5230 16292 5286 16294
rect 5310 16292 5366 16294
rect 5390 16292 5446 16294
rect 5150 15258 5206 15260
rect 5230 15258 5286 15260
rect 5310 15258 5366 15260
rect 5390 15258 5446 15260
rect 5150 15206 5176 15258
rect 5176 15206 5206 15258
rect 5230 15206 5240 15258
rect 5240 15206 5286 15258
rect 5310 15206 5356 15258
rect 5356 15206 5366 15258
rect 5390 15206 5420 15258
rect 5420 15206 5446 15258
rect 5150 15204 5206 15206
rect 5230 15204 5286 15206
rect 5310 15204 5366 15206
rect 5390 15204 5446 15206
rect 5150 14170 5206 14172
rect 5230 14170 5286 14172
rect 5310 14170 5366 14172
rect 5390 14170 5446 14172
rect 5150 14118 5176 14170
rect 5176 14118 5206 14170
rect 5230 14118 5240 14170
rect 5240 14118 5286 14170
rect 5310 14118 5356 14170
rect 5356 14118 5366 14170
rect 5390 14118 5420 14170
rect 5420 14118 5446 14170
rect 5150 14116 5206 14118
rect 5230 14116 5286 14118
rect 5310 14116 5366 14118
rect 5390 14116 5446 14118
rect 5150 13082 5206 13084
rect 5230 13082 5286 13084
rect 5310 13082 5366 13084
rect 5390 13082 5446 13084
rect 5150 13030 5176 13082
rect 5176 13030 5206 13082
rect 5230 13030 5240 13082
rect 5240 13030 5286 13082
rect 5310 13030 5356 13082
rect 5356 13030 5366 13082
rect 5390 13030 5420 13082
rect 5420 13030 5446 13082
rect 5150 13028 5206 13030
rect 5230 13028 5286 13030
rect 5310 13028 5366 13030
rect 5390 13028 5446 13030
rect 5150 11994 5206 11996
rect 5230 11994 5286 11996
rect 5310 11994 5366 11996
rect 5390 11994 5446 11996
rect 5150 11942 5176 11994
rect 5176 11942 5206 11994
rect 5230 11942 5240 11994
rect 5240 11942 5286 11994
rect 5310 11942 5356 11994
rect 5356 11942 5366 11994
rect 5390 11942 5420 11994
rect 5420 11942 5446 11994
rect 5150 11940 5206 11942
rect 5230 11940 5286 11942
rect 5310 11940 5366 11942
rect 5390 11940 5446 11942
rect 5150 10906 5206 10908
rect 5230 10906 5286 10908
rect 5310 10906 5366 10908
rect 5390 10906 5446 10908
rect 5150 10854 5176 10906
rect 5176 10854 5206 10906
rect 5230 10854 5240 10906
rect 5240 10854 5286 10906
rect 5310 10854 5356 10906
rect 5356 10854 5366 10906
rect 5390 10854 5420 10906
rect 5420 10854 5446 10906
rect 5150 10852 5206 10854
rect 5230 10852 5286 10854
rect 5310 10852 5366 10854
rect 5390 10852 5446 10854
rect 5150 9818 5206 9820
rect 5230 9818 5286 9820
rect 5310 9818 5366 9820
rect 5390 9818 5446 9820
rect 5150 9766 5176 9818
rect 5176 9766 5206 9818
rect 5230 9766 5240 9818
rect 5240 9766 5286 9818
rect 5310 9766 5356 9818
rect 5356 9766 5366 9818
rect 5390 9766 5420 9818
rect 5420 9766 5446 9818
rect 5150 9764 5206 9766
rect 5230 9764 5286 9766
rect 5310 9764 5366 9766
rect 5390 9764 5446 9766
rect 5150 8730 5206 8732
rect 5230 8730 5286 8732
rect 5310 8730 5366 8732
rect 5390 8730 5446 8732
rect 5150 8678 5176 8730
rect 5176 8678 5206 8730
rect 5230 8678 5240 8730
rect 5240 8678 5286 8730
rect 5310 8678 5356 8730
rect 5356 8678 5366 8730
rect 5390 8678 5420 8730
rect 5420 8678 5446 8730
rect 5150 8676 5206 8678
rect 5230 8676 5286 8678
rect 5310 8676 5366 8678
rect 5390 8676 5446 8678
rect 9022 19760 9078 19816
rect 9206 18672 9262 18728
rect 10954 24248 11010 24304
rect 10862 24112 10918 24168
rect 9817 23418 9873 23420
rect 9897 23418 9953 23420
rect 9977 23418 10033 23420
rect 10057 23418 10113 23420
rect 9817 23366 9843 23418
rect 9843 23366 9873 23418
rect 9897 23366 9907 23418
rect 9907 23366 9953 23418
rect 9977 23366 10023 23418
rect 10023 23366 10033 23418
rect 10057 23366 10087 23418
rect 10087 23366 10113 23418
rect 9817 23364 9873 23366
rect 9897 23364 9953 23366
rect 9977 23364 10033 23366
rect 10057 23364 10113 23366
rect 9817 22330 9873 22332
rect 9897 22330 9953 22332
rect 9977 22330 10033 22332
rect 10057 22330 10113 22332
rect 9817 22278 9843 22330
rect 9843 22278 9873 22330
rect 9897 22278 9907 22330
rect 9907 22278 9953 22330
rect 9977 22278 10023 22330
rect 10023 22278 10033 22330
rect 10057 22278 10087 22330
rect 10087 22278 10113 22330
rect 9817 22276 9873 22278
rect 9897 22276 9953 22278
rect 9977 22276 10033 22278
rect 10057 22276 10113 22278
rect 9817 21242 9873 21244
rect 9897 21242 9953 21244
rect 9977 21242 10033 21244
rect 10057 21242 10113 21244
rect 9817 21190 9843 21242
rect 9843 21190 9873 21242
rect 9897 21190 9907 21242
rect 9907 21190 9953 21242
rect 9977 21190 10023 21242
rect 10023 21190 10033 21242
rect 10057 21190 10087 21242
rect 10087 21190 10113 21242
rect 9817 21188 9873 21190
rect 9897 21188 9953 21190
rect 9977 21188 10033 21190
rect 10057 21188 10113 21190
rect 9482 18672 9538 18728
rect 9574 18572 9576 18592
rect 9576 18572 9628 18592
rect 9628 18572 9630 18592
rect 9574 18536 9630 18572
rect 9817 20154 9873 20156
rect 9897 20154 9953 20156
rect 9977 20154 10033 20156
rect 10057 20154 10113 20156
rect 9817 20102 9843 20154
rect 9843 20102 9873 20154
rect 9897 20102 9907 20154
rect 9907 20102 9953 20154
rect 9977 20102 10023 20154
rect 10023 20102 10033 20154
rect 10057 20102 10087 20154
rect 10087 20102 10113 20154
rect 9817 20100 9873 20102
rect 9897 20100 9953 20102
rect 9977 20100 10033 20102
rect 10057 20100 10113 20102
rect 9817 19066 9873 19068
rect 9897 19066 9953 19068
rect 9977 19066 10033 19068
rect 10057 19066 10113 19068
rect 9817 19014 9843 19066
rect 9843 19014 9873 19066
rect 9897 19014 9907 19066
rect 9907 19014 9953 19066
rect 9977 19014 10023 19066
rect 10023 19014 10033 19066
rect 10057 19014 10087 19066
rect 10087 19014 10113 19066
rect 9817 19012 9873 19014
rect 9897 19012 9953 19014
rect 9977 19012 10033 19014
rect 10057 19012 10113 19014
rect 9817 17978 9873 17980
rect 9897 17978 9953 17980
rect 9977 17978 10033 17980
rect 10057 17978 10113 17980
rect 9817 17926 9843 17978
rect 9843 17926 9873 17978
rect 9897 17926 9907 17978
rect 9907 17926 9953 17978
rect 9977 17926 10023 17978
rect 10023 17926 10033 17978
rect 10057 17926 10087 17978
rect 10087 17926 10113 17978
rect 9817 17924 9873 17926
rect 9897 17924 9953 17926
rect 9977 17924 10033 17926
rect 10057 17924 10113 17926
rect 9817 16890 9873 16892
rect 9897 16890 9953 16892
rect 9977 16890 10033 16892
rect 10057 16890 10113 16892
rect 9817 16838 9843 16890
rect 9843 16838 9873 16890
rect 9897 16838 9907 16890
rect 9907 16838 9953 16890
rect 9977 16838 10023 16890
rect 10023 16838 10033 16890
rect 10057 16838 10087 16890
rect 10087 16838 10113 16890
rect 9817 16836 9873 16838
rect 9897 16836 9953 16838
rect 9977 16836 10033 16838
rect 10057 16836 10113 16838
rect 10218 15852 10220 15872
rect 10220 15852 10272 15872
rect 10272 15852 10274 15872
rect 10218 15816 10274 15852
rect 9817 15802 9873 15804
rect 9897 15802 9953 15804
rect 9977 15802 10033 15804
rect 10057 15802 10113 15804
rect 9817 15750 9843 15802
rect 9843 15750 9873 15802
rect 9897 15750 9907 15802
rect 9907 15750 9953 15802
rect 9977 15750 10023 15802
rect 10023 15750 10033 15802
rect 10057 15750 10087 15802
rect 10087 15750 10113 15802
rect 9817 15748 9873 15750
rect 9897 15748 9953 15750
rect 9977 15748 10033 15750
rect 10057 15748 10113 15750
rect 9817 14714 9873 14716
rect 9897 14714 9953 14716
rect 9977 14714 10033 14716
rect 10057 14714 10113 14716
rect 9817 14662 9843 14714
rect 9843 14662 9873 14714
rect 9897 14662 9907 14714
rect 9907 14662 9953 14714
rect 9977 14662 10023 14714
rect 10023 14662 10033 14714
rect 10057 14662 10087 14714
rect 10087 14662 10113 14714
rect 9817 14660 9873 14662
rect 9897 14660 9953 14662
rect 9977 14660 10033 14662
rect 10057 14660 10113 14662
rect 9817 13626 9873 13628
rect 9897 13626 9953 13628
rect 9977 13626 10033 13628
rect 10057 13626 10113 13628
rect 9817 13574 9843 13626
rect 9843 13574 9873 13626
rect 9897 13574 9907 13626
rect 9907 13574 9953 13626
rect 9977 13574 10023 13626
rect 10023 13574 10033 13626
rect 10057 13574 10087 13626
rect 10087 13574 10113 13626
rect 9817 13572 9873 13574
rect 9897 13572 9953 13574
rect 9977 13572 10033 13574
rect 10057 13572 10113 13574
rect 9817 12538 9873 12540
rect 9897 12538 9953 12540
rect 9977 12538 10033 12540
rect 10057 12538 10113 12540
rect 9817 12486 9843 12538
rect 9843 12486 9873 12538
rect 9897 12486 9907 12538
rect 9907 12486 9953 12538
rect 9977 12486 10023 12538
rect 10023 12486 10033 12538
rect 10057 12486 10087 12538
rect 10087 12486 10113 12538
rect 9817 12484 9873 12486
rect 9897 12484 9953 12486
rect 9977 12484 10033 12486
rect 10057 12484 10113 12486
rect 9390 11600 9446 11656
rect 9817 11450 9873 11452
rect 9897 11450 9953 11452
rect 9977 11450 10033 11452
rect 10057 11450 10113 11452
rect 9817 11398 9843 11450
rect 9843 11398 9873 11450
rect 9897 11398 9907 11450
rect 9907 11398 9953 11450
rect 9977 11398 10023 11450
rect 10023 11398 10033 11450
rect 10057 11398 10087 11450
rect 10087 11398 10113 11450
rect 9817 11396 9873 11398
rect 9897 11396 9953 11398
rect 9977 11396 10033 11398
rect 10057 11396 10113 11398
rect 9817 10362 9873 10364
rect 9897 10362 9953 10364
rect 9977 10362 10033 10364
rect 10057 10362 10113 10364
rect 9817 10310 9843 10362
rect 9843 10310 9873 10362
rect 9897 10310 9907 10362
rect 9907 10310 9953 10362
rect 9977 10310 10023 10362
rect 10023 10310 10033 10362
rect 10057 10310 10087 10362
rect 10087 10310 10113 10362
rect 9817 10308 9873 10310
rect 9897 10308 9953 10310
rect 9977 10308 10033 10310
rect 10057 10308 10113 10310
rect 9817 9274 9873 9276
rect 9897 9274 9953 9276
rect 9977 9274 10033 9276
rect 10057 9274 10113 9276
rect 9817 9222 9843 9274
rect 9843 9222 9873 9274
rect 9897 9222 9907 9274
rect 9907 9222 9953 9274
rect 9977 9222 10023 9274
rect 10023 9222 10033 9274
rect 10057 9222 10087 9274
rect 10087 9222 10113 9274
rect 9817 9220 9873 9222
rect 9897 9220 9953 9222
rect 9977 9220 10033 9222
rect 10057 9220 10113 9222
rect 9817 8186 9873 8188
rect 9897 8186 9953 8188
rect 9977 8186 10033 8188
rect 10057 8186 10113 8188
rect 9817 8134 9843 8186
rect 9843 8134 9873 8186
rect 9897 8134 9907 8186
rect 9907 8134 9953 8186
rect 9977 8134 10023 8186
rect 10023 8134 10033 8186
rect 10057 8134 10087 8186
rect 10087 8134 10113 8186
rect 9817 8132 9873 8134
rect 9897 8132 9953 8134
rect 9977 8132 10033 8134
rect 10057 8132 10113 8134
rect 8194 7928 8250 7984
rect 5150 7642 5206 7644
rect 5230 7642 5286 7644
rect 5310 7642 5366 7644
rect 5390 7642 5446 7644
rect 5150 7590 5176 7642
rect 5176 7590 5206 7642
rect 5230 7590 5240 7642
rect 5240 7590 5286 7642
rect 5310 7590 5356 7642
rect 5356 7590 5366 7642
rect 5390 7590 5420 7642
rect 5420 7590 5446 7642
rect 5150 7588 5206 7590
rect 5230 7588 5286 7590
rect 5310 7588 5366 7590
rect 5390 7588 5446 7590
rect 9817 7098 9873 7100
rect 9897 7098 9953 7100
rect 9977 7098 10033 7100
rect 10057 7098 10113 7100
rect 9817 7046 9843 7098
rect 9843 7046 9873 7098
rect 9897 7046 9907 7098
rect 9907 7046 9953 7098
rect 9977 7046 10023 7098
rect 10023 7046 10033 7098
rect 10057 7046 10087 7098
rect 10087 7046 10113 7098
rect 9817 7044 9873 7046
rect 9897 7044 9953 7046
rect 9977 7044 10033 7046
rect 10057 7044 10113 7046
rect 5150 6554 5206 6556
rect 5230 6554 5286 6556
rect 5310 6554 5366 6556
rect 5390 6554 5446 6556
rect 5150 6502 5176 6554
rect 5176 6502 5206 6554
rect 5230 6502 5240 6554
rect 5240 6502 5286 6554
rect 5310 6502 5356 6554
rect 5356 6502 5366 6554
rect 5390 6502 5420 6554
rect 5420 6502 5446 6554
rect 5150 6500 5206 6502
rect 5230 6500 5286 6502
rect 5310 6500 5366 6502
rect 5390 6500 5446 6502
rect 9817 6010 9873 6012
rect 9897 6010 9953 6012
rect 9977 6010 10033 6012
rect 10057 6010 10113 6012
rect 9817 5958 9843 6010
rect 9843 5958 9873 6010
rect 9897 5958 9907 6010
rect 9907 5958 9953 6010
rect 9977 5958 10023 6010
rect 10023 5958 10033 6010
rect 10057 5958 10087 6010
rect 10087 5958 10113 6010
rect 9817 5956 9873 5958
rect 9897 5956 9953 5958
rect 9977 5956 10033 5958
rect 10057 5956 10113 5958
rect 8286 5752 8342 5808
rect 5150 5466 5206 5468
rect 5230 5466 5286 5468
rect 5310 5466 5366 5468
rect 5390 5466 5446 5468
rect 5150 5414 5176 5466
rect 5176 5414 5206 5466
rect 5230 5414 5240 5466
rect 5240 5414 5286 5466
rect 5310 5414 5356 5466
rect 5356 5414 5366 5466
rect 5390 5414 5420 5466
rect 5420 5414 5446 5466
rect 5150 5412 5206 5414
rect 5230 5412 5286 5414
rect 5310 5412 5366 5414
rect 5390 5412 5446 5414
rect 5150 4378 5206 4380
rect 5230 4378 5286 4380
rect 5310 4378 5366 4380
rect 5390 4378 5446 4380
rect 5150 4326 5176 4378
rect 5176 4326 5206 4378
rect 5230 4326 5240 4378
rect 5240 4326 5286 4378
rect 5310 4326 5356 4378
rect 5356 4326 5366 4378
rect 5390 4326 5420 4378
rect 5420 4326 5446 4378
rect 5150 4324 5206 4326
rect 5230 4324 5286 4326
rect 5310 4324 5366 4326
rect 5390 4324 5446 4326
rect 4790 3984 4846 4040
rect 1294 3440 1350 3496
rect 5150 3290 5206 3292
rect 5230 3290 5286 3292
rect 5310 3290 5366 3292
rect 5390 3290 5446 3292
rect 5150 3238 5176 3290
rect 5176 3238 5206 3290
rect 5230 3238 5240 3290
rect 5240 3238 5286 3290
rect 5310 3238 5356 3290
rect 5356 3238 5366 3290
rect 5390 3238 5420 3290
rect 5420 3238 5446 3290
rect 5150 3236 5206 3238
rect 5230 3236 5286 3238
rect 5310 3236 5366 3238
rect 5390 3236 5446 3238
rect 5150 2202 5206 2204
rect 5230 2202 5286 2204
rect 5310 2202 5366 2204
rect 5390 2202 5446 2204
rect 5150 2150 5176 2202
rect 5176 2150 5206 2202
rect 5230 2150 5240 2202
rect 5240 2150 5286 2202
rect 5310 2150 5356 2202
rect 5356 2150 5366 2202
rect 5390 2150 5420 2202
rect 5420 2150 5446 2202
rect 5150 2148 5206 2150
rect 5230 2148 5286 2150
rect 5310 2148 5366 2150
rect 5390 2148 5446 2150
rect 10402 16652 10458 16688
rect 10402 16632 10404 16652
rect 10404 16632 10456 16652
rect 10456 16632 10458 16652
rect 10770 16632 10826 16688
rect 10586 16088 10642 16144
rect 10586 15816 10642 15872
rect 10586 11464 10642 11520
rect 10586 11056 10642 11112
rect 10770 11056 10826 11112
rect 10310 5344 10366 5400
rect 9817 4922 9873 4924
rect 9897 4922 9953 4924
rect 9977 4922 10033 4924
rect 10057 4922 10113 4924
rect 9817 4870 9843 4922
rect 9843 4870 9873 4922
rect 9897 4870 9907 4922
rect 9907 4870 9953 4922
rect 9977 4870 10023 4922
rect 10023 4870 10033 4922
rect 10057 4870 10087 4922
rect 10087 4870 10113 4922
rect 9817 4868 9873 4870
rect 9897 4868 9953 4870
rect 9977 4868 10033 4870
rect 10057 4868 10113 4870
rect 9817 3834 9873 3836
rect 9897 3834 9953 3836
rect 9977 3834 10033 3836
rect 10057 3834 10113 3836
rect 9817 3782 9843 3834
rect 9843 3782 9873 3834
rect 9897 3782 9907 3834
rect 9907 3782 9953 3834
rect 9977 3782 10023 3834
rect 10023 3782 10033 3834
rect 10057 3782 10087 3834
rect 10087 3782 10113 3834
rect 9817 3780 9873 3782
rect 9897 3780 9953 3782
rect 9977 3780 10033 3782
rect 10057 3780 10113 3782
rect 11506 19252 11508 19272
rect 11508 19252 11560 19272
rect 11560 19252 11562 19272
rect 11506 19216 11562 19252
rect 11966 18708 11968 18728
rect 11968 18708 12020 18728
rect 12020 18708 12022 18728
rect 11966 18672 12022 18708
rect 14484 25050 14540 25052
rect 14564 25050 14620 25052
rect 14644 25050 14700 25052
rect 14724 25050 14780 25052
rect 14484 24998 14510 25050
rect 14510 24998 14540 25050
rect 14564 24998 14574 25050
rect 14574 24998 14620 25050
rect 14644 24998 14690 25050
rect 14690 24998 14700 25050
rect 14724 24998 14754 25050
rect 14754 24998 14780 25050
rect 14484 24996 14540 24998
rect 14564 24996 14620 24998
rect 14644 24996 14700 24998
rect 14724 24996 14780 24998
rect 14450 24656 14506 24712
rect 15002 24404 15058 24440
rect 15002 24384 15004 24404
rect 15004 24384 15056 24404
rect 15056 24384 15058 24404
rect 14082 23568 14138 23624
rect 12702 20304 12758 20360
rect 13162 19236 13218 19272
rect 13162 19216 13164 19236
rect 13164 19216 13216 19236
rect 13216 19216 13218 19236
rect 13806 18536 13862 18592
rect 14484 23962 14540 23964
rect 14564 23962 14620 23964
rect 14644 23962 14700 23964
rect 14724 23962 14780 23964
rect 14484 23910 14510 23962
rect 14510 23910 14540 23962
rect 14564 23910 14574 23962
rect 14574 23910 14620 23962
rect 14644 23910 14690 23962
rect 14690 23910 14700 23962
rect 14724 23910 14754 23962
rect 14754 23910 14780 23962
rect 14484 23908 14540 23910
rect 14564 23908 14620 23910
rect 14644 23908 14700 23910
rect 14724 23908 14780 23910
rect 14484 22874 14540 22876
rect 14564 22874 14620 22876
rect 14644 22874 14700 22876
rect 14724 22874 14780 22876
rect 14484 22822 14510 22874
rect 14510 22822 14540 22874
rect 14564 22822 14574 22874
rect 14574 22822 14620 22874
rect 14644 22822 14690 22874
rect 14690 22822 14700 22874
rect 14724 22822 14754 22874
rect 14754 22822 14780 22874
rect 14484 22820 14540 22822
rect 14564 22820 14620 22822
rect 14644 22820 14700 22822
rect 14724 22820 14780 22822
rect 14484 21786 14540 21788
rect 14564 21786 14620 21788
rect 14644 21786 14700 21788
rect 14724 21786 14780 21788
rect 14484 21734 14510 21786
rect 14510 21734 14540 21786
rect 14564 21734 14574 21786
rect 14574 21734 14620 21786
rect 14644 21734 14690 21786
rect 14690 21734 14700 21786
rect 14724 21734 14754 21786
rect 14754 21734 14780 21786
rect 14484 21732 14540 21734
rect 14564 21732 14620 21734
rect 14644 21732 14700 21734
rect 14724 21732 14780 21734
rect 14484 20698 14540 20700
rect 14564 20698 14620 20700
rect 14644 20698 14700 20700
rect 14724 20698 14780 20700
rect 14484 20646 14510 20698
rect 14510 20646 14540 20698
rect 14564 20646 14574 20698
rect 14574 20646 14620 20698
rect 14644 20646 14690 20698
rect 14690 20646 14700 20698
rect 14724 20646 14754 20698
rect 14754 20646 14780 20698
rect 14484 20644 14540 20646
rect 14564 20644 14620 20646
rect 14644 20644 14700 20646
rect 14724 20644 14780 20646
rect 14484 19610 14540 19612
rect 14564 19610 14620 19612
rect 14644 19610 14700 19612
rect 14724 19610 14780 19612
rect 14484 19558 14510 19610
rect 14510 19558 14540 19610
rect 14564 19558 14574 19610
rect 14574 19558 14620 19610
rect 14644 19558 14690 19610
rect 14690 19558 14700 19610
rect 14724 19558 14754 19610
rect 14754 19558 14780 19610
rect 14484 19556 14540 19558
rect 14564 19556 14620 19558
rect 14644 19556 14700 19558
rect 14724 19556 14780 19558
rect 15922 21564 15924 21584
rect 15924 21564 15976 21584
rect 15976 21564 15978 21584
rect 15922 21528 15978 21564
rect 14484 18522 14540 18524
rect 14564 18522 14620 18524
rect 14644 18522 14700 18524
rect 14724 18522 14780 18524
rect 14484 18470 14510 18522
rect 14510 18470 14540 18522
rect 14564 18470 14574 18522
rect 14574 18470 14620 18522
rect 14644 18470 14690 18522
rect 14690 18470 14700 18522
rect 14724 18470 14754 18522
rect 14754 18470 14780 18522
rect 14484 18468 14540 18470
rect 14564 18468 14620 18470
rect 14644 18468 14700 18470
rect 14724 18468 14780 18470
rect 13806 16632 13862 16688
rect 13162 16496 13218 16552
rect 14484 17434 14540 17436
rect 14564 17434 14620 17436
rect 14644 17434 14700 17436
rect 14724 17434 14780 17436
rect 14484 17382 14510 17434
rect 14510 17382 14540 17434
rect 14564 17382 14574 17434
rect 14574 17382 14620 17434
rect 14644 17382 14690 17434
rect 14690 17382 14700 17434
rect 14724 17382 14754 17434
rect 14754 17382 14780 17434
rect 14484 17380 14540 17382
rect 14564 17380 14620 17382
rect 14644 17380 14700 17382
rect 14724 17380 14780 17382
rect 14634 17212 14636 17232
rect 14636 17212 14688 17232
rect 14688 17212 14690 17232
rect 14634 17176 14690 17212
rect 14484 16346 14540 16348
rect 14564 16346 14620 16348
rect 14644 16346 14700 16348
rect 14724 16346 14780 16348
rect 14484 16294 14510 16346
rect 14510 16294 14540 16346
rect 14564 16294 14574 16346
rect 14574 16294 14620 16346
rect 14644 16294 14690 16346
rect 14690 16294 14700 16346
rect 14724 16294 14754 16346
rect 14754 16294 14780 16346
rect 14484 16292 14540 16294
rect 14564 16292 14620 16294
rect 14644 16292 14700 16294
rect 14724 16292 14780 16294
rect 15922 17448 15978 17504
rect 14910 16496 14966 16552
rect 16566 24112 16622 24168
rect 16658 23060 16660 23080
rect 16660 23060 16712 23080
rect 16712 23060 16714 23080
rect 16658 23024 16714 23060
rect 16198 17212 16200 17232
rect 16200 17212 16252 17232
rect 16252 17212 16254 17232
rect 16198 17176 16254 17212
rect 14174 15680 14230 15736
rect 14484 15258 14540 15260
rect 14564 15258 14620 15260
rect 14644 15258 14700 15260
rect 14724 15258 14780 15260
rect 14484 15206 14510 15258
rect 14510 15206 14540 15258
rect 14564 15206 14574 15258
rect 14574 15206 14620 15258
rect 14644 15206 14690 15258
rect 14690 15206 14700 15258
rect 14724 15206 14754 15258
rect 14754 15206 14780 15258
rect 14484 15204 14540 15206
rect 14564 15204 14620 15206
rect 14644 15204 14700 15206
rect 14724 15204 14780 15206
rect 14484 14170 14540 14172
rect 14564 14170 14620 14172
rect 14644 14170 14700 14172
rect 14724 14170 14780 14172
rect 14484 14118 14510 14170
rect 14510 14118 14540 14170
rect 14564 14118 14574 14170
rect 14574 14118 14620 14170
rect 14644 14118 14690 14170
rect 14690 14118 14700 14170
rect 14724 14118 14754 14170
rect 14754 14118 14780 14170
rect 14484 14116 14540 14118
rect 14564 14116 14620 14118
rect 14644 14116 14700 14118
rect 14724 14116 14780 14118
rect 13898 13404 13900 13424
rect 13900 13404 13952 13424
rect 13952 13404 13954 13424
rect 13898 13368 13954 13404
rect 14358 13232 14414 13288
rect 14484 13082 14540 13084
rect 14564 13082 14620 13084
rect 14644 13082 14700 13084
rect 14724 13082 14780 13084
rect 14484 13030 14510 13082
rect 14510 13030 14540 13082
rect 14564 13030 14574 13082
rect 14574 13030 14620 13082
rect 14644 13030 14690 13082
rect 14690 13030 14700 13082
rect 14724 13030 14754 13082
rect 14754 13030 14780 13082
rect 14484 13028 14540 13030
rect 14564 13028 14620 13030
rect 14644 13028 14700 13030
rect 14724 13028 14780 13030
rect 13714 11500 13716 11520
rect 13716 11500 13768 11520
rect 13768 11500 13770 11520
rect 13714 11464 13770 11500
rect 12242 9016 12298 9072
rect 13438 8200 13494 8256
rect 11782 7112 11838 7168
rect 11046 6840 11102 6896
rect 11598 5752 11654 5808
rect 10770 3984 10826 4040
rect 10586 3440 10642 3496
rect 9817 2746 9873 2748
rect 9897 2746 9953 2748
rect 9977 2746 10033 2748
rect 10057 2746 10113 2748
rect 9817 2694 9843 2746
rect 9843 2694 9873 2746
rect 9897 2694 9907 2746
rect 9907 2694 9953 2746
rect 9977 2694 10023 2746
rect 10023 2694 10033 2746
rect 10057 2694 10087 2746
rect 10087 2694 10113 2746
rect 9817 2692 9873 2694
rect 9897 2692 9953 2694
rect 9977 2692 10033 2694
rect 10057 2692 10113 2694
rect 14484 11994 14540 11996
rect 14564 11994 14620 11996
rect 14644 11994 14700 11996
rect 14724 11994 14780 11996
rect 14484 11942 14510 11994
rect 14510 11942 14540 11994
rect 14564 11942 14574 11994
rect 14574 11942 14620 11994
rect 14644 11942 14690 11994
rect 14690 11942 14700 11994
rect 14724 11942 14754 11994
rect 14754 11942 14780 11994
rect 14484 11940 14540 11942
rect 14564 11940 14620 11942
rect 14644 11940 14700 11942
rect 14724 11940 14780 11942
rect 14484 10906 14540 10908
rect 14564 10906 14620 10908
rect 14644 10906 14700 10908
rect 14724 10906 14780 10908
rect 14484 10854 14510 10906
rect 14510 10854 14540 10906
rect 14564 10854 14574 10906
rect 14574 10854 14620 10906
rect 14644 10854 14690 10906
rect 14690 10854 14700 10906
rect 14724 10854 14754 10906
rect 14754 10854 14780 10906
rect 14484 10852 14540 10854
rect 14564 10852 14620 10854
rect 14644 10852 14700 10854
rect 14724 10852 14780 10854
rect 14358 10648 14414 10704
rect 18498 24792 18554 24848
rect 17578 24384 17634 24440
rect 19150 25594 19206 25596
rect 19230 25594 19286 25596
rect 19310 25594 19366 25596
rect 19390 25594 19446 25596
rect 19150 25542 19176 25594
rect 19176 25542 19206 25594
rect 19230 25542 19240 25594
rect 19240 25542 19286 25594
rect 19310 25542 19356 25594
rect 19356 25542 19366 25594
rect 19390 25542 19420 25594
rect 19420 25542 19446 25594
rect 19150 25540 19206 25542
rect 19230 25540 19286 25542
rect 19310 25540 19366 25542
rect 19390 25540 19446 25542
rect 20706 24792 20762 24848
rect 19602 24656 19658 24712
rect 19150 24506 19206 24508
rect 19230 24506 19286 24508
rect 19310 24506 19366 24508
rect 19390 24506 19446 24508
rect 19150 24454 19176 24506
rect 19176 24454 19206 24506
rect 19230 24454 19240 24506
rect 19240 24454 19286 24506
rect 19310 24454 19356 24506
rect 19356 24454 19366 24506
rect 19390 24454 19420 24506
rect 19420 24454 19446 24506
rect 19150 24452 19206 24454
rect 19230 24452 19286 24454
rect 19310 24452 19366 24454
rect 19390 24452 19446 24454
rect 18590 24248 18646 24304
rect 19694 23860 19750 23896
rect 19694 23840 19696 23860
rect 19696 23840 19748 23860
rect 19748 23840 19750 23860
rect 20614 24248 20670 24304
rect 17670 23044 17726 23080
rect 17670 23024 17672 23044
rect 17672 23024 17724 23044
rect 17724 23024 17726 23044
rect 19150 23418 19206 23420
rect 19230 23418 19286 23420
rect 19310 23418 19366 23420
rect 19390 23418 19446 23420
rect 19150 23366 19176 23418
rect 19176 23366 19206 23418
rect 19230 23366 19240 23418
rect 19240 23366 19286 23418
rect 19310 23366 19356 23418
rect 19356 23366 19366 23418
rect 19390 23366 19420 23418
rect 19420 23366 19446 23418
rect 19150 23364 19206 23366
rect 19230 23364 19286 23366
rect 19310 23364 19366 23366
rect 19390 23364 19446 23366
rect 19150 22330 19206 22332
rect 19230 22330 19286 22332
rect 19310 22330 19366 22332
rect 19390 22330 19446 22332
rect 19150 22278 19176 22330
rect 19176 22278 19206 22330
rect 19230 22278 19240 22330
rect 19240 22278 19286 22330
rect 19310 22278 19356 22330
rect 19356 22278 19366 22330
rect 19390 22278 19420 22330
rect 19420 22278 19446 22330
rect 19150 22276 19206 22278
rect 19230 22276 19286 22278
rect 19310 22276 19366 22278
rect 19390 22276 19446 22278
rect 18590 21412 18646 21448
rect 18590 21392 18592 21412
rect 18592 21392 18644 21412
rect 18644 21392 18646 21412
rect 18498 20984 18554 21040
rect 17670 20576 17726 20632
rect 17670 19916 17726 19952
rect 17670 19896 17672 19916
rect 17672 19896 17724 19916
rect 17724 19896 17726 19916
rect 20798 24112 20854 24168
rect 20522 21972 20524 21992
rect 20524 21972 20576 21992
rect 20576 21972 20578 21992
rect 20522 21936 20578 21972
rect 21442 23196 21444 23216
rect 21444 23196 21496 23216
rect 21496 23196 21498 23216
rect 21442 23160 21498 23196
rect 20430 21392 20486 21448
rect 19150 21242 19206 21244
rect 19230 21242 19286 21244
rect 19310 21242 19366 21244
rect 19390 21242 19446 21244
rect 19150 21190 19176 21242
rect 19176 21190 19206 21242
rect 19230 21190 19240 21242
rect 19240 21190 19286 21242
rect 19310 21190 19356 21242
rect 19356 21190 19366 21242
rect 19390 21190 19420 21242
rect 19420 21190 19446 21242
rect 19150 21188 19206 21190
rect 19230 21188 19286 21190
rect 19310 21188 19366 21190
rect 19390 21188 19446 21190
rect 19150 20154 19206 20156
rect 19230 20154 19286 20156
rect 19310 20154 19366 20156
rect 19390 20154 19446 20156
rect 19150 20102 19176 20154
rect 19176 20102 19206 20154
rect 19230 20102 19240 20154
rect 19240 20102 19286 20154
rect 19310 20102 19356 20154
rect 19356 20102 19366 20154
rect 19390 20102 19420 20154
rect 19420 20102 19446 20154
rect 19150 20100 19206 20102
rect 19230 20100 19286 20102
rect 19310 20100 19366 20102
rect 19390 20100 19446 20102
rect 19150 19066 19206 19068
rect 19230 19066 19286 19068
rect 19310 19066 19366 19068
rect 19390 19066 19446 19068
rect 19150 19014 19176 19066
rect 19176 19014 19206 19066
rect 19230 19014 19240 19066
rect 19240 19014 19286 19066
rect 19310 19014 19356 19066
rect 19356 19014 19366 19066
rect 19390 19014 19420 19066
rect 19420 19014 19446 19066
rect 19150 19012 19206 19014
rect 19230 19012 19286 19014
rect 19310 19012 19366 19014
rect 19390 19012 19446 19014
rect 20522 20596 20578 20632
rect 20522 20576 20524 20596
rect 20524 20576 20576 20596
rect 20576 20576 20578 20596
rect 22270 24404 22326 24440
rect 22270 24384 22272 24404
rect 22272 24384 22324 24404
rect 22324 24384 22326 24404
rect 24294 26288 24350 26344
rect 23817 25050 23873 25052
rect 23897 25050 23953 25052
rect 23977 25050 24033 25052
rect 24057 25050 24113 25052
rect 23817 24998 23843 25050
rect 23843 24998 23873 25050
rect 23897 24998 23907 25050
rect 23907 24998 23953 25050
rect 23977 24998 24023 25050
rect 24023 24998 24033 25050
rect 24057 24998 24087 25050
rect 24087 24998 24113 25050
rect 23817 24996 23873 24998
rect 23897 24996 23953 24998
rect 23977 24996 24033 24998
rect 24057 24996 24113 24998
rect 24570 25336 24626 25392
rect 23742 24384 23798 24440
rect 23817 23962 23873 23964
rect 23897 23962 23953 23964
rect 23977 23962 24033 23964
rect 24057 23962 24113 23964
rect 23817 23910 23843 23962
rect 23843 23910 23873 23962
rect 23897 23910 23907 23962
rect 23907 23910 23953 23962
rect 23977 23910 24023 23962
rect 24023 23910 24033 23962
rect 24057 23910 24087 23962
rect 24087 23910 24113 23962
rect 23817 23908 23873 23910
rect 23897 23908 23953 23910
rect 23977 23908 24033 23910
rect 24057 23908 24113 23910
rect 22730 23840 22786 23896
rect 24478 24248 24534 24304
rect 25398 27376 25454 27432
rect 24294 23432 24350 23488
rect 23817 22874 23873 22876
rect 23897 22874 23953 22876
rect 23977 22874 24033 22876
rect 24057 22874 24113 22876
rect 23817 22822 23843 22874
rect 23843 22822 23873 22874
rect 23897 22822 23907 22874
rect 23907 22822 23953 22874
rect 23977 22822 24023 22874
rect 24023 22822 24033 22874
rect 24057 22822 24087 22874
rect 24087 22822 24113 22874
rect 23817 22820 23873 22822
rect 23897 22820 23953 22822
rect 23977 22820 24033 22822
rect 24057 22820 24113 22822
rect 23817 21786 23873 21788
rect 23897 21786 23953 21788
rect 23977 21786 24033 21788
rect 24057 21786 24113 21788
rect 23817 21734 23843 21786
rect 23843 21734 23873 21786
rect 23897 21734 23907 21786
rect 23907 21734 23953 21786
rect 23977 21734 24023 21786
rect 24023 21734 24033 21786
rect 24057 21734 24087 21786
rect 24087 21734 24113 21786
rect 23817 21732 23873 21734
rect 23897 21732 23953 21734
rect 23977 21732 24033 21734
rect 24057 21732 24113 21734
rect 19150 17978 19206 17980
rect 19230 17978 19286 17980
rect 19310 17978 19366 17980
rect 19390 17978 19446 17980
rect 19150 17926 19176 17978
rect 19176 17926 19206 17978
rect 19230 17926 19240 17978
rect 19240 17926 19286 17978
rect 19310 17926 19356 17978
rect 19356 17926 19366 17978
rect 19390 17926 19420 17978
rect 19420 17926 19446 17978
rect 19150 17924 19206 17926
rect 19230 17924 19286 17926
rect 19310 17924 19366 17926
rect 19390 17924 19446 17926
rect 17302 15852 17304 15872
rect 17304 15852 17356 15872
rect 17356 15852 17358 15872
rect 17302 15816 17358 15852
rect 17670 15680 17726 15736
rect 15922 13776 15978 13832
rect 14484 9818 14540 9820
rect 14564 9818 14620 9820
rect 14644 9818 14700 9820
rect 14724 9818 14780 9820
rect 14484 9766 14510 9818
rect 14510 9766 14540 9818
rect 14564 9766 14574 9818
rect 14574 9766 14620 9818
rect 14644 9766 14690 9818
rect 14690 9766 14700 9818
rect 14724 9766 14754 9818
rect 14754 9766 14780 9818
rect 14484 9764 14540 9766
rect 14564 9764 14620 9766
rect 14644 9764 14700 9766
rect 14724 9764 14780 9766
rect 13622 7148 13624 7168
rect 13624 7148 13676 7168
rect 13676 7148 13678 7168
rect 13622 7112 13678 7148
rect 13990 5364 14046 5400
rect 13990 5344 13992 5364
rect 13992 5344 14044 5364
rect 14044 5344 14046 5364
rect 14484 8730 14540 8732
rect 14564 8730 14620 8732
rect 14644 8730 14700 8732
rect 14724 8730 14780 8732
rect 14484 8678 14510 8730
rect 14510 8678 14540 8730
rect 14564 8678 14574 8730
rect 14574 8678 14620 8730
rect 14644 8678 14690 8730
rect 14690 8678 14700 8730
rect 14724 8678 14754 8730
rect 14754 8678 14780 8730
rect 14484 8676 14540 8678
rect 14564 8676 14620 8678
rect 14644 8676 14700 8678
rect 14724 8676 14780 8678
rect 14910 8200 14966 8256
rect 16198 11192 16254 11248
rect 14358 7792 14414 7848
rect 14484 7642 14540 7644
rect 14564 7642 14620 7644
rect 14644 7642 14700 7644
rect 14724 7642 14780 7644
rect 14484 7590 14510 7642
rect 14510 7590 14540 7642
rect 14564 7590 14574 7642
rect 14574 7590 14620 7642
rect 14644 7590 14690 7642
rect 14690 7590 14700 7642
rect 14724 7590 14754 7642
rect 14754 7590 14780 7642
rect 14484 7588 14540 7590
rect 14564 7588 14620 7590
rect 14644 7588 14700 7590
rect 14724 7588 14780 7590
rect 14484 6554 14540 6556
rect 14564 6554 14620 6556
rect 14644 6554 14700 6556
rect 14724 6554 14780 6556
rect 14484 6502 14510 6554
rect 14510 6502 14540 6554
rect 14564 6502 14574 6554
rect 14574 6502 14620 6554
rect 14644 6502 14690 6554
rect 14690 6502 14700 6554
rect 14724 6502 14754 6554
rect 14754 6502 14780 6554
rect 14484 6500 14540 6502
rect 14564 6500 14620 6502
rect 14644 6500 14700 6502
rect 14724 6500 14780 6502
rect 14484 5466 14540 5468
rect 14564 5466 14620 5468
rect 14644 5466 14700 5468
rect 14724 5466 14780 5468
rect 14484 5414 14510 5466
rect 14510 5414 14540 5466
rect 14564 5414 14574 5466
rect 14574 5414 14620 5466
rect 14644 5414 14690 5466
rect 14690 5414 14700 5466
rect 14724 5414 14754 5466
rect 14754 5414 14780 5466
rect 14484 5412 14540 5414
rect 14564 5412 14620 5414
rect 14644 5412 14700 5414
rect 14724 5412 14780 5414
rect 14484 4378 14540 4380
rect 14564 4378 14620 4380
rect 14644 4378 14700 4380
rect 14724 4378 14780 4380
rect 14484 4326 14510 4378
rect 14510 4326 14540 4378
rect 14564 4326 14574 4378
rect 14574 4326 14620 4378
rect 14644 4326 14690 4378
rect 14690 4326 14700 4378
rect 14724 4326 14754 4378
rect 14754 4326 14780 4378
rect 14484 4324 14540 4326
rect 14564 4324 14620 4326
rect 14644 4324 14700 4326
rect 14724 4324 14780 4326
rect 14266 3984 14322 4040
rect 14484 3290 14540 3292
rect 14564 3290 14620 3292
rect 14644 3290 14700 3292
rect 14724 3290 14780 3292
rect 14484 3238 14510 3290
rect 14510 3238 14540 3290
rect 14564 3238 14574 3290
rect 14574 3238 14620 3290
rect 14644 3238 14690 3290
rect 14690 3238 14700 3290
rect 14724 3238 14754 3290
rect 14754 3238 14780 3290
rect 14484 3236 14540 3238
rect 14564 3236 14620 3238
rect 14644 3236 14700 3238
rect 14724 3236 14780 3238
rect 14484 2202 14540 2204
rect 14564 2202 14620 2204
rect 14644 2202 14700 2204
rect 14724 2202 14780 2204
rect 14484 2150 14510 2202
rect 14510 2150 14540 2202
rect 14564 2150 14574 2202
rect 14574 2150 14620 2202
rect 14644 2150 14690 2202
rect 14690 2150 14700 2202
rect 14724 2150 14754 2202
rect 14754 2150 14780 2202
rect 14484 2148 14540 2150
rect 14564 2148 14620 2150
rect 14644 2148 14700 2150
rect 14724 2148 14780 2150
rect 20154 17484 20156 17504
rect 20156 17484 20208 17504
rect 20208 17484 20210 17504
rect 20154 17448 20210 17484
rect 19150 16890 19206 16892
rect 19230 16890 19286 16892
rect 19310 16890 19366 16892
rect 19390 16890 19446 16892
rect 19150 16838 19176 16890
rect 19176 16838 19206 16890
rect 19230 16838 19240 16890
rect 19240 16838 19286 16890
rect 19310 16838 19356 16890
rect 19356 16838 19366 16890
rect 19390 16838 19420 16890
rect 19420 16838 19446 16890
rect 19150 16836 19206 16838
rect 19230 16836 19286 16838
rect 19310 16836 19366 16838
rect 19390 16836 19446 16838
rect 20154 16632 20210 16688
rect 18222 15700 18278 15736
rect 18222 15680 18224 15700
rect 18224 15680 18276 15700
rect 18276 15680 18278 15700
rect 19150 15802 19206 15804
rect 19230 15802 19286 15804
rect 19310 15802 19366 15804
rect 19390 15802 19446 15804
rect 19150 15750 19176 15802
rect 19176 15750 19206 15802
rect 19230 15750 19240 15802
rect 19240 15750 19286 15802
rect 19310 15750 19356 15802
rect 19356 15750 19366 15802
rect 19390 15750 19420 15802
rect 19420 15750 19446 15802
rect 19150 15748 19206 15750
rect 19230 15748 19286 15750
rect 19310 15748 19366 15750
rect 19390 15748 19446 15750
rect 18130 13812 18132 13832
rect 18132 13812 18184 13832
rect 18184 13812 18186 13832
rect 18130 13776 18186 13812
rect 19150 14714 19206 14716
rect 19230 14714 19286 14716
rect 19310 14714 19366 14716
rect 19390 14714 19446 14716
rect 19150 14662 19176 14714
rect 19176 14662 19206 14714
rect 19230 14662 19240 14714
rect 19240 14662 19286 14714
rect 19310 14662 19356 14714
rect 19356 14662 19366 14714
rect 19390 14662 19420 14714
rect 19420 14662 19446 14714
rect 19150 14660 19206 14662
rect 19230 14660 19286 14662
rect 19310 14660 19366 14662
rect 19390 14660 19446 14662
rect 20706 14728 20762 14784
rect 19150 13626 19206 13628
rect 19230 13626 19286 13628
rect 19310 13626 19366 13628
rect 19390 13626 19446 13628
rect 19150 13574 19176 13626
rect 19176 13574 19206 13626
rect 19230 13574 19240 13626
rect 19240 13574 19286 13626
rect 19310 13574 19356 13626
rect 19356 13574 19366 13626
rect 19390 13574 19420 13626
rect 19420 13574 19446 13626
rect 19150 13572 19206 13574
rect 19230 13572 19286 13574
rect 19310 13572 19366 13574
rect 19390 13572 19446 13574
rect 18774 12044 18776 12064
rect 18776 12044 18828 12064
rect 18828 12044 18830 12064
rect 18774 12008 18830 12044
rect 19150 12538 19206 12540
rect 19230 12538 19286 12540
rect 19310 12538 19366 12540
rect 19390 12538 19446 12540
rect 19150 12486 19176 12538
rect 19176 12486 19206 12538
rect 19230 12486 19240 12538
rect 19240 12486 19286 12538
rect 19310 12486 19356 12538
rect 19356 12486 19366 12538
rect 19390 12486 19420 12538
rect 19420 12486 19446 12538
rect 19150 12484 19206 12486
rect 19230 12484 19286 12486
rect 19310 12484 19366 12486
rect 19390 12484 19446 12486
rect 24478 23024 24534 23080
rect 24478 22208 24534 22264
rect 24386 21528 24442 21584
rect 24294 21120 24350 21176
rect 23817 20698 23873 20700
rect 23897 20698 23953 20700
rect 23977 20698 24033 20700
rect 24057 20698 24113 20700
rect 23817 20646 23843 20698
rect 23843 20646 23873 20698
rect 23897 20646 23907 20698
rect 23907 20646 23953 20698
rect 23977 20646 24023 20698
rect 24023 20646 24033 20698
rect 24057 20646 24087 20698
rect 24087 20646 24113 20698
rect 23817 20644 23873 20646
rect 23897 20644 23953 20646
rect 23977 20644 24033 20646
rect 24057 20644 24113 20646
rect 24478 20984 24534 21040
rect 23006 20304 23062 20360
rect 24386 19780 24442 19816
rect 24386 19760 24388 19780
rect 24388 19760 24440 19780
rect 24440 19760 24442 19780
rect 23817 19610 23873 19612
rect 23897 19610 23953 19612
rect 23977 19610 24033 19612
rect 24057 19610 24113 19612
rect 23817 19558 23843 19610
rect 23843 19558 23873 19610
rect 23897 19558 23907 19610
rect 23907 19558 23953 19610
rect 23977 19558 24023 19610
rect 24023 19558 24033 19610
rect 24057 19558 24087 19610
rect 24087 19558 24113 19610
rect 23817 19556 23873 19558
rect 23897 19556 23953 19558
rect 23977 19556 24033 19558
rect 24057 19556 24113 19558
rect 23742 19080 23798 19136
rect 23190 16652 23246 16688
rect 23817 18522 23873 18524
rect 23897 18522 23953 18524
rect 23977 18522 24033 18524
rect 24057 18522 24113 18524
rect 23817 18470 23843 18522
rect 23843 18470 23873 18522
rect 23897 18470 23907 18522
rect 23907 18470 23953 18522
rect 23977 18470 24023 18522
rect 24023 18470 24033 18522
rect 24057 18470 24087 18522
rect 24087 18470 24113 18522
rect 23817 18468 23873 18470
rect 23897 18468 23953 18470
rect 23977 18468 24033 18470
rect 24057 18468 24113 18470
rect 23926 17992 23982 18048
rect 23817 17434 23873 17436
rect 23897 17434 23953 17436
rect 23977 17434 24033 17436
rect 24057 17434 24113 17436
rect 23817 17382 23843 17434
rect 23843 17382 23873 17434
rect 23897 17382 23907 17434
rect 23907 17382 23953 17434
rect 23977 17382 24023 17434
rect 24023 17382 24033 17434
rect 24057 17382 24087 17434
rect 24087 17382 24113 17434
rect 23817 17380 23873 17382
rect 23897 17380 23953 17382
rect 23977 17380 24033 17382
rect 24057 17380 24113 17382
rect 24478 17992 24534 18048
rect 24938 17040 24994 17096
rect 23190 16632 23192 16652
rect 23192 16632 23244 16652
rect 23244 16632 23246 16652
rect 23817 16346 23873 16348
rect 23897 16346 23953 16348
rect 23977 16346 24033 16348
rect 24057 16346 24113 16348
rect 23817 16294 23843 16346
rect 23843 16294 23873 16346
rect 23897 16294 23907 16346
rect 23907 16294 23953 16346
rect 23977 16294 24023 16346
rect 24023 16294 24033 16346
rect 24057 16294 24087 16346
rect 24087 16294 24113 16346
rect 23817 16292 23873 16294
rect 23897 16292 23953 16294
rect 23977 16292 24033 16294
rect 24057 16292 24113 16294
rect 23006 16088 23062 16144
rect 25306 24248 25362 24304
rect 25858 23432 25914 23488
rect 25306 23160 25362 23216
rect 25398 20032 25454 20088
rect 25490 17992 25546 18048
rect 24202 15952 24258 16008
rect 21074 13388 21130 13424
rect 21074 13368 21076 13388
rect 21076 13368 21128 13388
rect 21128 13368 21130 13388
rect 20890 13232 20946 13288
rect 23817 15258 23873 15260
rect 23897 15258 23953 15260
rect 23977 15258 24033 15260
rect 24057 15258 24113 15260
rect 23817 15206 23843 15258
rect 23843 15206 23873 15258
rect 23897 15206 23907 15258
rect 23907 15206 23953 15258
rect 23977 15206 24023 15258
rect 24023 15206 24033 15258
rect 24057 15206 24087 15258
rect 24087 15206 24113 15258
rect 23817 15204 23873 15206
rect 23897 15204 23953 15206
rect 23977 15204 24033 15206
rect 24057 15204 24113 15206
rect 24938 14864 24994 14920
rect 24846 14764 24848 14784
rect 24848 14764 24900 14784
rect 24900 14764 24902 14784
rect 24846 14728 24902 14764
rect 19150 11450 19206 11452
rect 19230 11450 19286 11452
rect 19310 11450 19366 11452
rect 19390 11450 19446 11452
rect 19150 11398 19176 11450
rect 19176 11398 19206 11450
rect 19230 11398 19240 11450
rect 19240 11398 19286 11450
rect 19310 11398 19356 11450
rect 19356 11398 19366 11450
rect 19390 11398 19420 11450
rect 19420 11398 19446 11450
rect 19150 11396 19206 11398
rect 19230 11396 19286 11398
rect 19310 11396 19366 11398
rect 19390 11396 19446 11398
rect 19694 10668 19750 10704
rect 19694 10648 19696 10668
rect 19696 10648 19748 10668
rect 19748 10648 19750 10668
rect 19150 10362 19206 10364
rect 19230 10362 19286 10364
rect 19310 10362 19366 10364
rect 19390 10362 19446 10364
rect 19150 10310 19176 10362
rect 19176 10310 19206 10362
rect 19230 10310 19240 10362
rect 19240 10310 19286 10362
rect 19310 10310 19356 10362
rect 19356 10310 19366 10362
rect 19390 10310 19420 10362
rect 19420 10310 19446 10362
rect 19150 10308 19206 10310
rect 19230 10308 19286 10310
rect 19310 10308 19366 10310
rect 19390 10308 19446 10310
rect 20614 11228 20616 11248
rect 20616 11228 20668 11248
rect 20668 11228 20670 11248
rect 20614 11192 20670 11228
rect 23817 14170 23873 14172
rect 23897 14170 23953 14172
rect 23977 14170 24033 14172
rect 24057 14170 24113 14172
rect 23817 14118 23843 14170
rect 23843 14118 23873 14170
rect 23897 14118 23907 14170
rect 23907 14118 23953 14170
rect 23977 14118 24023 14170
rect 24023 14118 24033 14170
rect 24057 14118 24087 14170
rect 24087 14118 24113 14170
rect 23817 14116 23873 14118
rect 23897 14116 23953 14118
rect 23977 14116 24033 14118
rect 24057 14116 24113 14118
rect 23817 13082 23873 13084
rect 23897 13082 23953 13084
rect 23977 13082 24033 13084
rect 24057 13082 24113 13084
rect 23817 13030 23843 13082
rect 23843 13030 23873 13082
rect 23897 13030 23907 13082
rect 23907 13030 23953 13082
rect 23977 13030 24023 13082
rect 24023 13030 24033 13082
rect 24057 13030 24087 13082
rect 24087 13030 24113 13082
rect 23817 13028 23873 13030
rect 23897 13028 23953 13030
rect 23977 13028 24033 13030
rect 24057 13028 24113 13030
rect 24846 12824 24902 12880
rect 23190 12008 23246 12064
rect 17946 9696 18002 9752
rect 16106 8200 16162 8256
rect 17118 6976 17174 7032
rect 18406 9016 18462 9072
rect 19694 9444 19750 9480
rect 19694 9424 19696 9444
rect 19696 9424 19748 9444
rect 19748 9424 19750 9444
rect 19150 9274 19206 9276
rect 19230 9274 19286 9276
rect 19310 9274 19366 9276
rect 19390 9274 19446 9276
rect 19150 9222 19176 9274
rect 19176 9222 19206 9274
rect 19230 9222 19240 9274
rect 19240 9222 19286 9274
rect 19310 9222 19356 9274
rect 19356 9222 19366 9274
rect 19390 9222 19420 9274
rect 19420 9222 19446 9274
rect 19150 9220 19206 9222
rect 19230 9220 19286 9222
rect 19310 9220 19366 9222
rect 19390 9220 19446 9222
rect 22914 10512 22970 10568
rect 22086 9460 22088 9480
rect 22088 9460 22140 9480
rect 22140 9460 22142 9480
rect 22086 9424 22142 9460
rect 19150 8186 19206 8188
rect 19230 8186 19286 8188
rect 19310 8186 19366 8188
rect 19390 8186 19446 8188
rect 19150 8134 19176 8186
rect 19176 8134 19206 8186
rect 19230 8134 19240 8186
rect 19240 8134 19286 8186
rect 19310 8134 19356 8186
rect 19356 8134 19366 8186
rect 19390 8134 19420 8186
rect 19420 8134 19446 8186
rect 19150 8132 19206 8134
rect 19230 8132 19286 8134
rect 19310 8132 19366 8134
rect 19390 8132 19446 8134
rect 20982 7928 21038 7984
rect 22270 7792 22326 7848
rect 19602 7148 19604 7168
rect 19604 7148 19656 7168
rect 19656 7148 19658 7168
rect 19602 7112 19658 7148
rect 19150 7098 19206 7100
rect 19230 7098 19286 7100
rect 19310 7098 19366 7100
rect 19390 7098 19446 7100
rect 19150 7046 19176 7098
rect 19176 7046 19206 7098
rect 19230 7046 19240 7098
rect 19240 7046 19286 7098
rect 19310 7046 19356 7098
rect 19356 7046 19366 7098
rect 19390 7046 19420 7098
rect 19420 7046 19446 7098
rect 19150 7044 19206 7046
rect 19230 7044 19286 7046
rect 19310 7044 19366 7046
rect 19390 7044 19446 7046
rect 18958 6976 19014 7032
rect 18498 6860 18554 6896
rect 18498 6840 18500 6860
rect 18500 6840 18552 6860
rect 18552 6840 18554 6860
rect 17946 6296 18002 6352
rect 17394 5480 17450 5536
rect 19694 6024 19750 6080
rect 19150 6010 19206 6012
rect 19230 6010 19286 6012
rect 19310 6010 19366 6012
rect 19390 6010 19446 6012
rect 19150 5958 19176 6010
rect 19176 5958 19206 6010
rect 19230 5958 19240 6010
rect 19240 5958 19286 6010
rect 19310 5958 19356 6010
rect 19356 5958 19366 6010
rect 19390 5958 19420 6010
rect 19420 5958 19446 6010
rect 19150 5956 19206 5958
rect 19230 5956 19286 5958
rect 19310 5956 19366 5958
rect 19390 5956 19446 5958
rect 19150 4922 19206 4924
rect 19230 4922 19286 4924
rect 19310 4922 19366 4924
rect 19390 4922 19446 4924
rect 19150 4870 19176 4922
rect 19176 4870 19206 4922
rect 19230 4870 19240 4922
rect 19240 4870 19286 4922
rect 19310 4870 19356 4922
rect 19356 4870 19366 4922
rect 19390 4870 19420 4922
rect 19420 4870 19446 4922
rect 19150 4868 19206 4870
rect 19230 4868 19286 4870
rect 19310 4868 19366 4870
rect 19390 4868 19446 4870
rect 18774 3984 18830 4040
rect 19602 3984 19658 4040
rect 16290 2932 16292 2952
rect 16292 2932 16344 2952
rect 16344 2932 16346 2952
rect 16290 2896 16346 2932
rect 19150 3834 19206 3836
rect 19230 3834 19286 3836
rect 19310 3834 19366 3836
rect 19390 3834 19446 3836
rect 19150 3782 19176 3834
rect 19176 3782 19206 3834
rect 19230 3782 19240 3834
rect 19240 3782 19286 3834
rect 19310 3782 19356 3834
rect 19356 3782 19366 3834
rect 19390 3782 19420 3834
rect 19420 3782 19446 3834
rect 19150 3780 19206 3782
rect 19230 3780 19286 3782
rect 19310 3780 19366 3782
rect 19390 3780 19446 3782
rect 19150 2746 19206 2748
rect 19230 2746 19286 2748
rect 19310 2746 19366 2748
rect 19390 2746 19446 2748
rect 19150 2694 19176 2746
rect 19176 2694 19206 2746
rect 19230 2694 19240 2746
rect 19240 2694 19286 2746
rect 19310 2694 19356 2746
rect 19356 2694 19366 2746
rect 19390 2694 19420 2746
rect 19420 2694 19446 2746
rect 19150 2692 19206 2694
rect 19230 2692 19286 2694
rect 19310 2692 19366 2694
rect 19390 2692 19446 2694
rect 23282 11620 23338 11656
rect 23282 11600 23284 11620
rect 23284 11600 23336 11620
rect 23336 11600 23338 11620
rect 23817 11994 23873 11996
rect 23897 11994 23953 11996
rect 23977 11994 24033 11996
rect 24057 11994 24113 11996
rect 23817 11942 23843 11994
rect 23843 11942 23873 11994
rect 23897 11942 23907 11994
rect 23907 11942 23953 11994
rect 23977 11942 24023 11994
rect 24023 11942 24033 11994
rect 24057 11942 24087 11994
rect 24087 11942 24113 11994
rect 23817 11940 23873 11942
rect 23897 11940 23953 11942
rect 23977 11940 24033 11942
rect 24057 11940 24113 11942
rect 23374 8472 23430 8528
rect 23190 8064 23246 8120
rect 23190 7112 23246 7168
rect 23006 6316 23062 6352
rect 23006 6296 23008 6316
rect 23008 6296 23060 6316
rect 23060 6296 23062 6316
rect 23098 5480 23154 5536
rect 23006 4004 23062 4040
rect 23006 3984 23008 4004
rect 23008 3984 23060 4004
rect 23060 3984 23062 4004
rect 23817 10906 23873 10908
rect 23897 10906 23953 10908
rect 23977 10906 24033 10908
rect 24057 10906 24113 10908
rect 23817 10854 23843 10906
rect 23843 10854 23873 10906
rect 23897 10854 23907 10906
rect 23907 10854 23953 10906
rect 23977 10854 24023 10906
rect 24023 10854 24033 10906
rect 24057 10854 24087 10906
rect 24087 10854 24113 10906
rect 23817 10852 23873 10854
rect 23897 10852 23953 10854
rect 23977 10852 24033 10854
rect 24057 10852 24113 10854
rect 23817 9818 23873 9820
rect 23897 9818 23953 9820
rect 23977 9818 24033 9820
rect 24057 9818 24113 9820
rect 23817 9766 23843 9818
rect 23843 9766 23873 9818
rect 23897 9766 23907 9818
rect 23907 9766 23953 9818
rect 23977 9766 24023 9818
rect 24023 9766 24033 9818
rect 24057 9766 24087 9818
rect 24087 9766 24113 9818
rect 23817 9764 23873 9766
rect 23897 9764 23953 9766
rect 23977 9764 24033 9766
rect 24057 9764 24113 9766
rect 23650 9560 23706 9616
rect 24294 9696 24350 9752
rect 24662 9696 24718 9752
rect 23650 7928 23706 7984
rect 23817 8730 23873 8732
rect 23897 8730 23953 8732
rect 23977 8730 24033 8732
rect 24057 8730 24113 8732
rect 23817 8678 23843 8730
rect 23843 8678 23873 8730
rect 23897 8678 23907 8730
rect 23907 8678 23953 8730
rect 23977 8678 24023 8730
rect 24023 8678 24033 8730
rect 24057 8678 24087 8730
rect 24087 8678 24113 8730
rect 23817 8676 23873 8678
rect 23897 8676 23953 8678
rect 23977 8676 24033 8678
rect 24057 8676 24113 8678
rect 23817 7642 23873 7644
rect 23897 7642 23953 7644
rect 23977 7642 24033 7644
rect 24057 7642 24113 7644
rect 23817 7590 23843 7642
rect 23843 7590 23873 7642
rect 23897 7590 23907 7642
rect 23907 7590 23953 7642
rect 23977 7590 24023 7642
rect 24023 7590 24033 7642
rect 24057 7590 24087 7642
rect 24087 7590 24113 7642
rect 23817 7588 23873 7590
rect 23897 7588 23953 7590
rect 23977 7588 24033 7590
rect 24057 7588 24113 7590
rect 25766 11736 25822 11792
rect 25122 10804 25178 10840
rect 25122 10784 25124 10804
rect 25124 10784 25176 10804
rect 25176 10784 25178 10804
rect 24938 10548 24940 10568
rect 24940 10548 24992 10568
rect 24992 10548 24994 10568
rect 24938 10512 24994 10548
rect 23817 6554 23873 6556
rect 23897 6554 23953 6556
rect 23977 6554 24033 6556
rect 24057 6554 24113 6556
rect 23817 6502 23843 6554
rect 23843 6502 23873 6554
rect 23897 6502 23907 6554
rect 23907 6502 23953 6554
rect 23977 6502 24023 6554
rect 24023 6502 24033 6554
rect 24057 6502 24087 6554
rect 24087 6502 24113 6554
rect 23817 6500 23873 6502
rect 23897 6500 23953 6502
rect 23977 6500 24033 6502
rect 24057 6500 24113 6502
rect 24938 8744 24994 8800
rect 24754 8472 24810 8528
rect 24754 7656 24810 7712
rect 25030 6568 25086 6624
rect 24662 5480 24718 5536
rect 23817 5466 23873 5468
rect 23897 5466 23953 5468
rect 23977 5466 24033 5468
rect 24057 5466 24113 5468
rect 23817 5414 23843 5466
rect 23843 5414 23873 5466
rect 23897 5414 23907 5466
rect 23907 5414 23953 5466
rect 23977 5414 24023 5466
rect 24023 5414 24033 5466
rect 24057 5414 24087 5466
rect 24087 5414 24113 5466
rect 23817 5412 23873 5414
rect 23897 5412 23953 5414
rect 23977 5412 24033 5414
rect 24057 5412 24113 5414
rect 24202 4528 24258 4584
rect 25030 4528 25086 4584
rect 23817 4378 23873 4380
rect 23897 4378 23953 4380
rect 23977 4378 24033 4380
rect 24057 4378 24113 4380
rect 23817 4326 23843 4378
rect 23843 4326 23873 4378
rect 23897 4326 23907 4378
rect 23907 4326 23953 4378
rect 23977 4326 24023 4378
rect 24023 4326 24033 4378
rect 24057 4326 24087 4378
rect 24087 4326 24113 4378
rect 23817 4324 23873 4326
rect 23897 4324 23953 4326
rect 23977 4324 24033 4326
rect 24057 4324 24113 4326
rect 24662 3440 24718 3496
rect 23817 3290 23873 3292
rect 23897 3290 23953 3292
rect 23977 3290 24033 3292
rect 24057 3290 24113 3292
rect 23817 3238 23843 3290
rect 23843 3238 23873 3290
rect 23897 3238 23907 3290
rect 23907 3238 23953 3290
rect 23977 3238 24023 3290
rect 24023 3238 24033 3290
rect 24057 3238 24087 3290
rect 24087 3238 24113 3290
rect 23817 3236 23873 3238
rect 23897 3236 23953 3238
rect 23977 3236 24033 3238
rect 24057 3236 24113 3238
rect 23817 2202 23873 2204
rect 23897 2202 23953 2204
rect 23977 2202 24033 2204
rect 24057 2202 24113 2204
rect 23817 2150 23843 2202
rect 23843 2150 23873 2202
rect 23897 2150 23907 2202
rect 23907 2150 23953 2202
rect 23977 2150 24023 2202
rect 24023 2150 24033 2202
rect 24057 2150 24087 2202
rect 24087 2150 24113 2202
rect 23817 2148 23873 2150
rect 23897 2148 23953 2150
rect 23977 2148 24033 2150
rect 24057 2148 24113 2150
rect 24662 1400 24718 1456
rect 25766 6024 25822 6080
rect 25122 448 25178 504
<< metal3 >>
rect 25393 27434 25459 27437
rect 27048 27434 27528 27464
rect 25393 27432 27528 27434
rect 25393 27376 25398 27432
rect 25454 27376 27528 27432
rect 25393 27374 27528 27376
rect 25393 27371 25459 27374
rect 27048 27344 27528 27374
rect 24289 26346 24355 26349
rect 27048 26346 27528 26376
rect 24289 26344 27528 26346
rect 24289 26288 24294 26344
rect 24350 26288 27528 26344
rect 24289 26286 27528 26288
rect 24289 26283 24355 26286
rect 27048 26256 27528 26286
rect 9805 25600 10125 25601
rect 9805 25536 9813 25600
rect 9877 25536 9893 25600
rect 9957 25536 9973 25600
rect 10037 25536 10053 25600
rect 10117 25536 10125 25600
rect 9805 25535 10125 25536
rect 19138 25600 19458 25601
rect 19138 25536 19146 25600
rect 19210 25536 19226 25600
rect 19290 25536 19306 25600
rect 19370 25536 19386 25600
rect 19450 25536 19458 25600
rect 19138 25535 19458 25536
rect 24565 25394 24631 25397
rect 27048 25394 27528 25424
rect 24565 25392 27528 25394
rect 24565 25336 24570 25392
rect 24626 25336 27528 25392
rect 24565 25334 27528 25336
rect 24565 25331 24631 25334
rect 27048 25304 27528 25334
rect 5138 25056 5458 25057
rect 5138 24992 5146 25056
rect 5210 24992 5226 25056
rect 5290 24992 5306 25056
rect 5370 24992 5386 25056
rect 5450 24992 5458 25056
rect 5138 24991 5458 24992
rect 14472 25056 14792 25057
rect 14472 24992 14480 25056
rect 14544 24992 14560 25056
rect 14624 24992 14640 25056
rect 14704 24992 14720 25056
rect 14784 24992 14792 25056
rect 14472 24991 14792 24992
rect 23805 25056 24125 25057
rect 23805 24992 23813 25056
rect 23877 24992 23893 25056
rect 23957 24992 23973 25056
rect 24037 24992 24053 25056
rect 24117 24992 24125 25056
rect 23805 24991 24125 24992
rect 18493 24850 18559 24853
rect 20701 24850 20767 24853
rect 18493 24848 20767 24850
rect 18493 24792 18498 24848
rect 18554 24792 20706 24848
rect 20762 24792 20767 24848
rect 18493 24790 20767 24792
rect 18493 24787 18559 24790
rect 20701 24787 20767 24790
rect 14445 24714 14511 24717
rect 19597 24714 19663 24717
rect 14445 24712 19663 24714
rect 14445 24656 14450 24712
rect 14506 24656 19602 24712
rect 19658 24656 19663 24712
rect 14445 24654 19663 24656
rect 14445 24651 14511 24654
rect 19597 24651 19663 24654
rect 9805 24512 10125 24513
rect 9805 24448 9813 24512
rect 9877 24448 9893 24512
rect 9957 24448 9973 24512
rect 10037 24448 10053 24512
rect 10117 24448 10125 24512
rect 9805 24447 10125 24448
rect 19138 24512 19458 24513
rect 19138 24448 19146 24512
rect 19210 24448 19226 24512
rect 19290 24448 19306 24512
rect 19370 24448 19386 24512
rect 19450 24448 19458 24512
rect 19138 24447 19458 24448
rect 14997 24442 15063 24445
rect 17573 24442 17639 24445
rect 14997 24440 17639 24442
rect 14997 24384 15002 24440
rect 15058 24384 17578 24440
rect 17634 24384 17639 24440
rect 14997 24382 17639 24384
rect 14997 24379 15063 24382
rect 17573 24379 17639 24382
rect 22265 24442 22331 24445
rect 23737 24442 23803 24445
rect 22265 24440 23803 24442
rect 22265 24384 22270 24440
rect 22326 24384 23742 24440
rect 23798 24384 23803 24440
rect 22265 24382 23803 24384
rect 22265 24379 22331 24382
rect 23737 24379 23803 24382
rect 1 24306 67 24309
rect 8373 24306 8439 24309
rect 1 24304 8439 24306
rect 1 24248 6 24304
rect 62 24248 8378 24304
rect 8434 24248 8439 24304
rect 1 24246 8439 24248
rect 1 24243 67 24246
rect 8373 24243 8439 24246
rect 10949 24306 11015 24309
rect 18585 24306 18651 24309
rect 10949 24304 18651 24306
rect 10949 24248 10954 24304
rect 11010 24248 18590 24304
rect 18646 24248 18651 24304
rect 10949 24246 18651 24248
rect 10949 24243 11015 24246
rect 18585 24243 18651 24246
rect 20609 24306 20675 24309
rect 24473 24306 24539 24309
rect 20609 24304 24539 24306
rect 20609 24248 20614 24304
rect 20670 24248 24478 24304
rect 24534 24248 24539 24304
rect 20609 24246 24539 24248
rect 20609 24243 20675 24246
rect 24473 24243 24539 24246
rect 25301 24306 25367 24309
rect 27048 24306 27528 24336
rect 25301 24304 27528 24306
rect 25301 24248 25306 24304
rect 25362 24248 27528 24304
rect 25301 24246 27528 24248
rect 25301 24243 25367 24246
rect 27048 24216 27528 24246
rect 1933 24170 1999 24173
rect 10857 24170 10923 24173
rect 1933 24168 10923 24170
rect 1933 24112 1938 24168
rect 1994 24112 10862 24168
rect 10918 24112 10923 24168
rect 1933 24110 10923 24112
rect 1933 24107 1999 24110
rect 10857 24107 10923 24110
rect 16561 24170 16627 24173
rect 20793 24170 20859 24173
rect 16561 24168 20859 24170
rect 16561 24112 16566 24168
rect 16622 24112 20798 24168
rect 20854 24112 20859 24168
rect 16561 24110 20859 24112
rect 16561 24107 16627 24110
rect 20793 24107 20859 24110
rect 5138 23968 5458 23969
rect 5138 23904 5146 23968
rect 5210 23904 5226 23968
rect 5290 23904 5306 23968
rect 5370 23904 5386 23968
rect 5450 23904 5458 23968
rect 5138 23903 5458 23904
rect 14472 23968 14792 23969
rect 14472 23904 14480 23968
rect 14544 23904 14560 23968
rect 14624 23904 14640 23968
rect 14704 23904 14720 23968
rect 14784 23904 14792 23968
rect 14472 23903 14792 23904
rect 23805 23968 24125 23969
rect 23805 23904 23813 23968
rect 23877 23904 23893 23968
rect 23957 23904 23973 23968
rect 24037 23904 24053 23968
rect 24117 23904 24125 23968
rect 23805 23903 24125 23904
rect 19689 23898 19755 23901
rect 22725 23898 22791 23901
rect 19689 23896 22791 23898
rect 19689 23840 19694 23896
rect 19750 23840 22730 23896
rect 22786 23840 22791 23896
rect 19689 23838 22791 23840
rect 19689 23835 19755 23838
rect 22725 23835 22791 23838
rect 3589 23626 3655 23629
rect 14077 23626 14143 23629
rect 3589 23624 14143 23626
rect 3589 23568 3594 23624
rect 3650 23568 14082 23624
rect 14138 23568 14143 23624
rect 3589 23566 14143 23568
rect 3589 23563 3655 23566
rect 14077 23563 14143 23566
rect 24289 23490 24355 23493
rect 25853 23490 25919 23493
rect 24289 23488 25919 23490
rect 24289 23432 24294 23488
rect 24350 23432 25858 23488
rect 25914 23432 25919 23488
rect 24289 23430 25919 23432
rect 24289 23427 24355 23430
rect 25853 23427 25919 23430
rect 9805 23424 10125 23425
rect 9805 23360 9813 23424
rect 9877 23360 9893 23424
rect 9957 23360 9973 23424
rect 10037 23360 10053 23424
rect 10117 23360 10125 23424
rect 9805 23359 10125 23360
rect 19138 23424 19458 23425
rect 19138 23360 19146 23424
rect 19210 23360 19226 23424
rect 19290 23360 19306 23424
rect 19370 23360 19386 23424
rect 19450 23360 19458 23424
rect 19138 23359 19458 23360
rect 7729 23218 7795 23221
rect 21437 23218 21503 23221
rect 7729 23216 21503 23218
rect 7729 23160 7734 23216
rect 7790 23160 21442 23216
rect 21498 23160 21503 23216
rect 7729 23158 21503 23160
rect 7729 23155 7795 23158
rect 21437 23155 21503 23158
rect 25301 23218 25367 23221
rect 27048 23218 27528 23248
rect 25301 23216 27528 23218
rect 25301 23160 25306 23216
rect 25362 23160 27528 23216
rect 25301 23158 27528 23160
rect 25301 23155 25367 23158
rect 27048 23128 27528 23158
rect 4969 23082 5035 23085
rect 16653 23082 16719 23085
rect 4969 23080 16719 23082
rect 4969 23024 4974 23080
rect 5030 23024 16658 23080
rect 16714 23024 16719 23080
rect 4969 23022 16719 23024
rect 4969 23019 5035 23022
rect 16653 23019 16719 23022
rect 17665 23082 17731 23085
rect 24473 23082 24539 23085
rect 17665 23080 24539 23082
rect 17665 23024 17670 23080
rect 17726 23024 24478 23080
rect 24534 23024 24539 23080
rect 17665 23022 24539 23024
rect 17665 23019 17731 23022
rect 24473 23019 24539 23022
rect 5138 22880 5458 22881
rect 5138 22816 5146 22880
rect 5210 22816 5226 22880
rect 5290 22816 5306 22880
rect 5370 22816 5386 22880
rect 5450 22816 5458 22880
rect 5138 22815 5458 22816
rect 14472 22880 14792 22881
rect 14472 22816 14480 22880
rect 14544 22816 14560 22880
rect 14624 22816 14640 22880
rect 14704 22816 14720 22880
rect 14784 22816 14792 22880
rect 14472 22815 14792 22816
rect 23805 22880 24125 22881
rect 23805 22816 23813 22880
rect 23877 22816 23893 22880
rect 23957 22816 23973 22880
rect 24037 22816 24053 22880
rect 24117 22816 24125 22880
rect 23805 22815 24125 22816
rect 9805 22336 10125 22337
rect 9805 22272 9813 22336
rect 9877 22272 9893 22336
rect 9957 22272 9973 22336
rect 10037 22272 10053 22336
rect 10117 22272 10125 22336
rect 9805 22271 10125 22272
rect 19138 22336 19458 22337
rect 19138 22272 19146 22336
rect 19210 22272 19226 22336
rect 19290 22272 19306 22336
rect 19370 22272 19386 22336
rect 19450 22272 19458 22336
rect 19138 22271 19458 22272
rect 24473 22266 24539 22269
rect 27048 22266 27528 22296
rect 24473 22264 27528 22266
rect 24473 22208 24478 22264
rect 24534 22208 27528 22264
rect 24473 22206 27528 22208
rect 24473 22203 24539 22206
rect 27048 22176 27528 22206
rect 6257 21994 6323 21997
rect 20517 21994 20583 21997
rect 6257 21992 20583 21994
rect 6257 21936 6262 21992
rect 6318 21936 20522 21992
rect 20578 21936 20583 21992
rect 6257 21934 20583 21936
rect 6257 21931 6323 21934
rect 20517 21931 20583 21934
rect 5138 21792 5458 21793
rect 5138 21728 5146 21792
rect 5210 21728 5226 21792
rect 5290 21728 5306 21792
rect 5370 21728 5386 21792
rect 5450 21728 5458 21792
rect 5138 21727 5458 21728
rect 14472 21792 14792 21793
rect 14472 21728 14480 21792
rect 14544 21728 14560 21792
rect 14624 21728 14640 21792
rect 14704 21728 14720 21792
rect 14784 21728 14792 21792
rect 14472 21727 14792 21728
rect 23805 21792 24125 21793
rect 23805 21728 23813 21792
rect 23877 21728 23893 21792
rect 23957 21728 23973 21792
rect 24037 21728 24053 21792
rect 24117 21728 24125 21792
rect 23805 21727 24125 21728
rect 2209 21586 2275 21589
rect 7453 21586 7519 21589
rect 2209 21584 7519 21586
rect 2209 21528 2214 21584
rect 2270 21528 7458 21584
rect 7514 21528 7519 21584
rect 2209 21526 7519 21528
rect 2209 21523 2275 21526
rect 7453 21523 7519 21526
rect 15917 21586 15983 21589
rect 24381 21586 24447 21589
rect 15917 21584 24447 21586
rect 15917 21528 15922 21584
rect 15978 21528 24386 21584
rect 24442 21528 24447 21584
rect 15917 21526 24447 21528
rect 15917 21523 15983 21526
rect 24381 21523 24447 21526
rect 18585 21450 18651 21453
rect 20425 21450 20491 21453
rect 18585 21448 20491 21450
rect 18585 21392 18590 21448
rect 18646 21392 20430 21448
rect 20486 21392 20491 21448
rect 18585 21390 20491 21392
rect 18585 21387 18651 21390
rect 20425 21387 20491 21390
rect 9805 21248 10125 21249
rect 9805 21184 9813 21248
rect 9877 21184 9893 21248
rect 9957 21184 9973 21248
rect 10037 21184 10053 21248
rect 10117 21184 10125 21248
rect 9805 21183 10125 21184
rect 19138 21248 19458 21249
rect 19138 21184 19146 21248
rect 19210 21184 19226 21248
rect 19290 21184 19306 21248
rect 19370 21184 19386 21248
rect 19450 21184 19458 21248
rect 19138 21183 19458 21184
rect 24289 21178 24355 21181
rect 27048 21178 27528 21208
rect 24289 21176 27528 21178
rect 24289 21120 24294 21176
rect 24350 21120 27528 21176
rect 24289 21118 27528 21120
rect 24289 21115 24355 21118
rect 27048 21088 27528 21118
rect 18493 21042 18559 21045
rect 24473 21042 24539 21045
rect 18493 21040 24539 21042
rect 18493 20984 18498 21040
rect 18554 20984 24478 21040
rect 24534 20984 24539 21040
rect 18493 20982 24539 20984
rect 18493 20979 18559 20982
rect 24473 20979 24539 20982
rect 5138 20704 5458 20705
rect 5138 20640 5146 20704
rect 5210 20640 5226 20704
rect 5290 20640 5306 20704
rect 5370 20640 5386 20704
rect 5450 20640 5458 20704
rect 5138 20639 5458 20640
rect 14472 20704 14792 20705
rect 14472 20640 14480 20704
rect 14544 20640 14560 20704
rect 14624 20640 14640 20704
rect 14704 20640 14720 20704
rect 14784 20640 14792 20704
rect 14472 20639 14792 20640
rect 23805 20704 24125 20705
rect 23805 20640 23813 20704
rect 23877 20640 23893 20704
rect 23957 20640 23973 20704
rect 24037 20640 24053 20704
rect 24117 20640 24125 20704
rect 23805 20639 24125 20640
rect 17665 20634 17731 20637
rect 20517 20634 20583 20637
rect 17665 20632 20583 20634
rect 17665 20576 17670 20632
rect 17726 20576 20522 20632
rect 20578 20576 20583 20632
rect 17665 20574 20583 20576
rect 17665 20571 17731 20574
rect 20517 20571 20583 20574
rect 12697 20362 12763 20365
rect 23001 20362 23067 20365
rect 12697 20360 23067 20362
rect 12697 20304 12702 20360
rect 12758 20304 23006 20360
rect 23062 20304 23067 20360
rect 12697 20302 23067 20304
rect 12697 20299 12763 20302
rect 23001 20299 23067 20302
rect 9805 20160 10125 20161
rect 9805 20096 9813 20160
rect 9877 20096 9893 20160
rect 9957 20096 9973 20160
rect 10037 20096 10053 20160
rect 10117 20096 10125 20160
rect 9805 20095 10125 20096
rect 19138 20160 19458 20161
rect 19138 20096 19146 20160
rect 19210 20096 19226 20160
rect 19290 20096 19306 20160
rect 19370 20096 19386 20160
rect 19450 20096 19458 20160
rect 19138 20095 19458 20096
rect 25393 20090 25459 20093
rect 27048 20090 27528 20120
rect 25393 20088 27528 20090
rect 25393 20032 25398 20088
rect 25454 20032 27528 20088
rect 25393 20030 27528 20032
rect 25393 20027 25459 20030
rect 27048 20000 27528 20030
rect 4969 19954 5035 19957
rect 17665 19954 17731 19957
rect 4969 19952 17731 19954
rect 4969 19896 4974 19952
rect 5030 19896 17670 19952
rect 17726 19896 17731 19952
rect 4969 19894 17731 19896
rect 4969 19891 5035 19894
rect 17665 19891 17731 19894
rect 9017 19818 9083 19821
rect 24381 19818 24447 19821
rect 9017 19816 24447 19818
rect 9017 19760 9022 19816
rect 9078 19760 24386 19816
rect 24442 19760 24447 19816
rect 9017 19758 24447 19760
rect 9017 19755 9083 19758
rect 24381 19755 24447 19758
rect 5138 19616 5458 19617
rect 5138 19552 5146 19616
rect 5210 19552 5226 19616
rect 5290 19552 5306 19616
rect 5370 19552 5386 19616
rect 5450 19552 5458 19616
rect 5138 19551 5458 19552
rect 14472 19616 14792 19617
rect 14472 19552 14480 19616
rect 14544 19552 14560 19616
rect 14624 19552 14640 19616
rect 14704 19552 14720 19616
rect 14784 19552 14792 19616
rect 14472 19551 14792 19552
rect 23805 19616 24125 19617
rect 23805 19552 23813 19616
rect 23877 19552 23893 19616
rect 23957 19552 23973 19616
rect 24037 19552 24053 19616
rect 24117 19552 24125 19616
rect 23805 19551 24125 19552
rect 11501 19274 11567 19277
rect 13157 19274 13223 19277
rect 11501 19272 13223 19274
rect 11501 19216 11506 19272
rect 11562 19216 13162 19272
rect 13218 19216 13223 19272
rect 11501 19214 13223 19216
rect 11501 19211 11567 19214
rect 13157 19211 13223 19214
rect 23737 19138 23803 19141
rect 27048 19138 27528 19168
rect 23737 19136 27528 19138
rect 23737 19080 23742 19136
rect 23798 19080 27528 19136
rect 23737 19078 27528 19080
rect 23737 19075 23803 19078
rect 9805 19072 10125 19073
rect 9805 19008 9813 19072
rect 9877 19008 9893 19072
rect 9957 19008 9973 19072
rect 10037 19008 10053 19072
rect 10117 19008 10125 19072
rect 9805 19007 10125 19008
rect 19138 19072 19458 19073
rect 19138 19008 19146 19072
rect 19210 19008 19226 19072
rect 19290 19008 19306 19072
rect 19370 19008 19386 19072
rect 19450 19008 19458 19072
rect 27048 19048 27528 19078
rect 19138 19007 19458 19008
rect 9201 18730 9267 18733
rect 9477 18730 9543 18733
rect 11961 18730 12027 18733
rect 9201 18728 12027 18730
rect 9201 18672 9206 18728
rect 9262 18672 9482 18728
rect 9538 18672 11966 18728
rect 12022 18672 12027 18728
rect 9201 18670 12027 18672
rect 9201 18667 9267 18670
rect 9477 18667 9543 18670
rect 11961 18667 12027 18670
rect 9569 18594 9635 18597
rect 13801 18594 13867 18597
rect 9569 18592 13867 18594
rect 9569 18536 9574 18592
rect 9630 18536 13806 18592
rect 13862 18536 13867 18592
rect 9569 18534 13867 18536
rect 9569 18531 9635 18534
rect 13801 18531 13867 18534
rect 5138 18528 5458 18529
rect 5138 18464 5146 18528
rect 5210 18464 5226 18528
rect 5290 18464 5306 18528
rect 5370 18464 5386 18528
rect 5450 18464 5458 18528
rect 5138 18463 5458 18464
rect 14472 18528 14792 18529
rect 14472 18464 14480 18528
rect 14544 18464 14560 18528
rect 14624 18464 14640 18528
rect 14704 18464 14720 18528
rect 14784 18464 14792 18528
rect 14472 18463 14792 18464
rect 23805 18528 24125 18529
rect 23805 18464 23813 18528
rect 23877 18464 23893 18528
rect 23957 18464 23973 18528
rect 24037 18464 24053 18528
rect 24117 18464 24125 18528
rect 23805 18463 24125 18464
rect 23921 18050 23987 18053
rect 24473 18050 24539 18053
rect 23921 18048 24539 18050
rect 23921 17992 23926 18048
rect 23982 17992 24478 18048
rect 24534 17992 24539 18048
rect 23921 17990 24539 17992
rect 23921 17987 23987 17990
rect 24473 17987 24539 17990
rect 25485 18050 25551 18053
rect 27048 18050 27528 18080
rect 25485 18048 27528 18050
rect 25485 17992 25490 18048
rect 25546 17992 27528 18048
rect 25485 17990 27528 17992
rect 25485 17987 25551 17990
rect 9805 17984 10125 17985
rect 9805 17920 9813 17984
rect 9877 17920 9893 17984
rect 9957 17920 9973 17984
rect 10037 17920 10053 17984
rect 10117 17920 10125 17984
rect 9805 17919 10125 17920
rect 19138 17984 19458 17985
rect 19138 17920 19146 17984
rect 19210 17920 19226 17984
rect 19290 17920 19306 17984
rect 19370 17920 19386 17984
rect 19450 17920 19458 17984
rect 27048 17960 27528 17990
rect 19138 17919 19458 17920
rect 15917 17506 15983 17509
rect 20149 17506 20215 17509
rect 15917 17504 20215 17506
rect 15917 17448 15922 17504
rect 15978 17448 20154 17504
rect 20210 17448 20215 17504
rect 15917 17446 20215 17448
rect 15917 17443 15983 17446
rect 20149 17443 20215 17446
rect 5138 17440 5458 17441
rect 5138 17376 5146 17440
rect 5210 17376 5226 17440
rect 5290 17376 5306 17440
rect 5370 17376 5386 17440
rect 5450 17376 5458 17440
rect 5138 17375 5458 17376
rect 14472 17440 14792 17441
rect 14472 17376 14480 17440
rect 14544 17376 14560 17440
rect 14624 17376 14640 17440
rect 14704 17376 14720 17440
rect 14784 17376 14792 17440
rect 14472 17375 14792 17376
rect 23805 17440 24125 17441
rect 23805 17376 23813 17440
rect 23877 17376 23893 17440
rect 23957 17376 23973 17440
rect 24037 17376 24053 17440
rect 24117 17376 24125 17440
rect 23805 17375 24125 17376
rect 14629 17234 14695 17237
rect 16193 17234 16259 17237
rect 14629 17232 16259 17234
rect 14629 17176 14634 17232
rect 14690 17176 16198 17232
rect 16254 17176 16259 17232
rect 14629 17174 16259 17176
rect 14629 17171 14695 17174
rect 16193 17171 16259 17174
rect 24933 17098 24999 17101
rect 27048 17098 27528 17128
rect 24933 17096 27528 17098
rect 24933 17040 24938 17096
rect 24994 17040 27528 17096
rect 24933 17038 27528 17040
rect 24933 17035 24999 17038
rect 27048 17008 27528 17038
rect 9805 16896 10125 16897
rect 9805 16832 9813 16896
rect 9877 16832 9893 16896
rect 9957 16832 9973 16896
rect 10037 16832 10053 16896
rect 10117 16832 10125 16896
rect 9805 16831 10125 16832
rect 19138 16896 19458 16897
rect 19138 16832 19146 16896
rect 19210 16832 19226 16896
rect 19290 16832 19306 16896
rect 19370 16832 19386 16896
rect 19450 16832 19458 16896
rect 19138 16831 19458 16832
rect 10397 16690 10463 16693
rect 10765 16690 10831 16693
rect 13801 16690 13867 16693
rect 10397 16688 13867 16690
rect 10397 16632 10402 16688
rect 10458 16632 10770 16688
rect 10826 16632 13806 16688
rect 13862 16632 13867 16688
rect 10397 16630 13867 16632
rect 10397 16627 10463 16630
rect 10765 16627 10831 16630
rect 13801 16627 13867 16630
rect 20149 16690 20215 16693
rect 23185 16690 23251 16693
rect 20149 16688 23251 16690
rect 20149 16632 20154 16688
rect 20210 16632 23190 16688
rect 23246 16632 23251 16688
rect 20149 16630 23251 16632
rect 20149 16627 20215 16630
rect 23185 16627 23251 16630
rect 13157 16554 13223 16557
rect 14905 16554 14971 16557
rect 13157 16552 14971 16554
rect 13157 16496 13162 16552
rect 13218 16496 14910 16552
rect 14966 16496 14971 16552
rect 13157 16494 14971 16496
rect 13157 16491 13223 16494
rect 14905 16491 14971 16494
rect 5138 16352 5458 16353
rect 5138 16288 5146 16352
rect 5210 16288 5226 16352
rect 5290 16288 5306 16352
rect 5370 16288 5386 16352
rect 5450 16288 5458 16352
rect 5138 16287 5458 16288
rect 14472 16352 14792 16353
rect 14472 16288 14480 16352
rect 14544 16288 14560 16352
rect 14624 16288 14640 16352
rect 14704 16288 14720 16352
rect 14784 16288 14792 16352
rect 14472 16287 14792 16288
rect 23805 16352 24125 16353
rect 23805 16288 23813 16352
rect 23877 16288 23893 16352
rect 23957 16288 23973 16352
rect 24037 16288 24053 16352
rect 24117 16288 24125 16352
rect 23805 16287 24125 16288
rect 10581 16146 10647 16149
rect 23001 16146 23067 16149
rect 10581 16144 23067 16146
rect 10581 16088 10586 16144
rect 10642 16088 23006 16144
rect 23062 16088 23067 16144
rect 10581 16086 23067 16088
rect 10581 16083 10647 16086
rect 23001 16083 23067 16086
rect 24197 16010 24263 16013
rect 27048 16010 27528 16040
rect 24197 16008 27528 16010
rect 24197 15952 24202 16008
rect 24258 15952 27528 16008
rect 24197 15950 27528 15952
rect 24197 15947 24263 15950
rect 27048 15920 27528 15950
rect 10213 15874 10279 15877
rect 10581 15874 10647 15877
rect 17297 15874 17363 15877
rect 10213 15872 17363 15874
rect 10213 15816 10218 15872
rect 10274 15816 10586 15872
rect 10642 15816 17302 15872
rect 17358 15816 17363 15872
rect 10213 15814 17363 15816
rect 10213 15811 10279 15814
rect 10581 15811 10647 15814
rect 17297 15811 17363 15814
rect 9805 15808 10125 15809
rect 9805 15744 9813 15808
rect 9877 15744 9893 15808
rect 9957 15744 9973 15808
rect 10037 15744 10053 15808
rect 10117 15744 10125 15808
rect 9805 15743 10125 15744
rect 19138 15808 19458 15809
rect 19138 15744 19146 15808
rect 19210 15744 19226 15808
rect 19290 15744 19306 15808
rect 19370 15744 19386 15808
rect 19450 15744 19458 15808
rect 19138 15743 19458 15744
rect 14169 15738 14235 15741
rect 17665 15738 17731 15741
rect 18217 15738 18283 15741
rect 14169 15736 18283 15738
rect 14169 15680 14174 15736
rect 14230 15680 17670 15736
rect 17726 15680 18222 15736
rect 18278 15680 18283 15736
rect 14169 15678 18283 15680
rect 14169 15675 14235 15678
rect 17665 15675 17731 15678
rect 18217 15675 18283 15678
rect 5138 15264 5458 15265
rect 5138 15200 5146 15264
rect 5210 15200 5226 15264
rect 5290 15200 5306 15264
rect 5370 15200 5386 15264
rect 5450 15200 5458 15264
rect 5138 15199 5458 15200
rect 14472 15264 14792 15265
rect 14472 15200 14480 15264
rect 14544 15200 14560 15264
rect 14624 15200 14640 15264
rect 14704 15200 14720 15264
rect 14784 15200 14792 15264
rect 14472 15199 14792 15200
rect 23805 15264 24125 15265
rect 23805 15200 23813 15264
rect 23877 15200 23893 15264
rect 23957 15200 23973 15264
rect 24037 15200 24053 15264
rect 24117 15200 24125 15264
rect 23805 15199 24125 15200
rect 24933 14922 24999 14925
rect 27048 14922 27528 14952
rect 24933 14920 27528 14922
rect 24933 14864 24938 14920
rect 24994 14864 27528 14920
rect 24933 14862 27528 14864
rect 24933 14859 24999 14862
rect 27048 14832 27528 14862
rect 20701 14786 20767 14789
rect 24841 14786 24907 14789
rect 20701 14784 24907 14786
rect 20701 14728 20706 14784
rect 20762 14728 24846 14784
rect 24902 14728 24907 14784
rect 20701 14726 24907 14728
rect 20701 14723 20767 14726
rect 24841 14723 24907 14726
rect 9805 14720 10125 14721
rect 9805 14656 9813 14720
rect 9877 14656 9893 14720
rect 9957 14656 9973 14720
rect 10037 14656 10053 14720
rect 10117 14656 10125 14720
rect 9805 14655 10125 14656
rect 19138 14720 19458 14721
rect 19138 14656 19146 14720
rect 19210 14656 19226 14720
rect 19290 14656 19306 14720
rect 19370 14656 19386 14720
rect 19450 14656 19458 14720
rect 19138 14655 19458 14656
rect 5138 14176 5458 14177
rect 5138 14112 5146 14176
rect 5210 14112 5226 14176
rect 5290 14112 5306 14176
rect 5370 14112 5386 14176
rect 5450 14112 5458 14176
rect 5138 14111 5458 14112
rect 14472 14176 14792 14177
rect 14472 14112 14480 14176
rect 14544 14112 14560 14176
rect 14624 14112 14640 14176
rect 14704 14112 14720 14176
rect 14784 14112 14792 14176
rect 14472 14111 14792 14112
rect 23805 14176 24125 14177
rect 23805 14112 23813 14176
rect 23877 14112 23893 14176
rect 23957 14112 23973 14176
rect 24037 14112 24053 14176
rect 24117 14112 24125 14176
rect 23805 14111 24125 14112
rect 24238 13908 24244 13972
rect 24308 13970 24314 13972
rect 27048 13970 27528 14000
rect 24308 13910 27528 13970
rect 24308 13908 24314 13910
rect 27048 13880 27528 13910
rect 15917 13834 15983 13837
rect 18125 13834 18191 13837
rect 15917 13832 18191 13834
rect 15917 13776 15922 13832
rect 15978 13776 18130 13832
rect 18186 13776 18191 13832
rect 15917 13774 18191 13776
rect 15917 13771 15983 13774
rect 18125 13771 18191 13774
rect 9805 13632 10125 13633
rect 9805 13568 9813 13632
rect 9877 13568 9893 13632
rect 9957 13568 9973 13632
rect 10037 13568 10053 13632
rect 10117 13568 10125 13632
rect 9805 13567 10125 13568
rect 19138 13632 19458 13633
rect 19138 13568 19146 13632
rect 19210 13568 19226 13632
rect 19290 13568 19306 13632
rect 19370 13568 19386 13632
rect 19450 13568 19458 13632
rect 19138 13567 19458 13568
rect 13893 13426 13959 13429
rect 21069 13426 21135 13429
rect 13893 13424 21135 13426
rect 13893 13368 13898 13424
rect 13954 13368 21074 13424
rect 21130 13368 21135 13424
rect 13893 13366 21135 13368
rect 13893 13363 13959 13366
rect 21069 13363 21135 13366
rect 14353 13290 14419 13293
rect 20885 13290 20951 13293
rect 14353 13288 20951 13290
rect 14353 13232 14358 13288
rect 14414 13232 20890 13288
rect 20946 13232 20951 13288
rect 14353 13230 20951 13232
rect 14353 13227 14419 13230
rect 20885 13227 20951 13230
rect 5138 13088 5458 13089
rect 5138 13024 5146 13088
rect 5210 13024 5226 13088
rect 5290 13024 5306 13088
rect 5370 13024 5386 13088
rect 5450 13024 5458 13088
rect 5138 13023 5458 13024
rect 14472 13088 14792 13089
rect 14472 13024 14480 13088
rect 14544 13024 14560 13088
rect 14624 13024 14640 13088
rect 14704 13024 14720 13088
rect 14784 13024 14792 13088
rect 14472 13023 14792 13024
rect 23805 13088 24125 13089
rect 23805 13024 23813 13088
rect 23877 13024 23893 13088
rect 23957 13024 23973 13088
rect 24037 13024 24053 13088
rect 24117 13024 24125 13088
rect 23805 13023 24125 13024
rect 24841 12882 24907 12885
rect 27048 12882 27528 12912
rect 24841 12880 27528 12882
rect 24841 12824 24846 12880
rect 24902 12824 27528 12880
rect 24841 12822 27528 12824
rect 24841 12819 24907 12822
rect 27048 12792 27528 12822
rect 9805 12544 10125 12545
rect 9805 12480 9813 12544
rect 9877 12480 9893 12544
rect 9957 12480 9973 12544
rect 10037 12480 10053 12544
rect 10117 12480 10125 12544
rect 9805 12479 10125 12480
rect 19138 12544 19458 12545
rect 19138 12480 19146 12544
rect 19210 12480 19226 12544
rect 19290 12480 19306 12544
rect 19370 12480 19386 12544
rect 19450 12480 19458 12544
rect 19138 12479 19458 12480
rect 18769 12066 18835 12069
rect 23185 12066 23251 12069
rect 18769 12064 23251 12066
rect 18769 12008 18774 12064
rect 18830 12008 23190 12064
rect 23246 12008 23251 12064
rect 18769 12006 23251 12008
rect 18769 12003 18835 12006
rect 23185 12003 23251 12006
rect 5138 12000 5458 12001
rect 5138 11936 5146 12000
rect 5210 11936 5226 12000
rect 5290 11936 5306 12000
rect 5370 11936 5386 12000
rect 5450 11936 5458 12000
rect 5138 11935 5458 11936
rect 14472 12000 14792 12001
rect 14472 11936 14480 12000
rect 14544 11936 14560 12000
rect 14624 11936 14640 12000
rect 14704 11936 14720 12000
rect 14784 11936 14792 12000
rect 14472 11935 14792 11936
rect 23805 12000 24125 12001
rect 23805 11936 23813 12000
rect 23877 11936 23893 12000
rect 23957 11936 23973 12000
rect 24037 11936 24053 12000
rect 24117 11936 24125 12000
rect 23805 11935 24125 11936
rect 25761 11794 25827 11797
rect 27048 11794 27528 11824
rect 25761 11792 27528 11794
rect 25761 11736 25766 11792
rect 25822 11736 27528 11792
rect 25761 11734 27528 11736
rect 25761 11731 25827 11734
rect 27048 11704 27528 11734
rect 9385 11658 9451 11661
rect 23277 11658 23343 11661
rect 9385 11656 23343 11658
rect 9385 11600 9390 11656
rect 9446 11600 23282 11656
rect 23338 11600 23343 11656
rect 9385 11598 23343 11600
rect 9385 11595 9451 11598
rect 23277 11595 23343 11598
rect 10581 11522 10647 11525
rect 13709 11522 13775 11525
rect 10581 11520 13775 11522
rect 10581 11464 10586 11520
rect 10642 11464 13714 11520
rect 13770 11464 13775 11520
rect 10581 11462 13775 11464
rect 10581 11459 10647 11462
rect 13709 11459 13775 11462
rect 9805 11456 10125 11457
rect 9805 11392 9813 11456
rect 9877 11392 9893 11456
rect 9957 11392 9973 11456
rect 10037 11392 10053 11456
rect 10117 11392 10125 11456
rect 9805 11391 10125 11392
rect 19138 11456 19458 11457
rect 19138 11392 19146 11456
rect 19210 11392 19226 11456
rect 19290 11392 19306 11456
rect 19370 11392 19386 11456
rect 19450 11392 19458 11456
rect 19138 11391 19458 11392
rect 16193 11250 16259 11253
rect 20609 11250 20675 11253
rect 16193 11248 20675 11250
rect 16193 11192 16198 11248
rect 16254 11192 20614 11248
rect 20670 11192 20675 11248
rect 16193 11190 20675 11192
rect 16193 11187 16259 11190
rect 20609 11187 20675 11190
rect 10581 11114 10647 11117
rect 10765 11114 10831 11117
rect 10581 11112 10831 11114
rect 10581 11056 10586 11112
rect 10642 11056 10770 11112
rect 10826 11056 10831 11112
rect 10581 11054 10831 11056
rect 10581 11051 10647 11054
rect 10765 11051 10831 11054
rect 5138 10912 5458 10913
rect 5138 10848 5146 10912
rect 5210 10848 5226 10912
rect 5290 10848 5306 10912
rect 5370 10848 5386 10912
rect 5450 10848 5458 10912
rect 5138 10847 5458 10848
rect 14472 10912 14792 10913
rect 14472 10848 14480 10912
rect 14544 10848 14560 10912
rect 14624 10848 14640 10912
rect 14704 10848 14720 10912
rect 14784 10848 14792 10912
rect 14472 10847 14792 10848
rect 23805 10912 24125 10913
rect 23805 10848 23813 10912
rect 23877 10848 23893 10912
rect 23957 10848 23973 10912
rect 24037 10848 24053 10912
rect 24117 10848 24125 10912
rect 23805 10847 24125 10848
rect 25117 10842 25183 10845
rect 27048 10842 27528 10872
rect 25117 10840 27528 10842
rect 25117 10784 25122 10840
rect 25178 10784 27528 10840
rect 25117 10782 27528 10784
rect 25117 10779 25183 10782
rect 27048 10752 27528 10782
rect 14353 10706 14419 10709
rect 19689 10706 19755 10709
rect 14353 10704 19755 10706
rect 14353 10648 14358 10704
rect 14414 10648 19694 10704
rect 19750 10648 19755 10704
rect 14353 10646 19755 10648
rect 14353 10643 14419 10646
rect 19689 10643 19755 10646
rect 22909 10570 22975 10573
rect 24933 10570 24999 10573
rect 22909 10568 24999 10570
rect 22909 10512 22914 10568
rect 22970 10512 24938 10568
rect 24994 10512 24999 10568
rect 22909 10510 24999 10512
rect 22909 10507 22975 10510
rect 24933 10507 24999 10510
rect 9805 10368 10125 10369
rect 9805 10304 9813 10368
rect 9877 10304 9893 10368
rect 9957 10304 9973 10368
rect 10037 10304 10053 10368
rect 10117 10304 10125 10368
rect 9805 10303 10125 10304
rect 19138 10368 19458 10369
rect 19138 10304 19146 10368
rect 19210 10304 19226 10368
rect 19290 10304 19306 10368
rect 19370 10304 19386 10368
rect 19450 10304 19458 10368
rect 19138 10303 19458 10304
rect 5138 9824 5458 9825
rect 5138 9760 5146 9824
rect 5210 9760 5226 9824
rect 5290 9760 5306 9824
rect 5370 9760 5386 9824
rect 5450 9760 5458 9824
rect 5138 9759 5458 9760
rect 14472 9824 14792 9825
rect 14472 9760 14480 9824
rect 14544 9760 14560 9824
rect 14624 9760 14640 9824
rect 14704 9760 14720 9824
rect 14784 9760 14792 9824
rect 14472 9759 14792 9760
rect 23805 9824 24125 9825
rect 23805 9760 23813 9824
rect 23877 9760 23893 9824
rect 23957 9760 23973 9824
rect 24037 9760 24053 9824
rect 24117 9760 24125 9824
rect 23805 9759 24125 9760
rect 17941 9754 18007 9757
rect 24289 9756 24355 9757
rect 24238 9754 24244 9756
rect 17941 9752 23570 9754
rect 17941 9696 17946 9752
rect 18002 9696 23570 9752
rect 17941 9694 23570 9696
rect 24198 9694 24244 9754
rect 24308 9752 24355 9756
rect 24350 9696 24355 9752
rect 17941 9691 18007 9694
rect 23510 9618 23570 9694
rect 24238 9692 24244 9694
rect 24308 9692 24355 9696
rect 24289 9691 24355 9692
rect 24657 9754 24723 9757
rect 27048 9754 27528 9784
rect 24657 9752 27528 9754
rect 24657 9696 24662 9752
rect 24718 9696 27528 9752
rect 24657 9694 27528 9696
rect 24657 9691 24723 9694
rect 27048 9664 27528 9694
rect 23645 9618 23711 9621
rect 23510 9616 23711 9618
rect 23510 9560 23650 9616
rect 23706 9560 23711 9616
rect 23510 9558 23711 9560
rect 23645 9555 23711 9558
rect 19689 9482 19755 9485
rect 22081 9482 22147 9485
rect 19689 9480 22147 9482
rect 19689 9424 19694 9480
rect 19750 9424 22086 9480
rect 22142 9424 22147 9480
rect 19689 9422 22147 9424
rect 19689 9419 19755 9422
rect 22081 9419 22147 9422
rect 9805 9280 10125 9281
rect 9805 9216 9813 9280
rect 9877 9216 9893 9280
rect 9957 9216 9973 9280
rect 10037 9216 10053 9280
rect 10117 9216 10125 9280
rect 9805 9215 10125 9216
rect 19138 9280 19458 9281
rect 19138 9216 19146 9280
rect 19210 9216 19226 9280
rect 19290 9216 19306 9280
rect 19370 9216 19386 9280
rect 19450 9216 19458 9280
rect 19138 9215 19458 9216
rect 12237 9074 12303 9077
rect 18401 9074 18467 9077
rect 12237 9072 18467 9074
rect 12237 9016 12242 9072
rect 12298 9016 18406 9072
rect 18462 9016 18467 9072
rect 12237 9014 18467 9016
rect 12237 9011 12303 9014
rect 18401 9011 18467 9014
rect 24933 8802 24999 8805
rect 27048 8802 27528 8832
rect 24933 8800 27528 8802
rect 24933 8744 24938 8800
rect 24994 8744 27528 8800
rect 24933 8742 27528 8744
rect 24933 8739 24999 8742
rect 5138 8736 5458 8737
rect 5138 8672 5146 8736
rect 5210 8672 5226 8736
rect 5290 8672 5306 8736
rect 5370 8672 5386 8736
rect 5450 8672 5458 8736
rect 5138 8671 5458 8672
rect 14472 8736 14792 8737
rect 14472 8672 14480 8736
rect 14544 8672 14560 8736
rect 14624 8672 14640 8736
rect 14704 8672 14720 8736
rect 14784 8672 14792 8736
rect 14472 8671 14792 8672
rect 23805 8736 24125 8737
rect 23805 8672 23813 8736
rect 23877 8672 23893 8736
rect 23957 8672 23973 8736
rect 24037 8672 24053 8736
rect 24117 8672 24125 8736
rect 27048 8712 27528 8742
rect 23805 8671 24125 8672
rect 23369 8530 23435 8533
rect 24749 8530 24815 8533
rect 23369 8528 24815 8530
rect 23369 8472 23374 8528
rect 23430 8472 24754 8528
rect 24810 8472 24815 8528
rect 23369 8470 24815 8472
rect 23369 8467 23435 8470
rect 24749 8467 24815 8470
rect 13433 8258 13499 8261
rect 14905 8258 14971 8261
rect 16101 8258 16167 8261
rect 13433 8256 16167 8258
rect 13433 8200 13438 8256
rect 13494 8200 14910 8256
rect 14966 8200 16106 8256
rect 16162 8200 16167 8256
rect 13433 8198 16167 8200
rect 13433 8195 13499 8198
rect 14905 8195 14971 8198
rect 16101 8195 16167 8198
rect 9805 8192 10125 8193
rect 9805 8128 9813 8192
rect 9877 8128 9893 8192
rect 9957 8128 9973 8192
rect 10037 8128 10053 8192
rect 10117 8128 10125 8192
rect 9805 8127 10125 8128
rect 19138 8192 19458 8193
rect 19138 8128 19146 8192
rect 19210 8128 19226 8192
rect 19290 8128 19306 8192
rect 19370 8128 19386 8192
rect 19450 8128 19458 8192
rect 19138 8127 19458 8128
rect 23185 8122 23251 8125
rect 23185 8120 23386 8122
rect 23185 8064 23190 8120
rect 23246 8064 23386 8120
rect 23185 8062 23386 8064
rect 23185 8059 23251 8062
rect 8189 7986 8255 7989
rect 20977 7986 21043 7989
rect 8189 7984 21043 7986
rect 8189 7928 8194 7984
rect 8250 7928 20982 7984
rect 21038 7928 21043 7984
rect 8189 7926 21043 7928
rect 23326 7986 23386 8062
rect 23645 7986 23711 7989
rect 23326 7984 23711 7986
rect 23326 7928 23650 7984
rect 23706 7928 23711 7984
rect 23326 7926 23711 7928
rect 8189 7923 8255 7926
rect 20977 7923 21043 7926
rect 23645 7923 23711 7926
rect 14353 7850 14419 7853
rect 22265 7850 22331 7853
rect 14353 7848 22331 7850
rect 14353 7792 14358 7848
rect 14414 7792 22270 7848
rect 22326 7792 22331 7848
rect 14353 7790 22331 7792
rect 14353 7787 14419 7790
rect 22265 7787 22331 7790
rect 24749 7714 24815 7717
rect 27048 7714 27528 7744
rect 24749 7712 27528 7714
rect 24749 7656 24754 7712
rect 24810 7656 27528 7712
rect 24749 7654 27528 7656
rect 24749 7651 24815 7654
rect 5138 7648 5458 7649
rect 5138 7584 5146 7648
rect 5210 7584 5226 7648
rect 5290 7584 5306 7648
rect 5370 7584 5386 7648
rect 5450 7584 5458 7648
rect 5138 7583 5458 7584
rect 14472 7648 14792 7649
rect 14472 7584 14480 7648
rect 14544 7584 14560 7648
rect 14624 7584 14640 7648
rect 14704 7584 14720 7648
rect 14784 7584 14792 7648
rect 14472 7583 14792 7584
rect 23805 7648 24125 7649
rect 23805 7584 23813 7648
rect 23877 7584 23893 7648
rect 23957 7584 23973 7648
rect 24037 7584 24053 7648
rect 24117 7584 24125 7648
rect 27048 7624 27528 7654
rect 23805 7583 24125 7584
rect 11777 7170 11843 7173
rect 13617 7170 13683 7173
rect 11777 7168 13683 7170
rect 11777 7112 11782 7168
rect 11838 7112 13622 7168
rect 13678 7112 13683 7168
rect 11777 7110 13683 7112
rect 11777 7107 11843 7110
rect 13617 7107 13683 7110
rect 19597 7170 19663 7173
rect 23185 7170 23251 7173
rect 19597 7168 23251 7170
rect 19597 7112 19602 7168
rect 19658 7112 23190 7168
rect 23246 7112 23251 7168
rect 19597 7110 23251 7112
rect 19597 7107 19663 7110
rect 23185 7107 23251 7110
rect 9805 7104 10125 7105
rect 9805 7040 9813 7104
rect 9877 7040 9893 7104
rect 9957 7040 9973 7104
rect 10037 7040 10053 7104
rect 10117 7040 10125 7104
rect 9805 7039 10125 7040
rect 19138 7104 19458 7105
rect 19138 7040 19146 7104
rect 19210 7040 19226 7104
rect 19290 7040 19306 7104
rect 19370 7040 19386 7104
rect 19450 7040 19458 7104
rect 19138 7039 19458 7040
rect 17113 7034 17179 7037
rect 18953 7034 19019 7037
rect 17113 7032 19019 7034
rect 17113 6976 17118 7032
rect 17174 6976 18958 7032
rect 19014 6976 19019 7032
rect 17113 6974 19019 6976
rect 17113 6971 17179 6974
rect 18953 6971 19019 6974
rect 11041 6898 11107 6901
rect 18493 6898 18559 6901
rect 11041 6896 18559 6898
rect 11041 6840 11046 6896
rect 11102 6840 18498 6896
rect 18554 6840 18559 6896
rect 11041 6838 18559 6840
rect 11041 6835 11107 6838
rect 18493 6835 18559 6838
rect 25025 6626 25091 6629
rect 27048 6626 27528 6656
rect 25025 6624 27528 6626
rect 25025 6568 25030 6624
rect 25086 6568 27528 6624
rect 25025 6566 27528 6568
rect 25025 6563 25091 6566
rect 5138 6560 5458 6561
rect 5138 6496 5146 6560
rect 5210 6496 5226 6560
rect 5290 6496 5306 6560
rect 5370 6496 5386 6560
rect 5450 6496 5458 6560
rect 5138 6495 5458 6496
rect 14472 6560 14792 6561
rect 14472 6496 14480 6560
rect 14544 6496 14560 6560
rect 14624 6496 14640 6560
rect 14704 6496 14720 6560
rect 14784 6496 14792 6560
rect 14472 6495 14792 6496
rect 23805 6560 24125 6561
rect 23805 6496 23813 6560
rect 23877 6496 23893 6560
rect 23957 6496 23973 6560
rect 24037 6496 24053 6560
rect 24117 6496 24125 6560
rect 27048 6536 27528 6566
rect 23805 6495 24125 6496
rect 17941 6354 18007 6357
rect 23001 6354 23067 6357
rect 17941 6352 23067 6354
rect 17941 6296 17946 6352
rect 18002 6296 23006 6352
rect 23062 6296 23067 6352
rect 17941 6294 23067 6296
rect 17941 6291 18007 6294
rect 23001 6291 23067 6294
rect 19689 6082 19755 6085
rect 25761 6082 25827 6085
rect 19689 6080 25827 6082
rect 19689 6024 19694 6080
rect 19750 6024 25766 6080
rect 25822 6024 25827 6080
rect 19689 6022 25827 6024
rect 19689 6019 19755 6022
rect 25761 6019 25827 6022
rect 9805 6016 10125 6017
rect 9805 5952 9813 6016
rect 9877 5952 9893 6016
rect 9957 5952 9973 6016
rect 10037 5952 10053 6016
rect 10117 5952 10125 6016
rect 9805 5951 10125 5952
rect 19138 6016 19458 6017
rect 19138 5952 19146 6016
rect 19210 5952 19226 6016
rect 19290 5952 19306 6016
rect 19370 5952 19386 6016
rect 19450 5952 19458 6016
rect 19138 5951 19458 5952
rect 8281 5810 8347 5813
rect 11593 5810 11659 5813
rect 8281 5808 11659 5810
rect 8281 5752 8286 5808
rect 8342 5752 11598 5808
rect 11654 5752 11659 5808
rect 8281 5750 11659 5752
rect 8281 5747 8347 5750
rect 11593 5747 11659 5750
rect 27048 5674 27528 5704
rect 24798 5614 27528 5674
rect 17389 5538 17455 5541
rect 23093 5538 23159 5541
rect 17389 5536 23159 5538
rect 17389 5480 17394 5536
rect 17450 5480 23098 5536
rect 23154 5480 23159 5536
rect 17389 5478 23159 5480
rect 17389 5475 17455 5478
rect 23093 5475 23159 5478
rect 24657 5538 24723 5541
rect 24798 5538 24858 5614
rect 27048 5584 27528 5614
rect 24657 5536 24858 5538
rect 24657 5480 24662 5536
rect 24718 5480 24858 5536
rect 24657 5478 24858 5480
rect 24657 5475 24723 5478
rect 5138 5472 5458 5473
rect 5138 5408 5146 5472
rect 5210 5408 5226 5472
rect 5290 5408 5306 5472
rect 5370 5408 5386 5472
rect 5450 5408 5458 5472
rect 5138 5407 5458 5408
rect 14472 5472 14792 5473
rect 14472 5408 14480 5472
rect 14544 5408 14560 5472
rect 14624 5408 14640 5472
rect 14704 5408 14720 5472
rect 14784 5408 14792 5472
rect 14472 5407 14792 5408
rect 23805 5472 24125 5473
rect 23805 5408 23813 5472
rect 23877 5408 23893 5472
rect 23957 5408 23973 5472
rect 24037 5408 24053 5472
rect 24117 5408 24125 5472
rect 23805 5407 24125 5408
rect 10305 5402 10371 5405
rect 13985 5402 14051 5405
rect 10305 5400 14051 5402
rect 10305 5344 10310 5400
rect 10366 5344 13990 5400
rect 14046 5344 14051 5400
rect 10305 5342 14051 5344
rect 10305 5339 10371 5342
rect 13985 5339 14051 5342
rect 9805 4928 10125 4929
rect 9805 4864 9813 4928
rect 9877 4864 9893 4928
rect 9957 4864 9973 4928
rect 10037 4864 10053 4928
rect 10117 4864 10125 4928
rect 9805 4863 10125 4864
rect 19138 4928 19458 4929
rect 19138 4864 19146 4928
rect 19210 4864 19226 4928
rect 19290 4864 19306 4928
rect 19370 4864 19386 4928
rect 19450 4864 19458 4928
rect 19138 4863 19458 4864
rect 24197 4586 24263 4589
rect 25025 4586 25091 4589
rect 27048 4586 27528 4616
rect 24197 4584 27528 4586
rect 24197 4528 24202 4584
rect 24258 4528 25030 4584
rect 25086 4528 27528 4584
rect 24197 4526 27528 4528
rect 24197 4523 24263 4526
rect 25025 4523 25091 4526
rect 27048 4496 27528 4526
rect 5138 4384 5458 4385
rect 5138 4320 5146 4384
rect 5210 4320 5226 4384
rect 5290 4320 5306 4384
rect 5370 4320 5386 4384
rect 5450 4320 5458 4384
rect 5138 4319 5458 4320
rect 14472 4384 14792 4385
rect 14472 4320 14480 4384
rect 14544 4320 14560 4384
rect 14624 4320 14640 4384
rect 14704 4320 14720 4384
rect 14784 4320 14792 4384
rect 14472 4319 14792 4320
rect 23805 4384 24125 4385
rect 23805 4320 23813 4384
rect 23877 4320 23893 4384
rect 23957 4320 23973 4384
rect 24037 4320 24053 4384
rect 24117 4320 24125 4384
rect 23805 4319 24125 4320
rect 4785 4042 4851 4045
rect 10765 4042 10831 4045
rect 4785 4040 10831 4042
rect 4785 3984 4790 4040
rect 4846 3984 10770 4040
rect 10826 3984 10831 4040
rect 4785 3982 10831 3984
rect 4785 3979 4851 3982
rect 10765 3979 10831 3982
rect 14261 4042 14327 4045
rect 18769 4042 18835 4045
rect 14261 4040 18835 4042
rect 14261 3984 14266 4040
rect 14322 3984 18774 4040
rect 18830 3984 18835 4040
rect 14261 3982 18835 3984
rect 14261 3979 14327 3982
rect 18769 3979 18835 3982
rect 19597 4042 19663 4045
rect 23001 4042 23067 4045
rect 19597 4040 23067 4042
rect 19597 3984 19602 4040
rect 19658 3984 23006 4040
rect 23062 3984 23067 4040
rect 19597 3982 23067 3984
rect 19597 3979 19663 3982
rect 23001 3979 23067 3982
rect 9805 3840 10125 3841
rect 9805 3776 9813 3840
rect 9877 3776 9893 3840
rect 9957 3776 9973 3840
rect 10037 3776 10053 3840
rect 10117 3776 10125 3840
rect 9805 3775 10125 3776
rect 19138 3840 19458 3841
rect 19138 3776 19146 3840
rect 19210 3776 19226 3840
rect 19290 3776 19306 3840
rect 19370 3776 19386 3840
rect 19450 3776 19458 3840
rect 19138 3775 19458 3776
rect 1289 3498 1355 3501
rect 10581 3498 10647 3501
rect 1289 3496 10647 3498
rect 1289 3440 1294 3496
rect 1350 3440 10586 3496
rect 10642 3440 10647 3496
rect 1289 3438 10647 3440
rect 1289 3435 1355 3438
rect 10581 3435 10647 3438
rect 24657 3498 24723 3501
rect 27048 3498 27528 3528
rect 24657 3496 27528 3498
rect 24657 3440 24662 3496
rect 24718 3440 27528 3496
rect 24657 3438 27528 3440
rect 24657 3435 24723 3438
rect 27048 3408 27528 3438
rect 5138 3296 5458 3297
rect 5138 3232 5146 3296
rect 5210 3232 5226 3296
rect 5290 3232 5306 3296
rect 5370 3232 5386 3296
rect 5450 3232 5458 3296
rect 5138 3231 5458 3232
rect 14472 3296 14792 3297
rect 14472 3232 14480 3296
rect 14544 3232 14560 3296
rect 14624 3232 14640 3296
rect 14704 3232 14720 3296
rect 14784 3232 14792 3296
rect 14472 3231 14792 3232
rect 23805 3296 24125 3297
rect 23805 3232 23813 3296
rect 23877 3232 23893 3296
rect 23957 3232 23973 3296
rect 24037 3232 24053 3296
rect 24117 3232 24125 3296
rect 23805 3231 24125 3232
rect 16285 2954 16351 2957
rect 16285 2952 23202 2954
rect 16285 2896 16290 2952
rect 16346 2896 23202 2952
rect 16285 2894 23202 2896
rect 16285 2891 16351 2894
rect 9805 2752 10125 2753
rect 9805 2688 9813 2752
rect 9877 2688 9893 2752
rect 9957 2688 9973 2752
rect 10037 2688 10053 2752
rect 10117 2688 10125 2752
rect 9805 2687 10125 2688
rect 19138 2752 19458 2753
rect 19138 2688 19146 2752
rect 19210 2688 19226 2752
rect 19290 2688 19306 2752
rect 19370 2688 19386 2752
rect 19450 2688 19458 2752
rect 19138 2687 19458 2688
rect 23142 2546 23202 2894
rect 27048 2546 27528 2576
rect 23142 2486 27528 2546
rect 27048 2456 27528 2486
rect 5138 2208 5458 2209
rect 5138 2144 5146 2208
rect 5210 2144 5226 2208
rect 5290 2144 5306 2208
rect 5370 2144 5386 2208
rect 5450 2144 5458 2208
rect 5138 2143 5458 2144
rect 14472 2208 14792 2209
rect 14472 2144 14480 2208
rect 14544 2144 14560 2208
rect 14624 2144 14640 2208
rect 14704 2144 14720 2208
rect 14784 2144 14792 2208
rect 14472 2143 14792 2144
rect 23805 2208 24125 2209
rect 23805 2144 23813 2208
rect 23877 2144 23893 2208
rect 23957 2144 23973 2208
rect 24037 2144 24053 2208
rect 24117 2144 24125 2208
rect 23805 2143 24125 2144
rect 24657 1458 24723 1461
rect 27048 1458 27528 1488
rect 24657 1456 27528 1458
rect 24657 1400 24662 1456
rect 24718 1400 27528 1456
rect 24657 1398 27528 1400
rect 24657 1395 24723 1398
rect 27048 1368 27528 1398
rect 25117 506 25183 509
rect 27048 506 27528 536
rect 25117 504 27528 506
rect 25117 448 25122 504
rect 25178 448 27528 504
rect 25117 446 27528 448
rect 25117 443 25183 446
rect 27048 416 27528 446
<< via3 >>
rect 9813 25596 9877 25600
rect 9813 25540 9817 25596
rect 9817 25540 9873 25596
rect 9873 25540 9877 25596
rect 9813 25536 9877 25540
rect 9893 25596 9957 25600
rect 9893 25540 9897 25596
rect 9897 25540 9953 25596
rect 9953 25540 9957 25596
rect 9893 25536 9957 25540
rect 9973 25596 10037 25600
rect 9973 25540 9977 25596
rect 9977 25540 10033 25596
rect 10033 25540 10037 25596
rect 9973 25536 10037 25540
rect 10053 25596 10117 25600
rect 10053 25540 10057 25596
rect 10057 25540 10113 25596
rect 10113 25540 10117 25596
rect 10053 25536 10117 25540
rect 19146 25596 19210 25600
rect 19146 25540 19150 25596
rect 19150 25540 19206 25596
rect 19206 25540 19210 25596
rect 19146 25536 19210 25540
rect 19226 25596 19290 25600
rect 19226 25540 19230 25596
rect 19230 25540 19286 25596
rect 19286 25540 19290 25596
rect 19226 25536 19290 25540
rect 19306 25596 19370 25600
rect 19306 25540 19310 25596
rect 19310 25540 19366 25596
rect 19366 25540 19370 25596
rect 19306 25536 19370 25540
rect 19386 25596 19450 25600
rect 19386 25540 19390 25596
rect 19390 25540 19446 25596
rect 19446 25540 19450 25596
rect 19386 25536 19450 25540
rect 5146 25052 5210 25056
rect 5146 24996 5150 25052
rect 5150 24996 5206 25052
rect 5206 24996 5210 25052
rect 5146 24992 5210 24996
rect 5226 25052 5290 25056
rect 5226 24996 5230 25052
rect 5230 24996 5286 25052
rect 5286 24996 5290 25052
rect 5226 24992 5290 24996
rect 5306 25052 5370 25056
rect 5306 24996 5310 25052
rect 5310 24996 5366 25052
rect 5366 24996 5370 25052
rect 5306 24992 5370 24996
rect 5386 25052 5450 25056
rect 5386 24996 5390 25052
rect 5390 24996 5446 25052
rect 5446 24996 5450 25052
rect 5386 24992 5450 24996
rect 14480 25052 14544 25056
rect 14480 24996 14484 25052
rect 14484 24996 14540 25052
rect 14540 24996 14544 25052
rect 14480 24992 14544 24996
rect 14560 25052 14624 25056
rect 14560 24996 14564 25052
rect 14564 24996 14620 25052
rect 14620 24996 14624 25052
rect 14560 24992 14624 24996
rect 14640 25052 14704 25056
rect 14640 24996 14644 25052
rect 14644 24996 14700 25052
rect 14700 24996 14704 25052
rect 14640 24992 14704 24996
rect 14720 25052 14784 25056
rect 14720 24996 14724 25052
rect 14724 24996 14780 25052
rect 14780 24996 14784 25052
rect 14720 24992 14784 24996
rect 23813 25052 23877 25056
rect 23813 24996 23817 25052
rect 23817 24996 23873 25052
rect 23873 24996 23877 25052
rect 23813 24992 23877 24996
rect 23893 25052 23957 25056
rect 23893 24996 23897 25052
rect 23897 24996 23953 25052
rect 23953 24996 23957 25052
rect 23893 24992 23957 24996
rect 23973 25052 24037 25056
rect 23973 24996 23977 25052
rect 23977 24996 24033 25052
rect 24033 24996 24037 25052
rect 23973 24992 24037 24996
rect 24053 25052 24117 25056
rect 24053 24996 24057 25052
rect 24057 24996 24113 25052
rect 24113 24996 24117 25052
rect 24053 24992 24117 24996
rect 9813 24508 9877 24512
rect 9813 24452 9817 24508
rect 9817 24452 9873 24508
rect 9873 24452 9877 24508
rect 9813 24448 9877 24452
rect 9893 24508 9957 24512
rect 9893 24452 9897 24508
rect 9897 24452 9953 24508
rect 9953 24452 9957 24508
rect 9893 24448 9957 24452
rect 9973 24508 10037 24512
rect 9973 24452 9977 24508
rect 9977 24452 10033 24508
rect 10033 24452 10037 24508
rect 9973 24448 10037 24452
rect 10053 24508 10117 24512
rect 10053 24452 10057 24508
rect 10057 24452 10113 24508
rect 10113 24452 10117 24508
rect 10053 24448 10117 24452
rect 19146 24508 19210 24512
rect 19146 24452 19150 24508
rect 19150 24452 19206 24508
rect 19206 24452 19210 24508
rect 19146 24448 19210 24452
rect 19226 24508 19290 24512
rect 19226 24452 19230 24508
rect 19230 24452 19286 24508
rect 19286 24452 19290 24508
rect 19226 24448 19290 24452
rect 19306 24508 19370 24512
rect 19306 24452 19310 24508
rect 19310 24452 19366 24508
rect 19366 24452 19370 24508
rect 19306 24448 19370 24452
rect 19386 24508 19450 24512
rect 19386 24452 19390 24508
rect 19390 24452 19446 24508
rect 19446 24452 19450 24508
rect 19386 24448 19450 24452
rect 5146 23964 5210 23968
rect 5146 23908 5150 23964
rect 5150 23908 5206 23964
rect 5206 23908 5210 23964
rect 5146 23904 5210 23908
rect 5226 23964 5290 23968
rect 5226 23908 5230 23964
rect 5230 23908 5286 23964
rect 5286 23908 5290 23964
rect 5226 23904 5290 23908
rect 5306 23964 5370 23968
rect 5306 23908 5310 23964
rect 5310 23908 5366 23964
rect 5366 23908 5370 23964
rect 5306 23904 5370 23908
rect 5386 23964 5450 23968
rect 5386 23908 5390 23964
rect 5390 23908 5446 23964
rect 5446 23908 5450 23964
rect 5386 23904 5450 23908
rect 14480 23964 14544 23968
rect 14480 23908 14484 23964
rect 14484 23908 14540 23964
rect 14540 23908 14544 23964
rect 14480 23904 14544 23908
rect 14560 23964 14624 23968
rect 14560 23908 14564 23964
rect 14564 23908 14620 23964
rect 14620 23908 14624 23964
rect 14560 23904 14624 23908
rect 14640 23964 14704 23968
rect 14640 23908 14644 23964
rect 14644 23908 14700 23964
rect 14700 23908 14704 23964
rect 14640 23904 14704 23908
rect 14720 23964 14784 23968
rect 14720 23908 14724 23964
rect 14724 23908 14780 23964
rect 14780 23908 14784 23964
rect 14720 23904 14784 23908
rect 23813 23964 23877 23968
rect 23813 23908 23817 23964
rect 23817 23908 23873 23964
rect 23873 23908 23877 23964
rect 23813 23904 23877 23908
rect 23893 23964 23957 23968
rect 23893 23908 23897 23964
rect 23897 23908 23953 23964
rect 23953 23908 23957 23964
rect 23893 23904 23957 23908
rect 23973 23964 24037 23968
rect 23973 23908 23977 23964
rect 23977 23908 24033 23964
rect 24033 23908 24037 23964
rect 23973 23904 24037 23908
rect 24053 23964 24117 23968
rect 24053 23908 24057 23964
rect 24057 23908 24113 23964
rect 24113 23908 24117 23964
rect 24053 23904 24117 23908
rect 9813 23420 9877 23424
rect 9813 23364 9817 23420
rect 9817 23364 9873 23420
rect 9873 23364 9877 23420
rect 9813 23360 9877 23364
rect 9893 23420 9957 23424
rect 9893 23364 9897 23420
rect 9897 23364 9953 23420
rect 9953 23364 9957 23420
rect 9893 23360 9957 23364
rect 9973 23420 10037 23424
rect 9973 23364 9977 23420
rect 9977 23364 10033 23420
rect 10033 23364 10037 23420
rect 9973 23360 10037 23364
rect 10053 23420 10117 23424
rect 10053 23364 10057 23420
rect 10057 23364 10113 23420
rect 10113 23364 10117 23420
rect 10053 23360 10117 23364
rect 19146 23420 19210 23424
rect 19146 23364 19150 23420
rect 19150 23364 19206 23420
rect 19206 23364 19210 23420
rect 19146 23360 19210 23364
rect 19226 23420 19290 23424
rect 19226 23364 19230 23420
rect 19230 23364 19286 23420
rect 19286 23364 19290 23420
rect 19226 23360 19290 23364
rect 19306 23420 19370 23424
rect 19306 23364 19310 23420
rect 19310 23364 19366 23420
rect 19366 23364 19370 23420
rect 19306 23360 19370 23364
rect 19386 23420 19450 23424
rect 19386 23364 19390 23420
rect 19390 23364 19446 23420
rect 19446 23364 19450 23420
rect 19386 23360 19450 23364
rect 5146 22876 5210 22880
rect 5146 22820 5150 22876
rect 5150 22820 5206 22876
rect 5206 22820 5210 22876
rect 5146 22816 5210 22820
rect 5226 22876 5290 22880
rect 5226 22820 5230 22876
rect 5230 22820 5286 22876
rect 5286 22820 5290 22876
rect 5226 22816 5290 22820
rect 5306 22876 5370 22880
rect 5306 22820 5310 22876
rect 5310 22820 5366 22876
rect 5366 22820 5370 22876
rect 5306 22816 5370 22820
rect 5386 22876 5450 22880
rect 5386 22820 5390 22876
rect 5390 22820 5446 22876
rect 5446 22820 5450 22876
rect 5386 22816 5450 22820
rect 14480 22876 14544 22880
rect 14480 22820 14484 22876
rect 14484 22820 14540 22876
rect 14540 22820 14544 22876
rect 14480 22816 14544 22820
rect 14560 22876 14624 22880
rect 14560 22820 14564 22876
rect 14564 22820 14620 22876
rect 14620 22820 14624 22876
rect 14560 22816 14624 22820
rect 14640 22876 14704 22880
rect 14640 22820 14644 22876
rect 14644 22820 14700 22876
rect 14700 22820 14704 22876
rect 14640 22816 14704 22820
rect 14720 22876 14784 22880
rect 14720 22820 14724 22876
rect 14724 22820 14780 22876
rect 14780 22820 14784 22876
rect 14720 22816 14784 22820
rect 23813 22876 23877 22880
rect 23813 22820 23817 22876
rect 23817 22820 23873 22876
rect 23873 22820 23877 22876
rect 23813 22816 23877 22820
rect 23893 22876 23957 22880
rect 23893 22820 23897 22876
rect 23897 22820 23953 22876
rect 23953 22820 23957 22876
rect 23893 22816 23957 22820
rect 23973 22876 24037 22880
rect 23973 22820 23977 22876
rect 23977 22820 24033 22876
rect 24033 22820 24037 22876
rect 23973 22816 24037 22820
rect 24053 22876 24117 22880
rect 24053 22820 24057 22876
rect 24057 22820 24113 22876
rect 24113 22820 24117 22876
rect 24053 22816 24117 22820
rect 9813 22332 9877 22336
rect 9813 22276 9817 22332
rect 9817 22276 9873 22332
rect 9873 22276 9877 22332
rect 9813 22272 9877 22276
rect 9893 22332 9957 22336
rect 9893 22276 9897 22332
rect 9897 22276 9953 22332
rect 9953 22276 9957 22332
rect 9893 22272 9957 22276
rect 9973 22332 10037 22336
rect 9973 22276 9977 22332
rect 9977 22276 10033 22332
rect 10033 22276 10037 22332
rect 9973 22272 10037 22276
rect 10053 22332 10117 22336
rect 10053 22276 10057 22332
rect 10057 22276 10113 22332
rect 10113 22276 10117 22332
rect 10053 22272 10117 22276
rect 19146 22332 19210 22336
rect 19146 22276 19150 22332
rect 19150 22276 19206 22332
rect 19206 22276 19210 22332
rect 19146 22272 19210 22276
rect 19226 22332 19290 22336
rect 19226 22276 19230 22332
rect 19230 22276 19286 22332
rect 19286 22276 19290 22332
rect 19226 22272 19290 22276
rect 19306 22332 19370 22336
rect 19306 22276 19310 22332
rect 19310 22276 19366 22332
rect 19366 22276 19370 22332
rect 19306 22272 19370 22276
rect 19386 22332 19450 22336
rect 19386 22276 19390 22332
rect 19390 22276 19446 22332
rect 19446 22276 19450 22332
rect 19386 22272 19450 22276
rect 5146 21788 5210 21792
rect 5146 21732 5150 21788
rect 5150 21732 5206 21788
rect 5206 21732 5210 21788
rect 5146 21728 5210 21732
rect 5226 21788 5290 21792
rect 5226 21732 5230 21788
rect 5230 21732 5286 21788
rect 5286 21732 5290 21788
rect 5226 21728 5290 21732
rect 5306 21788 5370 21792
rect 5306 21732 5310 21788
rect 5310 21732 5366 21788
rect 5366 21732 5370 21788
rect 5306 21728 5370 21732
rect 5386 21788 5450 21792
rect 5386 21732 5390 21788
rect 5390 21732 5446 21788
rect 5446 21732 5450 21788
rect 5386 21728 5450 21732
rect 14480 21788 14544 21792
rect 14480 21732 14484 21788
rect 14484 21732 14540 21788
rect 14540 21732 14544 21788
rect 14480 21728 14544 21732
rect 14560 21788 14624 21792
rect 14560 21732 14564 21788
rect 14564 21732 14620 21788
rect 14620 21732 14624 21788
rect 14560 21728 14624 21732
rect 14640 21788 14704 21792
rect 14640 21732 14644 21788
rect 14644 21732 14700 21788
rect 14700 21732 14704 21788
rect 14640 21728 14704 21732
rect 14720 21788 14784 21792
rect 14720 21732 14724 21788
rect 14724 21732 14780 21788
rect 14780 21732 14784 21788
rect 14720 21728 14784 21732
rect 23813 21788 23877 21792
rect 23813 21732 23817 21788
rect 23817 21732 23873 21788
rect 23873 21732 23877 21788
rect 23813 21728 23877 21732
rect 23893 21788 23957 21792
rect 23893 21732 23897 21788
rect 23897 21732 23953 21788
rect 23953 21732 23957 21788
rect 23893 21728 23957 21732
rect 23973 21788 24037 21792
rect 23973 21732 23977 21788
rect 23977 21732 24033 21788
rect 24033 21732 24037 21788
rect 23973 21728 24037 21732
rect 24053 21788 24117 21792
rect 24053 21732 24057 21788
rect 24057 21732 24113 21788
rect 24113 21732 24117 21788
rect 24053 21728 24117 21732
rect 9813 21244 9877 21248
rect 9813 21188 9817 21244
rect 9817 21188 9873 21244
rect 9873 21188 9877 21244
rect 9813 21184 9877 21188
rect 9893 21244 9957 21248
rect 9893 21188 9897 21244
rect 9897 21188 9953 21244
rect 9953 21188 9957 21244
rect 9893 21184 9957 21188
rect 9973 21244 10037 21248
rect 9973 21188 9977 21244
rect 9977 21188 10033 21244
rect 10033 21188 10037 21244
rect 9973 21184 10037 21188
rect 10053 21244 10117 21248
rect 10053 21188 10057 21244
rect 10057 21188 10113 21244
rect 10113 21188 10117 21244
rect 10053 21184 10117 21188
rect 19146 21244 19210 21248
rect 19146 21188 19150 21244
rect 19150 21188 19206 21244
rect 19206 21188 19210 21244
rect 19146 21184 19210 21188
rect 19226 21244 19290 21248
rect 19226 21188 19230 21244
rect 19230 21188 19286 21244
rect 19286 21188 19290 21244
rect 19226 21184 19290 21188
rect 19306 21244 19370 21248
rect 19306 21188 19310 21244
rect 19310 21188 19366 21244
rect 19366 21188 19370 21244
rect 19306 21184 19370 21188
rect 19386 21244 19450 21248
rect 19386 21188 19390 21244
rect 19390 21188 19446 21244
rect 19446 21188 19450 21244
rect 19386 21184 19450 21188
rect 5146 20700 5210 20704
rect 5146 20644 5150 20700
rect 5150 20644 5206 20700
rect 5206 20644 5210 20700
rect 5146 20640 5210 20644
rect 5226 20700 5290 20704
rect 5226 20644 5230 20700
rect 5230 20644 5286 20700
rect 5286 20644 5290 20700
rect 5226 20640 5290 20644
rect 5306 20700 5370 20704
rect 5306 20644 5310 20700
rect 5310 20644 5366 20700
rect 5366 20644 5370 20700
rect 5306 20640 5370 20644
rect 5386 20700 5450 20704
rect 5386 20644 5390 20700
rect 5390 20644 5446 20700
rect 5446 20644 5450 20700
rect 5386 20640 5450 20644
rect 14480 20700 14544 20704
rect 14480 20644 14484 20700
rect 14484 20644 14540 20700
rect 14540 20644 14544 20700
rect 14480 20640 14544 20644
rect 14560 20700 14624 20704
rect 14560 20644 14564 20700
rect 14564 20644 14620 20700
rect 14620 20644 14624 20700
rect 14560 20640 14624 20644
rect 14640 20700 14704 20704
rect 14640 20644 14644 20700
rect 14644 20644 14700 20700
rect 14700 20644 14704 20700
rect 14640 20640 14704 20644
rect 14720 20700 14784 20704
rect 14720 20644 14724 20700
rect 14724 20644 14780 20700
rect 14780 20644 14784 20700
rect 14720 20640 14784 20644
rect 23813 20700 23877 20704
rect 23813 20644 23817 20700
rect 23817 20644 23873 20700
rect 23873 20644 23877 20700
rect 23813 20640 23877 20644
rect 23893 20700 23957 20704
rect 23893 20644 23897 20700
rect 23897 20644 23953 20700
rect 23953 20644 23957 20700
rect 23893 20640 23957 20644
rect 23973 20700 24037 20704
rect 23973 20644 23977 20700
rect 23977 20644 24033 20700
rect 24033 20644 24037 20700
rect 23973 20640 24037 20644
rect 24053 20700 24117 20704
rect 24053 20644 24057 20700
rect 24057 20644 24113 20700
rect 24113 20644 24117 20700
rect 24053 20640 24117 20644
rect 9813 20156 9877 20160
rect 9813 20100 9817 20156
rect 9817 20100 9873 20156
rect 9873 20100 9877 20156
rect 9813 20096 9877 20100
rect 9893 20156 9957 20160
rect 9893 20100 9897 20156
rect 9897 20100 9953 20156
rect 9953 20100 9957 20156
rect 9893 20096 9957 20100
rect 9973 20156 10037 20160
rect 9973 20100 9977 20156
rect 9977 20100 10033 20156
rect 10033 20100 10037 20156
rect 9973 20096 10037 20100
rect 10053 20156 10117 20160
rect 10053 20100 10057 20156
rect 10057 20100 10113 20156
rect 10113 20100 10117 20156
rect 10053 20096 10117 20100
rect 19146 20156 19210 20160
rect 19146 20100 19150 20156
rect 19150 20100 19206 20156
rect 19206 20100 19210 20156
rect 19146 20096 19210 20100
rect 19226 20156 19290 20160
rect 19226 20100 19230 20156
rect 19230 20100 19286 20156
rect 19286 20100 19290 20156
rect 19226 20096 19290 20100
rect 19306 20156 19370 20160
rect 19306 20100 19310 20156
rect 19310 20100 19366 20156
rect 19366 20100 19370 20156
rect 19306 20096 19370 20100
rect 19386 20156 19450 20160
rect 19386 20100 19390 20156
rect 19390 20100 19446 20156
rect 19446 20100 19450 20156
rect 19386 20096 19450 20100
rect 5146 19612 5210 19616
rect 5146 19556 5150 19612
rect 5150 19556 5206 19612
rect 5206 19556 5210 19612
rect 5146 19552 5210 19556
rect 5226 19612 5290 19616
rect 5226 19556 5230 19612
rect 5230 19556 5286 19612
rect 5286 19556 5290 19612
rect 5226 19552 5290 19556
rect 5306 19612 5370 19616
rect 5306 19556 5310 19612
rect 5310 19556 5366 19612
rect 5366 19556 5370 19612
rect 5306 19552 5370 19556
rect 5386 19612 5450 19616
rect 5386 19556 5390 19612
rect 5390 19556 5446 19612
rect 5446 19556 5450 19612
rect 5386 19552 5450 19556
rect 14480 19612 14544 19616
rect 14480 19556 14484 19612
rect 14484 19556 14540 19612
rect 14540 19556 14544 19612
rect 14480 19552 14544 19556
rect 14560 19612 14624 19616
rect 14560 19556 14564 19612
rect 14564 19556 14620 19612
rect 14620 19556 14624 19612
rect 14560 19552 14624 19556
rect 14640 19612 14704 19616
rect 14640 19556 14644 19612
rect 14644 19556 14700 19612
rect 14700 19556 14704 19612
rect 14640 19552 14704 19556
rect 14720 19612 14784 19616
rect 14720 19556 14724 19612
rect 14724 19556 14780 19612
rect 14780 19556 14784 19612
rect 14720 19552 14784 19556
rect 23813 19612 23877 19616
rect 23813 19556 23817 19612
rect 23817 19556 23873 19612
rect 23873 19556 23877 19612
rect 23813 19552 23877 19556
rect 23893 19612 23957 19616
rect 23893 19556 23897 19612
rect 23897 19556 23953 19612
rect 23953 19556 23957 19612
rect 23893 19552 23957 19556
rect 23973 19612 24037 19616
rect 23973 19556 23977 19612
rect 23977 19556 24033 19612
rect 24033 19556 24037 19612
rect 23973 19552 24037 19556
rect 24053 19612 24117 19616
rect 24053 19556 24057 19612
rect 24057 19556 24113 19612
rect 24113 19556 24117 19612
rect 24053 19552 24117 19556
rect 9813 19068 9877 19072
rect 9813 19012 9817 19068
rect 9817 19012 9873 19068
rect 9873 19012 9877 19068
rect 9813 19008 9877 19012
rect 9893 19068 9957 19072
rect 9893 19012 9897 19068
rect 9897 19012 9953 19068
rect 9953 19012 9957 19068
rect 9893 19008 9957 19012
rect 9973 19068 10037 19072
rect 9973 19012 9977 19068
rect 9977 19012 10033 19068
rect 10033 19012 10037 19068
rect 9973 19008 10037 19012
rect 10053 19068 10117 19072
rect 10053 19012 10057 19068
rect 10057 19012 10113 19068
rect 10113 19012 10117 19068
rect 10053 19008 10117 19012
rect 19146 19068 19210 19072
rect 19146 19012 19150 19068
rect 19150 19012 19206 19068
rect 19206 19012 19210 19068
rect 19146 19008 19210 19012
rect 19226 19068 19290 19072
rect 19226 19012 19230 19068
rect 19230 19012 19286 19068
rect 19286 19012 19290 19068
rect 19226 19008 19290 19012
rect 19306 19068 19370 19072
rect 19306 19012 19310 19068
rect 19310 19012 19366 19068
rect 19366 19012 19370 19068
rect 19306 19008 19370 19012
rect 19386 19068 19450 19072
rect 19386 19012 19390 19068
rect 19390 19012 19446 19068
rect 19446 19012 19450 19068
rect 19386 19008 19450 19012
rect 5146 18524 5210 18528
rect 5146 18468 5150 18524
rect 5150 18468 5206 18524
rect 5206 18468 5210 18524
rect 5146 18464 5210 18468
rect 5226 18524 5290 18528
rect 5226 18468 5230 18524
rect 5230 18468 5286 18524
rect 5286 18468 5290 18524
rect 5226 18464 5290 18468
rect 5306 18524 5370 18528
rect 5306 18468 5310 18524
rect 5310 18468 5366 18524
rect 5366 18468 5370 18524
rect 5306 18464 5370 18468
rect 5386 18524 5450 18528
rect 5386 18468 5390 18524
rect 5390 18468 5446 18524
rect 5446 18468 5450 18524
rect 5386 18464 5450 18468
rect 14480 18524 14544 18528
rect 14480 18468 14484 18524
rect 14484 18468 14540 18524
rect 14540 18468 14544 18524
rect 14480 18464 14544 18468
rect 14560 18524 14624 18528
rect 14560 18468 14564 18524
rect 14564 18468 14620 18524
rect 14620 18468 14624 18524
rect 14560 18464 14624 18468
rect 14640 18524 14704 18528
rect 14640 18468 14644 18524
rect 14644 18468 14700 18524
rect 14700 18468 14704 18524
rect 14640 18464 14704 18468
rect 14720 18524 14784 18528
rect 14720 18468 14724 18524
rect 14724 18468 14780 18524
rect 14780 18468 14784 18524
rect 14720 18464 14784 18468
rect 23813 18524 23877 18528
rect 23813 18468 23817 18524
rect 23817 18468 23873 18524
rect 23873 18468 23877 18524
rect 23813 18464 23877 18468
rect 23893 18524 23957 18528
rect 23893 18468 23897 18524
rect 23897 18468 23953 18524
rect 23953 18468 23957 18524
rect 23893 18464 23957 18468
rect 23973 18524 24037 18528
rect 23973 18468 23977 18524
rect 23977 18468 24033 18524
rect 24033 18468 24037 18524
rect 23973 18464 24037 18468
rect 24053 18524 24117 18528
rect 24053 18468 24057 18524
rect 24057 18468 24113 18524
rect 24113 18468 24117 18524
rect 24053 18464 24117 18468
rect 9813 17980 9877 17984
rect 9813 17924 9817 17980
rect 9817 17924 9873 17980
rect 9873 17924 9877 17980
rect 9813 17920 9877 17924
rect 9893 17980 9957 17984
rect 9893 17924 9897 17980
rect 9897 17924 9953 17980
rect 9953 17924 9957 17980
rect 9893 17920 9957 17924
rect 9973 17980 10037 17984
rect 9973 17924 9977 17980
rect 9977 17924 10033 17980
rect 10033 17924 10037 17980
rect 9973 17920 10037 17924
rect 10053 17980 10117 17984
rect 10053 17924 10057 17980
rect 10057 17924 10113 17980
rect 10113 17924 10117 17980
rect 10053 17920 10117 17924
rect 19146 17980 19210 17984
rect 19146 17924 19150 17980
rect 19150 17924 19206 17980
rect 19206 17924 19210 17980
rect 19146 17920 19210 17924
rect 19226 17980 19290 17984
rect 19226 17924 19230 17980
rect 19230 17924 19286 17980
rect 19286 17924 19290 17980
rect 19226 17920 19290 17924
rect 19306 17980 19370 17984
rect 19306 17924 19310 17980
rect 19310 17924 19366 17980
rect 19366 17924 19370 17980
rect 19306 17920 19370 17924
rect 19386 17980 19450 17984
rect 19386 17924 19390 17980
rect 19390 17924 19446 17980
rect 19446 17924 19450 17980
rect 19386 17920 19450 17924
rect 5146 17436 5210 17440
rect 5146 17380 5150 17436
rect 5150 17380 5206 17436
rect 5206 17380 5210 17436
rect 5146 17376 5210 17380
rect 5226 17436 5290 17440
rect 5226 17380 5230 17436
rect 5230 17380 5286 17436
rect 5286 17380 5290 17436
rect 5226 17376 5290 17380
rect 5306 17436 5370 17440
rect 5306 17380 5310 17436
rect 5310 17380 5366 17436
rect 5366 17380 5370 17436
rect 5306 17376 5370 17380
rect 5386 17436 5450 17440
rect 5386 17380 5390 17436
rect 5390 17380 5446 17436
rect 5446 17380 5450 17436
rect 5386 17376 5450 17380
rect 14480 17436 14544 17440
rect 14480 17380 14484 17436
rect 14484 17380 14540 17436
rect 14540 17380 14544 17436
rect 14480 17376 14544 17380
rect 14560 17436 14624 17440
rect 14560 17380 14564 17436
rect 14564 17380 14620 17436
rect 14620 17380 14624 17436
rect 14560 17376 14624 17380
rect 14640 17436 14704 17440
rect 14640 17380 14644 17436
rect 14644 17380 14700 17436
rect 14700 17380 14704 17436
rect 14640 17376 14704 17380
rect 14720 17436 14784 17440
rect 14720 17380 14724 17436
rect 14724 17380 14780 17436
rect 14780 17380 14784 17436
rect 14720 17376 14784 17380
rect 23813 17436 23877 17440
rect 23813 17380 23817 17436
rect 23817 17380 23873 17436
rect 23873 17380 23877 17436
rect 23813 17376 23877 17380
rect 23893 17436 23957 17440
rect 23893 17380 23897 17436
rect 23897 17380 23953 17436
rect 23953 17380 23957 17436
rect 23893 17376 23957 17380
rect 23973 17436 24037 17440
rect 23973 17380 23977 17436
rect 23977 17380 24033 17436
rect 24033 17380 24037 17436
rect 23973 17376 24037 17380
rect 24053 17436 24117 17440
rect 24053 17380 24057 17436
rect 24057 17380 24113 17436
rect 24113 17380 24117 17436
rect 24053 17376 24117 17380
rect 9813 16892 9877 16896
rect 9813 16836 9817 16892
rect 9817 16836 9873 16892
rect 9873 16836 9877 16892
rect 9813 16832 9877 16836
rect 9893 16892 9957 16896
rect 9893 16836 9897 16892
rect 9897 16836 9953 16892
rect 9953 16836 9957 16892
rect 9893 16832 9957 16836
rect 9973 16892 10037 16896
rect 9973 16836 9977 16892
rect 9977 16836 10033 16892
rect 10033 16836 10037 16892
rect 9973 16832 10037 16836
rect 10053 16892 10117 16896
rect 10053 16836 10057 16892
rect 10057 16836 10113 16892
rect 10113 16836 10117 16892
rect 10053 16832 10117 16836
rect 19146 16892 19210 16896
rect 19146 16836 19150 16892
rect 19150 16836 19206 16892
rect 19206 16836 19210 16892
rect 19146 16832 19210 16836
rect 19226 16892 19290 16896
rect 19226 16836 19230 16892
rect 19230 16836 19286 16892
rect 19286 16836 19290 16892
rect 19226 16832 19290 16836
rect 19306 16892 19370 16896
rect 19306 16836 19310 16892
rect 19310 16836 19366 16892
rect 19366 16836 19370 16892
rect 19306 16832 19370 16836
rect 19386 16892 19450 16896
rect 19386 16836 19390 16892
rect 19390 16836 19446 16892
rect 19446 16836 19450 16892
rect 19386 16832 19450 16836
rect 5146 16348 5210 16352
rect 5146 16292 5150 16348
rect 5150 16292 5206 16348
rect 5206 16292 5210 16348
rect 5146 16288 5210 16292
rect 5226 16348 5290 16352
rect 5226 16292 5230 16348
rect 5230 16292 5286 16348
rect 5286 16292 5290 16348
rect 5226 16288 5290 16292
rect 5306 16348 5370 16352
rect 5306 16292 5310 16348
rect 5310 16292 5366 16348
rect 5366 16292 5370 16348
rect 5306 16288 5370 16292
rect 5386 16348 5450 16352
rect 5386 16292 5390 16348
rect 5390 16292 5446 16348
rect 5446 16292 5450 16348
rect 5386 16288 5450 16292
rect 14480 16348 14544 16352
rect 14480 16292 14484 16348
rect 14484 16292 14540 16348
rect 14540 16292 14544 16348
rect 14480 16288 14544 16292
rect 14560 16348 14624 16352
rect 14560 16292 14564 16348
rect 14564 16292 14620 16348
rect 14620 16292 14624 16348
rect 14560 16288 14624 16292
rect 14640 16348 14704 16352
rect 14640 16292 14644 16348
rect 14644 16292 14700 16348
rect 14700 16292 14704 16348
rect 14640 16288 14704 16292
rect 14720 16348 14784 16352
rect 14720 16292 14724 16348
rect 14724 16292 14780 16348
rect 14780 16292 14784 16348
rect 14720 16288 14784 16292
rect 23813 16348 23877 16352
rect 23813 16292 23817 16348
rect 23817 16292 23873 16348
rect 23873 16292 23877 16348
rect 23813 16288 23877 16292
rect 23893 16348 23957 16352
rect 23893 16292 23897 16348
rect 23897 16292 23953 16348
rect 23953 16292 23957 16348
rect 23893 16288 23957 16292
rect 23973 16348 24037 16352
rect 23973 16292 23977 16348
rect 23977 16292 24033 16348
rect 24033 16292 24037 16348
rect 23973 16288 24037 16292
rect 24053 16348 24117 16352
rect 24053 16292 24057 16348
rect 24057 16292 24113 16348
rect 24113 16292 24117 16348
rect 24053 16288 24117 16292
rect 9813 15804 9877 15808
rect 9813 15748 9817 15804
rect 9817 15748 9873 15804
rect 9873 15748 9877 15804
rect 9813 15744 9877 15748
rect 9893 15804 9957 15808
rect 9893 15748 9897 15804
rect 9897 15748 9953 15804
rect 9953 15748 9957 15804
rect 9893 15744 9957 15748
rect 9973 15804 10037 15808
rect 9973 15748 9977 15804
rect 9977 15748 10033 15804
rect 10033 15748 10037 15804
rect 9973 15744 10037 15748
rect 10053 15804 10117 15808
rect 10053 15748 10057 15804
rect 10057 15748 10113 15804
rect 10113 15748 10117 15804
rect 10053 15744 10117 15748
rect 19146 15804 19210 15808
rect 19146 15748 19150 15804
rect 19150 15748 19206 15804
rect 19206 15748 19210 15804
rect 19146 15744 19210 15748
rect 19226 15804 19290 15808
rect 19226 15748 19230 15804
rect 19230 15748 19286 15804
rect 19286 15748 19290 15804
rect 19226 15744 19290 15748
rect 19306 15804 19370 15808
rect 19306 15748 19310 15804
rect 19310 15748 19366 15804
rect 19366 15748 19370 15804
rect 19306 15744 19370 15748
rect 19386 15804 19450 15808
rect 19386 15748 19390 15804
rect 19390 15748 19446 15804
rect 19446 15748 19450 15804
rect 19386 15744 19450 15748
rect 5146 15260 5210 15264
rect 5146 15204 5150 15260
rect 5150 15204 5206 15260
rect 5206 15204 5210 15260
rect 5146 15200 5210 15204
rect 5226 15260 5290 15264
rect 5226 15204 5230 15260
rect 5230 15204 5286 15260
rect 5286 15204 5290 15260
rect 5226 15200 5290 15204
rect 5306 15260 5370 15264
rect 5306 15204 5310 15260
rect 5310 15204 5366 15260
rect 5366 15204 5370 15260
rect 5306 15200 5370 15204
rect 5386 15260 5450 15264
rect 5386 15204 5390 15260
rect 5390 15204 5446 15260
rect 5446 15204 5450 15260
rect 5386 15200 5450 15204
rect 14480 15260 14544 15264
rect 14480 15204 14484 15260
rect 14484 15204 14540 15260
rect 14540 15204 14544 15260
rect 14480 15200 14544 15204
rect 14560 15260 14624 15264
rect 14560 15204 14564 15260
rect 14564 15204 14620 15260
rect 14620 15204 14624 15260
rect 14560 15200 14624 15204
rect 14640 15260 14704 15264
rect 14640 15204 14644 15260
rect 14644 15204 14700 15260
rect 14700 15204 14704 15260
rect 14640 15200 14704 15204
rect 14720 15260 14784 15264
rect 14720 15204 14724 15260
rect 14724 15204 14780 15260
rect 14780 15204 14784 15260
rect 14720 15200 14784 15204
rect 23813 15260 23877 15264
rect 23813 15204 23817 15260
rect 23817 15204 23873 15260
rect 23873 15204 23877 15260
rect 23813 15200 23877 15204
rect 23893 15260 23957 15264
rect 23893 15204 23897 15260
rect 23897 15204 23953 15260
rect 23953 15204 23957 15260
rect 23893 15200 23957 15204
rect 23973 15260 24037 15264
rect 23973 15204 23977 15260
rect 23977 15204 24033 15260
rect 24033 15204 24037 15260
rect 23973 15200 24037 15204
rect 24053 15260 24117 15264
rect 24053 15204 24057 15260
rect 24057 15204 24113 15260
rect 24113 15204 24117 15260
rect 24053 15200 24117 15204
rect 9813 14716 9877 14720
rect 9813 14660 9817 14716
rect 9817 14660 9873 14716
rect 9873 14660 9877 14716
rect 9813 14656 9877 14660
rect 9893 14716 9957 14720
rect 9893 14660 9897 14716
rect 9897 14660 9953 14716
rect 9953 14660 9957 14716
rect 9893 14656 9957 14660
rect 9973 14716 10037 14720
rect 9973 14660 9977 14716
rect 9977 14660 10033 14716
rect 10033 14660 10037 14716
rect 9973 14656 10037 14660
rect 10053 14716 10117 14720
rect 10053 14660 10057 14716
rect 10057 14660 10113 14716
rect 10113 14660 10117 14716
rect 10053 14656 10117 14660
rect 19146 14716 19210 14720
rect 19146 14660 19150 14716
rect 19150 14660 19206 14716
rect 19206 14660 19210 14716
rect 19146 14656 19210 14660
rect 19226 14716 19290 14720
rect 19226 14660 19230 14716
rect 19230 14660 19286 14716
rect 19286 14660 19290 14716
rect 19226 14656 19290 14660
rect 19306 14716 19370 14720
rect 19306 14660 19310 14716
rect 19310 14660 19366 14716
rect 19366 14660 19370 14716
rect 19306 14656 19370 14660
rect 19386 14716 19450 14720
rect 19386 14660 19390 14716
rect 19390 14660 19446 14716
rect 19446 14660 19450 14716
rect 19386 14656 19450 14660
rect 5146 14172 5210 14176
rect 5146 14116 5150 14172
rect 5150 14116 5206 14172
rect 5206 14116 5210 14172
rect 5146 14112 5210 14116
rect 5226 14172 5290 14176
rect 5226 14116 5230 14172
rect 5230 14116 5286 14172
rect 5286 14116 5290 14172
rect 5226 14112 5290 14116
rect 5306 14172 5370 14176
rect 5306 14116 5310 14172
rect 5310 14116 5366 14172
rect 5366 14116 5370 14172
rect 5306 14112 5370 14116
rect 5386 14172 5450 14176
rect 5386 14116 5390 14172
rect 5390 14116 5446 14172
rect 5446 14116 5450 14172
rect 5386 14112 5450 14116
rect 14480 14172 14544 14176
rect 14480 14116 14484 14172
rect 14484 14116 14540 14172
rect 14540 14116 14544 14172
rect 14480 14112 14544 14116
rect 14560 14172 14624 14176
rect 14560 14116 14564 14172
rect 14564 14116 14620 14172
rect 14620 14116 14624 14172
rect 14560 14112 14624 14116
rect 14640 14172 14704 14176
rect 14640 14116 14644 14172
rect 14644 14116 14700 14172
rect 14700 14116 14704 14172
rect 14640 14112 14704 14116
rect 14720 14172 14784 14176
rect 14720 14116 14724 14172
rect 14724 14116 14780 14172
rect 14780 14116 14784 14172
rect 14720 14112 14784 14116
rect 23813 14172 23877 14176
rect 23813 14116 23817 14172
rect 23817 14116 23873 14172
rect 23873 14116 23877 14172
rect 23813 14112 23877 14116
rect 23893 14172 23957 14176
rect 23893 14116 23897 14172
rect 23897 14116 23953 14172
rect 23953 14116 23957 14172
rect 23893 14112 23957 14116
rect 23973 14172 24037 14176
rect 23973 14116 23977 14172
rect 23977 14116 24033 14172
rect 24033 14116 24037 14172
rect 23973 14112 24037 14116
rect 24053 14172 24117 14176
rect 24053 14116 24057 14172
rect 24057 14116 24113 14172
rect 24113 14116 24117 14172
rect 24053 14112 24117 14116
rect 24244 13908 24308 13972
rect 9813 13628 9877 13632
rect 9813 13572 9817 13628
rect 9817 13572 9873 13628
rect 9873 13572 9877 13628
rect 9813 13568 9877 13572
rect 9893 13628 9957 13632
rect 9893 13572 9897 13628
rect 9897 13572 9953 13628
rect 9953 13572 9957 13628
rect 9893 13568 9957 13572
rect 9973 13628 10037 13632
rect 9973 13572 9977 13628
rect 9977 13572 10033 13628
rect 10033 13572 10037 13628
rect 9973 13568 10037 13572
rect 10053 13628 10117 13632
rect 10053 13572 10057 13628
rect 10057 13572 10113 13628
rect 10113 13572 10117 13628
rect 10053 13568 10117 13572
rect 19146 13628 19210 13632
rect 19146 13572 19150 13628
rect 19150 13572 19206 13628
rect 19206 13572 19210 13628
rect 19146 13568 19210 13572
rect 19226 13628 19290 13632
rect 19226 13572 19230 13628
rect 19230 13572 19286 13628
rect 19286 13572 19290 13628
rect 19226 13568 19290 13572
rect 19306 13628 19370 13632
rect 19306 13572 19310 13628
rect 19310 13572 19366 13628
rect 19366 13572 19370 13628
rect 19306 13568 19370 13572
rect 19386 13628 19450 13632
rect 19386 13572 19390 13628
rect 19390 13572 19446 13628
rect 19446 13572 19450 13628
rect 19386 13568 19450 13572
rect 5146 13084 5210 13088
rect 5146 13028 5150 13084
rect 5150 13028 5206 13084
rect 5206 13028 5210 13084
rect 5146 13024 5210 13028
rect 5226 13084 5290 13088
rect 5226 13028 5230 13084
rect 5230 13028 5286 13084
rect 5286 13028 5290 13084
rect 5226 13024 5290 13028
rect 5306 13084 5370 13088
rect 5306 13028 5310 13084
rect 5310 13028 5366 13084
rect 5366 13028 5370 13084
rect 5306 13024 5370 13028
rect 5386 13084 5450 13088
rect 5386 13028 5390 13084
rect 5390 13028 5446 13084
rect 5446 13028 5450 13084
rect 5386 13024 5450 13028
rect 14480 13084 14544 13088
rect 14480 13028 14484 13084
rect 14484 13028 14540 13084
rect 14540 13028 14544 13084
rect 14480 13024 14544 13028
rect 14560 13084 14624 13088
rect 14560 13028 14564 13084
rect 14564 13028 14620 13084
rect 14620 13028 14624 13084
rect 14560 13024 14624 13028
rect 14640 13084 14704 13088
rect 14640 13028 14644 13084
rect 14644 13028 14700 13084
rect 14700 13028 14704 13084
rect 14640 13024 14704 13028
rect 14720 13084 14784 13088
rect 14720 13028 14724 13084
rect 14724 13028 14780 13084
rect 14780 13028 14784 13084
rect 14720 13024 14784 13028
rect 23813 13084 23877 13088
rect 23813 13028 23817 13084
rect 23817 13028 23873 13084
rect 23873 13028 23877 13084
rect 23813 13024 23877 13028
rect 23893 13084 23957 13088
rect 23893 13028 23897 13084
rect 23897 13028 23953 13084
rect 23953 13028 23957 13084
rect 23893 13024 23957 13028
rect 23973 13084 24037 13088
rect 23973 13028 23977 13084
rect 23977 13028 24033 13084
rect 24033 13028 24037 13084
rect 23973 13024 24037 13028
rect 24053 13084 24117 13088
rect 24053 13028 24057 13084
rect 24057 13028 24113 13084
rect 24113 13028 24117 13084
rect 24053 13024 24117 13028
rect 9813 12540 9877 12544
rect 9813 12484 9817 12540
rect 9817 12484 9873 12540
rect 9873 12484 9877 12540
rect 9813 12480 9877 12484
rect 9893 12540 9957 12544
rect 9893 12484 9897 12540
rect 9897 12484 9953 12540
rect 9953 12484 9957 12540
rect 9893 12480 9957 12484
rect 9973 12540 10037 12544
rect 9973 12484 9977 12540
rect 9977 12484 10033 12540
rect 10033 12484 10037 12540
rect 9973 12480 10037 12484
rect 10053 12540 10117 12544
rect 10053 12484 10057 12540
rect 10057 12484 10113 12540
rect 10113 12484 10117 12540
rect 10053 12480 10117 12484
rect 19146 12540 19210 12544
rect 19146 12484 19150 12540
rect 19150 12484 19206 12540
rect 19206 12484 19210 12540
rect 19146 12480 19210 12484
rect 19226 12540 19290 12544
rect 19226 12484 19230 12540
rect 19230 12484 19286 12540
rect 19286 12484 19290 12540
rect 19226 12480 19290 12484
rect 19306 12540 19370 12544
rect 19306 12484 19310 12540
rect 19310 12484 19366 12540
rect 19366 12484 19370 12540
rect 19306 12480 19370 12484
rect 19386 12540 19450 12544
rect 19386 12484 19390 12540
rect 19390 12484 19446 12540
rect 19446 12484 19450 12540
rect 19386 12480 19450 12484
rect 5146 11996 5210 12000
rect 5146 11940 5150 11996
rect 5150 11940 5206 11996
rect 5206 11940 5210 11996
rect 5146 11936 5210 11940
rect 5226 11996 5290 12000
rect 5226 11940 5230 11996
rect 5230 11940 5286 11996
rect 5286 11940 5290 11996
rect 5226 11936 5290 11940
rect 5306 11996 5370 12000
rect 5306 11940 5310 11996
rect 5310 11940 5366 11996
rect 5366 11940 5370 11996
rect 5306 11936 5370 11940
rect 5386 11996 5450 12000
rect 5386 11940 5390 11996
rect 5390 11940 5446 11996
rect 5446 11940 5450 11996
rect 5386 11936 5450 11940
rect 14480 11996 14544 12000
rect 14480 11940 14484 11996
rect 14484 11940 14540 11996
rect 14540 11940 14544 11996
rect 14480 11936 14544 11940
rect 14560 11996 14624 12000
rect 14560 11940 14564 11996
rect 14564 11940 14620 11996
rect 14620 11940 14624 11996
rect 14560 11936 14624 11940
rect 14640 11996 14704 12000
rect 14640 11940 14644 11996
rect 14644 11940 14700 11996
rect 14700 11940 14704 11996
rect 14640 11936 14704 11940
rect 14720 11996 14784 12000
rect 14720 11940 14724 11996
rect 14724 11940 14780 11996
rect 14780 11940 14784 11996
rect 14720 11936 14784 11940
rect 23813 11996 23877 12000
rect 23813 11940 23817 11996
rect 23817 11940 23873 11996
rect 23873 11940 23877 11996
rect 23813 11936 23877 11940
rect 23893 11996 23957 12000
rect 23893 11940 23897 11996
rect 23897 11940 23953 11996
rect 23953 11940 23957 11996
rect 23893 11936 23957 11940
rect 23973 11996 24037 12000
rect 23973 11940 23977 11996
rect 23977 11940 24033 11996
rect 24033 11940 24037 11996
rect 23973 11936 24037 11940
rect 24053 11996 24117 12000
rect 24053 11940 24057 11996
rect 24057 11940 24113 11996
rect 24113 11940 24117 11996
rect 24053 11936 24117 11940
rect 9813 11452 9877 11456
rect 9813 11396 9817 11452
rect 9817 11396 9873 11452
rect 9873 11396 9877 11452
rect 9813 11392 9877 11396
rect 9893 11452 9957 11456
rect 9893 11396 9897 11452
rect 9897 11396 9953 11452
rect 9953 11396 9957 11452
rect 9893 11392 9957 11396
rect 9973 11452 10037 11456
rect 9973 11396 9977 11452
rect 9977 11396 10033 11452
rect 10033 11396 10037 11452
rect 9973 11392 10037 11396
rect 10053 11452 10117 11456
rect 10053 11396 10057 11452
rect 10057 11396 10113 11452
rect 10113 11396 10117 11452
rect 10053 11392 10117 11396
rect 19146 11452 19210 11456
rect 19146 11396 19150 11452
rect 19150 11396 19206 11452
rect 19206 11396 19210 11452
rect 19146 11392 19210 11396
rect 19226 11452 19290 11456
rect 19226 11396 19230 11452
rect 19230 11396 19286 11452
rect 19286 11396 19290 11452
rect 19226 11392 19290 11396
rect 19306 11452 19370 11456
rect 19306 11396 19310 11452
rect 19310 11396 19366 11452
rect 19366 11396 19370 11452
rect 19306 11392 19370 11396
rect 19386 11452 19450 11456
rect 19386 11396 19390 11452
rect 19390 11396 19446 11452
rect 19446 11396 19450 11452
rect 19386 11392 19450 11396
rect 5146 10908 5210 10912
rect 5146 10852 5150 10908
rect 5150 10852 5206 10908
rect 5206 10852 5210 10908
rect 5146 10848 5210 10852
rect 5226 10908 5290 10912
rect 5226 10852 5230 10908
rect 5230 10852 5286 10908
rect 5286 10852 5290 10908
rect 5226 10848 5290 10852
rect 5306 10908 5370 10912
rect 5306 10852 5310 10908
rect 5310 10852 5366 10908
rect 5366 10852 5370 10908
rect 5306 10848 5370 10852
rect 5386 10908 5450 10912
rect 5386 10852 5390 10908
rect 5390 10852 5446 10908
rect 5446 10852 5450 10908
rect 5386 10848 5450 10852
rect 14480 10908 14544 10912
rect 14480 10852 14484 10908
rect 14484 10852 14540 10908
rect 14540 10852 14544 10908
rect 14480 10848 14544 10852
rect 14560 10908 14624 10912
rect 14560 10852 14564 10908
rect 14564 10852 14620 10908
rect 14620 10852 14624 10908
rect 14560 10848 14624 10852
rect 14640 10908 14704 10912
rect 14640 10852 14644 10908
rect 14644 10852 14700 10908
rect 14700 10852 14704 10908
rect 14640 10848 14704 10852
rect 14720 10908 14784 10912
rect 14720 10852 14724 10908
rect 14724 10852 14780 10908
rect 14780 10852 14784 10908
rect 14720 10848 14784 10852
rect 23813 10908 23877 10912
rect 23813 10852 23817 10908
rect 23817 10852 23873 10908
rect 23873 10852 23877 10908
rect 23813 10848 23877 10852
rect 23893 10908 23957 10912
rect 23893 10852 23897 10908
rect 23897 10852 23953 10908
rect 23953 10852 23957 10908
rect 23893 10848 23957 10852
rect 23973 10908 24037 10912
rect 23973 10852 23977 10908
rect 23977 10852 24033 10908
rect 24033 10852 24037 10908
rect 23973 10848 24037 10852
rect 24053 10908 24117 10912
rect 24053 10852 24057 10908
rect 24057 10852 24113 10908
rect 24113 10852 24117 10908
rect 24053 10848 24117 10852
rect 9813 10364 9877 10368
rect 9813 10308 9817 10364
rect 9817 10308 9873 10364
rect 9873 10308 9877 10364
rect 9813 10304 9877 10308
rect 9893 10364 9957 10368
rect 9893 10308 9897 10364
rect 9897 10308 9953 10364
rect 9953 10308 9957 10364
rect 9893 10304 9957 10308
rect 9973 10364 10037 10368
rect 9973 10308 9977 10364
rect 9977 10308 10033 10364
rect 10033 10308 10037 10364
rect 9973 10304 10037 10308
rect 10053 10364 10117 10368
rect 10053 10308 10057 10364
rect 10057 10308 10113 10364
rect 10113 10308 10117 10364
rect 10053 10304 10117 10308
rect 19146 10364 19210 10368
rect 19146 10308 19150 10364
rect 19150 10308 19206 10364
rect 19206 10308 19210 10364
rect 19146 10304 19210 10308
rect 19226 10364 19290 10368
rect 19226 10308 19230 10364
rect 19230 10308 19286 10364
rect 19286 10308 19290 10364
rect 19226 10304 19290 10308
rect 19306 10364 19370 10368
rect 19306 10308 19310 10364
rect 19310 10308 19366 10364
rect 19366 10308 19370 10364
rect 19306 10304 19370 10308
rect 19386 10364 19450 10368
rect 19386 10308 19390 10364
rect 19390 10308 19446 10364
rect 19446 10308 19450 10364
rect 19386 10304 19450 10308
rect 5146 9820 5210 9824
rect 5146 9764 5150 9820
rect 5150 9764 5206 9820
rect 5206 9764 5210 9820
rect 5146 9760 5210 9764
rect 5226 9820 5290 9824
rect 5226 9764 5230 9820
rect 5230 9764 5286 9820
rect 5286 9764 5290 9820
rect 5226 9760 5290 9764
rect 5306 9820 5370 9824
rect 5306 9764 5310 9820
rect 5310 9764 5366 9820
rect 5366 9764 5370 9820
rect 5306 9760 5370 9764
rect 5386 9820 5450 9824
rect 5386 9764 5390 9820
rect 5390 9764 5446 9820
rect 5446 9764 5450 9820
rect 5386 9760 5450 9764
rect 14480 9820 14544 9824
rect 14480 9764 14484 9820
rect 14484 9764 14540 9820
rect 14540 9764 14544 9820
rect 14480 9760 14544 9764
rect 14560 9820 14624 9824
rect 14560 9764 14564 9820
rect 14564 9764 14620 9820
rect 14620 9764 14624 9820
rect 14560 9760 14624 9764
rect 14640 9820 14704 9824
rect 14640 9764 14644 9820
rect 14644 9764 14700 9820
rect 14700 9764 14704 9820
rect 14640 9760 14704 9764
rect 14720 9820 14784 9824
rect 14720 9764 14724 9820
rect 14724 9764 14780 9820
rect 14780 9764 14784 9820
rect 14720 9760 14784 9764
rect 23813 9820 23877 9824
rect 23813 9764 23817 9820
rect 23817 9764 23873 9820
rect 23873 9764 23877 9820
rect 23813 9760 23877 9764
rect 23893 9820 23957 9824
rect 23893 9764 23897 9820
rect 23897 9764 23953 9820
rect 23953 9764 23957 9820
rect 23893 9760 23957 9764
rect 23973 9820 24037 9824
rect 23973 9764 23977 9820
rect 23977 9764 24033 9820
rect 24033 9764 24037 9820
rect 23973 9760 24037 9764
rect 24053 9820 24117 9824
rect 24053 9764 24057 9820
rect 24057 9764 24113 9820
rect 24113 9764 24117 9820
rect 24053 9760 24117 9764
rect 24244 9752 24308 9756
rect 24244 9696 24294 9752
rect 24294 9696 24308 9752
rect 24244 9692 24308 9696
rect 9813 9276 9877 9280
rect 9813 9220 9817 9276
rect 9817 9220 9873 9276
rect 9873 9220 9877 9276
rect 9813 9216 9877 9220
rect 9893 9276 9957 9280
rect 9893 9220 9897 9276
rect 9897 9220 9953 9276
rect 9953 9220 9957 9276
rect 9893 9216 9957 9220
rect 9973 9276 10037 9280
rect 9973 9220 9977 9276
rect 9977 9220 10033 9276
rect 10033 9220 10037 9276
rect 9973 9216 10037 9220
rect 10053 9276 10117 9280
rect 10053 9220 10057 9276
rect 10057 9220 10113 9276
rect 10113 9220 10117 9276
rect 10053 9216 10117 9220
rect 19146 9276 19210 9280
rect 19146 9220 19150 9276
rect 19150 9220 19206 9276
rect 19206 9220 19210 9276
rect 19146 9216 19210 9220
rect 19226 9276 19290 9280
rect 19226 9220 19230 9276
rect 19230 9220 19286 9276
rect 19286 9220 19290 9276
rect 19226 9216 19290 9220
rect 19306 9276 19370 9280
rect 19306 9220 19310 9276
rect 19310 9220 19366 9276
rect 19366 9220 19370 9276
rect 19306 9216 19370 9220
rect 19386 9276 19450 9280
rect 19386 9220 19390 9276
rect 19390 9220 19446 9276
rect 19446 9220 19450 9276
rect 19386 9216 19450 9220
rect 5146 8732 5210 8736
rect 5146 8676 5150 8732
rect 5150 8676 5206 8732
rect 5206 8676 5210 8732
rect 5146 8672 5210 8676
rect 5226 8732 5290 8736
rect 5226 8676 5230 8732
rect 5230 8676 5286 8732
rect 5286 8676 5290 8732
rect 5226 8672 5290 8676
rect 5306 8732 5370 8736
rect 5306 8676 5310 8732
rect 5310 8676 5366 8732
rect 5366 8676 5370 8732
rect 5306 8672 5370 8676
rect 5386 8732 5450 8736
rect 5386 8676 5390 8732
rect 5390 8676 5446 8732
rect 5446 8676 5450 8732
rect 5386 8672 5450 8676
rect 14480 8732 14544 8736
rect 14480 8676 14484 8732
rect 14484 8676 14540 8732
rect 14540 8676 14544 8732
rect 14480 8672 14544 8676
rect 14560 8732 14624 8736
rect 14560 8676 14564 8732
rect 14564 8676 14620 8732
rect 14620 8676 14624 8732
rect 14560 8672 14624 8676
rect 14640 8732 14704 8736
rect 14640 8676 14644 8732
rect 14644 8676 14700 8732
rect 14700 8676 14704 8732
rect 14640 8672 14704 8676
rect 14720 8732 14784 8736
rect 14720 8676 14724 8732
rect 14724 8676 14780 8732
rect 14780 8676 14784 8732
rect 14720 8672 14784 8676
rect 23813 8732 23877 8736
rect 23813 8676 23817 8732
rect 23817 8676 23873 8732
rect 23873 8676 23877 8732
rect 23813 8672 23877 8676
rect 23893 8732 23957 8736
rect 23893 8676 23897 8732
rect 23897 8676 23953 8732
rect 23953 8676 23957 8732
rect 23893 8672 23957 8676
rect 23973 8732 24037 8736
rect 23973 8676 23977 8732
rect 23977 8676 24033 8732
rect 24033 8676 24037 8732
rect 23973 8672 24037 8676
rect 24053 8732 24117 8736
rect 24053 8676 24057 8732
rect 24057 8676 24113 8732
rect 24113 8676 24117 8732
rect 24053 8672 24117 8676
rect 9813 8188 9877 8192
rect 9813 8132 9817 8188
rect 9817 8132 9873 8188
rect 9873 8132 9877 8188
rect 9813 8128 9877 8132
rect 9893 8188 9957 8192
rect 9893 8132 9897 8188
rect 9897 8132 9953 8188
rect 9953 8132 9957 8188
rect 9893 8128 9957 8132
rect 9973 8188 10037 8192
rect 9973 8132 9977 8188
rect 9977 8132 10033 8188
rect 10033 8132 10037 8188
rect 9973 8128 10037 8132
rect 10053 8188 10117 8192
rect 10053 8132 10057 8188
rect 10057 8132 10113 8188
rect 10113 8132 10117 8188
rect 10053 8128 10117 8132
rect 19146 8188 19210 8192
rect 19146 8132 19150 8188
rect 19150 8132 19206 8188
rect 19206 8132 19210 8188
rect 19146 8128 19210 8132
rect 19226 8188 19290 8192
rect 19226 8132 19230 8188
rect 19230 8132 19286 8188
rect 19286 8132 19290 8188
rect 19226 8128 19290 8132
rect 19306 8188 19370 8192
rect 19306 8132 19310 8188
rect 19310 8132 19366 8188
rect 19366 8132 19370 8188
rect 19306 8128 19370 8132
rect 19386 8188 19450 8192
rect 19386 8132 19390 8188
rect 19390 8132 19446 8188
rect 19446 8132 19450 8188
rect 19386 8128 19450 8132
rect 5146 7644 5210 7648
rect 5146 7588 5150 7644
rect 5150 7588 5206 7644
rect 5206 7588 5210 7644
rect 5146 7584 5210 7588
rect 5226 7644 5290 7648
rect 5226 7588 5230 7644
rect 5230 7588 5286 7644
rect 5286 7588 5290 7644
rect 5226 7584 5290 7588
rect 5306 7644 5370 7648
rect 5306 7588 5310 7644
rect 5310 7588 5366 7644
rect 5366 7588 5370 7644
rect 5306 7584 5370 7588
rect 5386 7644 5450 7648
rect 5386 7588 5390 7644
rect 5390 7588 5446 7644
rect 5446 7588 5450 7644
rect 5386 7584 5450 7588
rect 14480 7644 14544 7648
rect 14480 7588 14484 7644
rect 14484 7588 14540 7644
rect 14540 7588 14544 7644
rect 14480 7584 14544 7588
rect 14560 7644 14624 7648
rect 14560 7588 14564 7644
rect 14564 7588 14620 7644
rect 14620 7588 14624 7644
rect 14560 7584 14624 7588
rect 14640 7644 14704 7648
rect 14640 7588 14644 7644
rect 14644 7588 14700 7644
rect 14700 7588 14704 7644
rect 14640 7584 14704 7588
rect 14720 7644 14784 7648
rect 14720 7588 14724 7644
rect 14724 7588 14780 7644
rect 14780 7588 14784 7644
rect 14720 7584 14784 7588
rect 23813 7644 23877 7648
rect 23813 7588 23817 7644
rect 23817 7588 23873 7644
rect 23873 7588 23877 7644
rect 23813 7584 23877 7588
rect 23893 7644 23957 7648
rect 23893 7588 23897 7644
rect 23897 7588 23953 7644
rect 23953 7588 23957 7644
rect 23893 7584 23957 7588
rect 23973 7644 24037 7648
rect 23973 7588 23977 7644
rect 23977 7588 24033 7644
rect 24033 7588 24037 7644
rect 23973 7584 24037 7588
rect 24053 7644 24117 7648
rect 24053 7588 24057 7644
rect 24057 7588 24113 7644
rect 24113 7588 24117 7644
rect 24053 7584 24117 7588
rect 9813 7100 9877 7104
rect 9813 7044 9817 7100
rect 9817 7044 9873 7100
rect 9873 7044 9877 7100
rect 9813 7040 9877 7044
rect 9893 7100 9957 7104
rect 9893 7044 9897 7100
rect 9897 7044 9953 7100
rect 9953 7044 9957 7100
rect 9893 7040 9957 7044
rect 9973 7100 10037 7104
rect 9973 7044 9977 7100
rect 9977 7044 10033 7100
rect 10033 7044 10037 7100
rect 9973 7040 10037 7044
rect 10053 7100 10117 7104
rect 10053 7044 10057 7100
rect 10057 7044 10113 7100
rect 10113 7044 10117 7100
rect 10053 7040 10117 7044
rect 19146 7100 19210 7104
rect 19146 7044 19150 7100
rect 19150 7044 19206 7100
rect 19206 7044 19210 7100
rect 19146 7040 19210 7044
rect 19226 7100 19290 7104
rect 19226 7044 19230 7100
rect 19230 7044 19286 7100
rect 19286 7044 19290 7100
rect 19226 7040 19290 7044
rect 19306 7100 19370 7104
rect 19306 7044 19310 7100
rect 19310 7044 19366 7100
rect 19366 7044 19370 7100
rect 19306 7040 19370 7044
rect 19386 7100 19450 7104
rect 19386 7044 19390 7100
rect 19390 7044 19446 7100
rect 19446 7044 19450 7100
rect 19386 7040 19450 7044
rect 5146 6556 5210 6560
rect 5146 6500 5150 6556
rect 5150 6500 5206 6556
rect 5206 6500 5210 6556
rect 5146 6496 5210 6500
rect 5226 6556 5290 6560
rect 5226 6500 5230 6556
rect 5230 6500 5286 6556
rect 5286 6500 5290 6556
rect 5226 6496 5290 6500
rect 5306 6556 5370 6560
rect 5306 6500 5310 6556
rect 5310 6500 5366 6556
rect 5366 6500 5370 6556
rect 5306 6496 5370 6500
rect 5386 6556 5450 6560
rect 5386 6500 5390 6556
rect 5390 6500 5446 6556
rect 5446 6500 5450 6556
rect 5386 6496 5450 6500
rect 14480 6556 14544 6560
rect 14480 6500 14484 6556
rect 14484 6500 14540 6556
rect 14540 6500 14544 6556
rect 14480 6496 14544 6500
rect 14560 6556 14624 6560
rect 14560 6500 14564 6556
rect 14564 6500 14620 6556
rect 14620 6500 14624 6556
rect 14560 6496 14624 6500
rect 14640 6556 14704 6560
rect 14640 6500 14644 6556
rect 14644 6500 14700 6556
rect 14700 6500 14704 6556
rect 14640 6496 14704 6500
rect 14720 6556 14784 6560
rect 14720 6500 14724 6556
rect 14724 6500 14780 6556
rect 14780 6500 14784 6556
rect 14720 6496 14784 6500
rect 23813 6556 23877 6560
rect 23813 6500 23817 6556
rect 23817 6500 23873 6556
rect 23873 6500 23877 6556
rect 23813 6496 23877 6500
rect 23893 6556 23957 6560
rect 23893 6500 23897 6556
rect 23897 6500 23953 6556
rect 23953 6500 23957 6556
rect 23893 6496 23957 6500
rect 23973 6556 24037 6560
rect 23973 6500 23977 6556
rect 23977 6500 24033 6556
rect 24033 6500 24037 6556
rect 23973 6496 24037 6500
rect 24053 6556 24117 6560
rect 24053 6500 24057 6556
rect 24057 6500 24113 6556
rect 24113 6500 24117 6556
rect 24053 6496 24117 6500
rect 9813 6012 9877 6016
rect 9813 5956 9817 6012
rect 9817 5956 9873 6012
rect 9873 5956 9877 6012
rect 9813 5952 9877 5956
rect 9893 6012 9957 6016
rect 9893 5956 9897 6012
rect 9897 5956 9953 6012
rect 9953 5956 9957 6012
rect 9893 5952 9957 5956
rect 9973 6012 10037 6016
rect 9973 5956 9977 6012
rect 9977 5956 10033 6012
rect 10033 5956 10037 6012
rect 9973 5952 10037 5956
rect 10053 6012 10117 6016
rect 10053 5956 10057 6012
rect 10057 5956 10113 6012
rect 10113 5956 10117 6012
rect 10053 5952 10117 5956
rect 19146 6012 19210 6016
rect 19146 5956 19150 6012
rect 19150 5956 19206 6012
rect 19206 5956 19210 6012
rect 19146 5952 19210 5956
rect 19226 6012 19290 6016
rect 19226 5956 19230 6012
rect 19230 5956 19286 6012
rect 19286 5956 19290 6012
rect 19226 5952 19290 5956
rect 19306 6012 19370 6016
rect 19306 5956 19310 6012
rect 19310 5956 19366 6012
rect 19366 5956 19370 6012
rect 19306 5952 19370 5956
rect 19386 6012 19450 6016
rect 19386 5956 19390 6012
rect 19390 5956 19446 6012
rect 19446 5956 19450 6012
rect 19386 5952 19450 5956
rect 5146 5468 5210 5472
rect 5146 5412 5150 5468
rect 5150 5412 5206 5468
rect 5206 5412 5210 5468
rect 5146 5408 5210 5412
rect 5226 5468 5290 5472
rect 5226 5412 5230 5468
rect 5230 5412 5286 5468
rect 5286 5412 5290 5468
rect 5226 5408 5290 5412
rect 5306 5468 5370 5472
rect 5306 5412 5310 5468
rect 5310 5412 5366 5468
rect 5366 5412 5370 5468
rect 5306 5408 5370 5412
rect 5386 5468 5450 5472
rect 5386 5412 5390 5468
rect 5390 5412 5446 5468
rect 5446 5412 5450 5468
rect 5386 5408 5450 5412
rect 14480 5468 14544 5472
rect 14480 5412 14484 5468
rect 14484 5412 14540 5468
rect 14540 5412 14544 5468
rect 14480 5408 14544 5412
rect 14560 5468 14624 5472
rect 14560 5412 14564 5468
rect 14564 5412 14620 5468
rect 14620 5412 14624 5468
rect 14560 5408 14624 5412
rect 14640 5468 14704 5472
rect 14640 5412 14644 5468
rect 14644 5412 14700 5468
rect 14700 5412 14704 5468
rect 14640 5408 14704 5412
rect 14720 5468 14784 5472
rect 14720 5412 14724 5468
rect 14724 5412 14780 5468
rect 14780 5412 14784 5468
rect 14720 5408 14784 5412
rect 23813 5468 23877 5472
rect 23813 5412 23817 5468
rect 23817 5412 23873 5468
rect 23873 5412 23877 5468
rect 23813 5408 23877 5412
rect 23893 5468 23957 5472
rect 23893 5412 23897 5468
rect 23897 5412 23953 5468
rect 23953 5412 23957 5468
rect 23893 5408 23957 5412
rect 23973 5468 24037 5472
rect 23973 5412 23977 5468
rect 23977 5412 24033 5468
rect 24033 5412 24037 5468
rect 23973 5408 24037 5412
rect 24053 5468 24117 5472
rect 24053 5412 24057 5468
rect 24057 5412 24113 5468
rect 24113 5412 24117 5468
rect 24053 5408 24117 5412
rect 9813 4924 9877 4928
rect 9813 4868 9817 4924
rect 9817 4868 9873 4924
rect 9873 4868 9877 4924
rect 9813 4864 9877 4868
rect 9893 4924 9957 4928
rect 9893 4868 9897 4924
rect 9897 4868 9953 4924
rect 9953 4868 9957 4924
rect 9893 4864 9957 4868
rect 9973 4924 10037 4928
rect 9973 4868 9977 4924
rect 9977 4868 10033 4924
rect 10033 4868 10037 4924
rect 9973 4864 10037 4868
rect 10053 4924 10117 4928
rect 10053 4868 10057 4924
rect 10057 4868 10113 4924
rect 10113 4868 10117 4924
rect 10053 4864 10117 4868
rect 19146 4924 19210 4928
rect 19146 4868 19150 4924
rect 19150 4868 19206 4924
rect 19206 4868 19210 4924
rect 19146 4864 19210 4868
rect 19226 4924 19290 4928
rect 19226 4868 19230 4924
rect 19230 4868 19286 4924
rect 19286 4868 19290 4924
rect 19226 4864 19290 4868
rect 19306 4924 19370 4928
rect 19306 4868 19310 4924
rect 19310 4868 19366 4924
rect 19366 4868 19370 4924
rect 19306 4864 19370 4868
rect 19386 4924 19450 4928
rect 19386 4868 19390 4924
rect 19390 4868 19446 4924
rect 19446 4868 19450 4924
rect 19386 4864 19450 4868
rect 5146 4380 5210 4384
rect 5146 4324 5150 4380
rect 5150 4324 5206 4380
rect 5206 4324 5210 4380
rect 5146 4320 5210 4324
rect 5226 4380 5290 4384
rect 5226 4324 5230 4380
rect 5230 4324 5286 4380
rect 5286 4324 5290 4380
rect 5226 4320 5290 4324
rect 5306 4380 5370 4384
rect 5306 4324 5310 4380
rect 5310 4324 5366 4380
rect 5366 4324 5370 4380
rect 5306 4320 5370 4324
rect 5386 4380 5450 4384
rect 5386 4324 5390 4380
rect 5390 4324 5446 4380
rect 5446 4324 5450 4380
rect 5386 4320 5450 4324
rect 14480 4380 14544 4384
rect 14480 4324 14484 4380
rect 14484 4324 14540 4380
rect 14540 4324 14544 4380
rect 14480 4320 14544 4324
rect 14560 4380 14624 4384
rect 14560 4324 14564 4380
rect 14564 4324 14620 4380
rect 14620 4324 14624 4380
rect 14560 4320 14624 4324
rect 14640 4380 14704 4384
rect 14640 4324 14644 4380
rect 14644 4324 14700 4380
rect 14700 4324 14704 4380
rect 14640 4320 14704 4324
rect 14720 4380 14784 4384
rect 14720 4324 14724 4380
rect 14724 4324 14780 4380
rect 14780 4324 14784 4380
rect 14720 4320 14784 4324
rect 23813 4380 23877 4384
rect 23813 4324 23817 4380
rect 23817 4324 23873 4380
rect 23873 4324 23877 4380
rect 23813 4320 23877 4324
rect 23893 4380 23957 4384
rect 23893 4324 23897 4380
rect 23897 4324 23953 4380
rect 23953 4324 23957 4380
rect 23893 4320 23957 4324
rect 23973 4380 24037 4384
rect 23973 4324 23977 4380
rect 23977 4324 24033 4380
rect 24033 4324 24037 4380
rect 23973 4320 24037 4324
rect 24053 4380 24117 4384
rect 24053 4324 24057 4380
rect 24057 4324 24113 4380
rect 24113 4324 24117 4380
rect 24053 4320 24117 4324
rect 9813 3836 9877 3840
rect 9813 3780 9817 3836
rect 9817 3780 9873 3836
rect 9873 3780 9877 3836
rect 9813 3776 9877 3780
rect 9893 3836 9957 3840
rect 9893 3780 9897 3836
rect 9897 3780 9953 3836
rect 9953 3780 9957 3836
rect 9893 3776 9957 3780
rect 9973 3836 10037 3840
rect 9973 3780 9977 3836
rect 9977 3780 10033 3836
rect 10033 3780 10037 3836
rect 9973 3776 10037 3780
rect 10053 3836 10117 3840
rect 10053 3780 10057 3836
rect 10057 3780 10113 3836
rect 10113 3780 10117 3836
rect 10053 3776 10117 3780
rect 19146 3836 19210 3840
rect 19146 3780 19150 3836
rect 19150 3780 19206 3836
rect 19206 3780 19210 3836
rect 19146 3776 19210 3780
rect 19226 3836 19290 3840
rect 19226 3780 19230 3836
rect 19230 3780 19286 3836
rect 19286 3780 19290 3836
rect 19226 3776 19290 3780
rect 19306 3836 19370 3840
rect 19306 3780 19310 3836
rect 19310 3780 19366 3836
rect 19366 3780 19370 3836
rect 19306 3776 19370 3780
rect 19386 3836 19450 3840
rect 19386 3780 19390 3836
rect 19390 3780 19446 3836
rect 19446 3780 19450 3836
rect 19386 3776 19450 3780
rect 5146 3292 5210 3296
rect 5146 3236 5150 3292
rect 5150 3236 5206 3292
rect 5206 3236 5210 3292
rect 5146 3232 5210 3236
rect 5226 3292 5290 3296
rect 5226 3236 5230 3292
rect 5230 3236 5286 3292
rect 5286 3236 5290 3292
rect 5226 3232 5290 3236
rect 5306 3292 5370 3296
rect 5306 3236 5310 3292
rect 5310 3236 5366 3292
rect 5366 3236 5370 3292
rect 5306 3232 5370 3236
rect 5386 3292 5450 3296
rect 5386 3236 5390 3292
rect 5390 3236 5446 3292
rect 5446 3236 5450 3292
rect 5386 3232 5450 3236
rect 14480 3292 14544 3296
rect 14480 3236 14484 3292
rect 14484 3236 14540 3292
rect 14540 3236 14544 3292
rect 14480 3232 14544 3236
rect 14560 3292 14624 3296
rect 14560 3236 14564 3292
rect 14564 3236 14620 3292
rect 14620 3236 14624 3292
rect 14560 3232 14624 3236
rect 14640 3292 14704 3296
rect 14640 3236 14644 3292
rect 14644 3236 14700 3292
rect 14700 3236 14704 3292
rect 14640 3232 14704 3236
rect 14720 3292 14784 3296
rect 14720 3236 14724 3292
rect 14724 3236 14780 3292
rect 14780 3236 14784 3292
rect 14720 3232 14784 3236
rect 23813 3292 23877 3296
rect 23813 3236 23817 3292
rect 23817 3236 23873 3292
rect 23873 3236 23877 3292
rect 23813 3232 23877 3236
rect 23893 3292 23957 3296
rect 23893 3236 23897 3292
rect 23897 3236 23953 3292
rect 23953 3236 23957 3292
rect 23893 3232 23957 3236
rect 23973 3292 24037 3296
rect 23973 3236 23977 3292
rect 23977 3236 24033 3292
rect 24033 3236 24037 3292
rect 23973 3232 24037 3236
rect 24053 3292 24117 3296
rect 24053 3236 24057 3292
rect 24057 3236 24113 3292
rect 24113 3236 24117 3292
rect 24053 3232 24117 3236
rect 9813 2748 9877 2752
rect 9813 2692 9817 2748
rect 9817 2692 9873 2748
rect 9873 2692 9877 2748
rect 9813 2688 9877 2692
rect 9893 2748 9957 2752
rect 9893 2692 9897 2748
rect 9897 2692 9953 2748
rect 9953 2692 9957 2748
rect 9893 2688 9957 2692
rect 9973 2748 10037 2752
rect 9973 2692 9977 2748
rect 9977 2692 10033 2748
rect 10033 2692 10037 2748
rect 9973 2688 10037 2692
rect 10053 2748 10117 2752
rect 10053 2692 10057 2748
rect 10057 2692 10113 2748
rect 10113 2692 10117 2748
rect 10053 2688 10117 2692
rect 19146 2748 19210 2752
rect 19146 2692 19150 2748
rect 19150 2692 19206 2748
rect 19206 2692 19210 2748
rect 19146 2688 19210 2692
rect 19226 2748 19290 2752
rect 19226 2692 19230 2748
rect 19230 2692 19286 2748
rect 19286 2692 19290 2748
rect 19226 2688 19290 2692
rect 19306 2748 19370 2752
rect 19306 2692 19310 2748
rect 19310 2692 19366 2748
rect 19366 2692 19370 2748
rect 19306 2688 19370 2692
rect 19386 2748 19450 2752
rect 19386 2692 19390 2748
rect 19390 2692 19446 2748
rect 19446 2692 19450 2748
rect 19386 2688 19450 2692
rect 5146 2204 5210 2208
rect 5146 2148 5150 2204
rect 5150 2148 5206 2204
rect 5206 2148 5210 2204
rect 5146 2144 5210 2148
rect 5226 2204 5290 2208
rect 5226 2148 5230 2204
rect 5230 2148 5286 2204
rect 5286 2148 5290 2204
rect 5226 2144 5290 2148
rect 5306 2204 5370 2208
rect 5306 2148 5310 2204
rect 5310 2148 5366 2204
rect 5366 2148 5370 2204
rect 5306 2144 5370 2148
rect 5386 2204 5450 2208
rect 5386 2148 5390 2204
rect 5390 2148 5446 2204
rect 5446 2148 5450 2204
rect 5386 2144 5450 2148
rect 14480 2204 14544 2208
rect 14480 2148 14484 2204
rect 14484 2148 14540 2204
rect 14540 2148 14544 2204
rect 14480 2144 14544 2148
rect 14560 2204 14624 2208
rect 14560 2148 14564 2204
rect 14564 2148 14620 2204
rect 14620 2148 14624 2204
rect 14560 2144 14624 2148
rect 14640 2204 14704 2208
rect 14640 2148 14644 2204
rect 14644 2148 14700 2204
rect 14700 2148 14704 2204
rect 14640 2144 14704 2148
rect 14720 2204 14784 2208
rect 14720 2148 14724 2204
rect 14724 2148 14780 2204
rect 14780 2148 14784 2204
rect 14720 2144 14784 2148
rect 23813 2204 23877 2208
rect 23813 2148 23817 2204
rect 23817 2148 23873 2204
rect 23873 2148 23877 2204
rect 23813 2144 23877 2148
rect 23893 2204 23957 2208
rect 23893 2148 23897 2204
rect 23897 2148 23953 2204
rect 23953 2148 23957 2204
rect 23893 2144 23957 2148
rect 23973 2204 24037 2208
rect 23973 2148 23977 2204
rect 23977 2148 24033 2204
rect 24033 2148 24037 2204
rect 23973 2144 24037 2148
rect 24053 2204 24117 2208
rect 24053 2148 24057 2204
rect 24057 2148 24113 2204
rect 24113 2148 24117 2204
rect 24053 2144 24117 2148
<< metal4 >>
rect 5138 25056 5459 25616
rect 5138 24992 5146 25056
rect 5210 24992 5226 25056
rect 5290 24992 5306 25056
rect 5370 24992 5386 25056
rect 5450 24992 5459 25056
rect 5138 23968 5459 24992
rect 5138 23904 5146 23968
rect 5210 23904 5226 23968
rect 5290 23904 5306 23968
rect 5370 23904 5386 23968
rect 5450 23904 5459 23968
rect 5138 22880 5459 23904
rect 5138 22816 5146 22880
rect 5210 22816 5226 22880
rect 5290 22816 5306 22880
rect 5370 22816 5386 22880
rect 5450 22816 5459 22880
rect 5138 21792 5459 22816
rect 5138 21728 5146 21792
rect 5210 21728 5226 21792
rect 5290 21728 5306 21792
rect 5370 21728 5386 21792
rect 5450 21728 5459 21792
rect 5138 20704 5459 21728
rect 5138 20640 5146 20704
rect 5210 20640 5226 20704
rect 5290 20640 5306 20704
rect 5370 20640 5386 20704
rect 5450 20640 5459 20704
rect 5138 19616 5459 20640
rect 5138 19552 5146 19616
rect 5210 19552 5226 19616
rect 5290 19552 5306 19616
rect 5370 19552 5386 19616
rect 5450 19552 5459 19616
rect 5138 18528 5459 19552
rect 5138 18464 5146 18528
rect 5210 18464 5226 18528
rect 5290 18464 5306 18528
rect 5370 18464 5386 18528
rect 5450 18464 5459 18528
rect 5138 17440 5459 18464
rect 5138 17376 5146 17440
rect 5210 17376 5226 17440
rect 5290 17376 5306 17440
rect 5370 17376 5386 17440
rect 5450 17376 5459 17440
rect 5138 16352 5459 17376
rect 5138 16288 5146 16352
rect 5210 16288 5226 16352
rect 5290 16288 5306 16352
rect 5370 16288 5386 16352
rect 5450 16288 5459 16352
rect 5138 15264 5459 16288
rect 5138 15200 5146 15264
rect 5210 15200 5226 15264
rect 5290 15200 5306 15264
rect 5370 15200 5386 15264
rect 5450 15200 5459 15264
rect 5138 14176 5459 15200
rect 5138 14112 5146 14176
rect 5210 14112 5226 14176
rect 5290 14112 5306 14176
rect 5370 14112 5386 14176
rect 5450 14112 5459 14176
rect 5138 13088 5459 14112
rect 5138 13024 5146 13088
rect 5210 13024 5226 13088
rect 5290 13024 5306 13088
rect 5370 13024 5386 13088
rect 5450 13024 5459 13088
rect 5138 12000 5459 13024
rect 5138 11936 5146 12000
rect 5210 11936 5226 12000
rect 5290 11936 5306 12000
rect 5370 11936 5386 12000
rect 5450 11936 5459 12000
rect 5138 10912 5459 11936
rect 5138 10848 5146 10912
rect 5210 10848 5226 10912
rect 5290 10848 5306 10912
rect 5370 10848 5386 10912
rect 5450 10848 5459 10912
rect 5138 9824 5459 10848
rect 5138 9760 5146 9824
rect 5210 9760 5226 9824
rect 5290 9760 5306 9824
rect 5370 9760 5386 9824
rect 5450 9760 5459 9824
rect 5138 8736 5459 9760
rect 5138 8672 5146 8736
rect 5210 8672 5226 8736
rect 5290 8672 5306 8736
rect 5370 8672 5386 8736
rect 5450 8672 5459 8736
rect 5138 7648 5459 8672
rect 5138 7584 5146 7648
rect 5210 7584 5226 7648
rect 5290 7584 5306 7648
rect 5370 7584 5386 7648
rect 5450 7584 5459 7648
rect 5138 6560 5459 7584
rect 5138 6496 5146 6560
rect 5210 6496 5226 6560
rect 5290 6496 5306 6560
rect 5370 6496 5386 6560
rect 5450 6496 5459 6560
rect 5138 5472 5459 6496
rect 5138 5408 5146 5472
rect 5210 5408 5226 5472
rect 5290 5408 5306 5472
rect 5370 5408 5386 5472
rect 5450 5408 5459 5472
rect 5138 4384 5459 5408
rect 5138 4320 5146 4384
rect 5210 4320 5226 4384
rect 5290 4320 5306 4384
rect 5370 4320 5386 4384
rect 5450 4320 5459 4384
rect 5138 3296 5459 4320
rect 5138 3232 5146 3296
rect 5210 3232 5226 3296
rect 5290 3232 5306 3296
rect 5370 3232 5386 3296
rect 5450 3232 5459 3296
rect 5138 2208 5459 3232
rect 5138 2144 5146 2208
rect 5210 2144 5226 2208
rect 5290 2144 5306 2208
rect 5370 2144 5386 2208
rect 5450 2144 5459 2208
rect 5138 2128 5459 2144
rect 9805 25600 10125 25616
rect 9805 25536 9813 25600
rect 9877 25536 9893 25600
rect 9957 25536 9973 25600
rect 10037 25536 10053 25600
rect 10117 25536 10125 25600
rect 9805 24512 10125 25536
rect 9805 24448 9813 24512
rect 9877 24448 9893 24512
rect 9957 24448 9973 24512
rect 10037 24448 10053 24512
rect 10117 24448 10125 24512
rect 9805 23424 10125 24448
rect 9805 23360 9813 23424
rect 9877 23360 9893 23424
rect 9957 23360 9973 23424
rect 10037 23360 10053 23424
rect 10117 23360 10125 23424
rect 9805 22336 10125 23360
rect 9805 22272 9813 22336
rect 9877 22272 9893 22336
rect 9957 22272 9973 22336
rect 10037 22272 10053 22336
rect 10117 22272 10125 22336
rect 9805 21248 10125 22272
rect 9805 21184 9813 21248
rect 9877 21184 9893 21248
rect 9957 21184 9973 21248
rect 10037 21184 10053 21248
rect 10117 21184 10125 21248
rect 9805 20160 10125 21184
rect 9805 20096 9813 20160
rect 9877 20096 9893 20160
rect 9957 20096 9973 20160
rect 10037 20096 10053 20160
rect 10117 20096 10125 20160
rect 9805 19072 10125 20096
rect 9805 19008 9813 19072
rect 9877 19008 9893 19072
rect 9957 19008 9973 19072
rect 10037 19008 10053 19072
rect 10117 19008 10125 19072
rect 9805 17984 10125 19008
rect 9805 17920 9813 17984
rect 9877 17920 9893 17984
rect 9957 17920 9973 17984
rect 10037 17920 10053 17984
rect 10117 17920 10125 17984
rect 9805 16896 10125 17920
rect 9805 16832 9813 16896
rect 9877 16832 9893 16896
rect 9957 16832 9973 16896
rect 10037 16832 10053 16896
rect 10117 16832 10125 16896
rect 9805 15808 10125 16832
rect 9805 15744 9813 15808
rect 9877 15744 9893 15808
rect 9957 15744 9973 15808
rect 10037 15744 10053 15808
rect 10117 15744 10125 15808
rect 9805 14720 10125 15744
rect 9805 14656 9813 14720
rect 9877 14656 9893 14720
rect 9957 14656 9973 14720
rect 10037 14656 10053 14720
rect 10117 14656 10125 14720
rect 9805 13632 10125 14656
rect 9805 13568 9813 13632
rect 9877 13568 9893 13632
rect 9957 13568 9973 13632
rect 10037 13568 10053 13632
rect 10117 13568 10125 13632
rect 9805 12544 10125 13568
rect 9805 12480 9813 12544
rect 9877 12480 9893 12544
rect 9957 12480 9973 12544
rect 10037 12480 10053 12544
rect 10117 12480 10125 12544
rect 9805 11456 10125 12480
rect 9805 11392 9813 11456
rect 9877 11392 9893 11456
rect 9957 11392 9973 11456
rect 10037 11392 10053 11456
rect 10117 11392 10125 11456
rect 9805 10368 10125 11392
rect 9805 10304 9813 10368
rect 9877 10304 9893 10368
rect 9957 10304 9973 10368
rect 10037 10304 10053 10368
rect 10117 10304 10125 10368
rect 9805 9280 10125 10304
rect 9805 9216 9813 9280
rect 9877 9216 9893 9280
rect 9957 9216 9973 9280
rect 10037 9216 10053 9280
rect 10117 9216 10125 9280
rect 9805 8192 10125 9216
rect 9805 8128 9813 8192
rect 9877 8128 9893 8192
rect 9957 8128 9973 8192
rect 10037 8128 10053 8192
rect 10117 8128 10125 8192
rect 9805 7104 10125 8128
rect 9805 7040 9813 7104
rect 9877 7040 9893 7104
rect 9957 7040 9973 7104
rect 10037 7040 10053 7104
rect 10117 7040 10125 7104
rect 9805 6016 10125 7040
rect 9805 5952 9813 6016
rect 9877 5952 9893 6016
rect 9957 5952 9973 6016
rect 10037 5952 10053 6016
rect 10117 5952 10125 6016
rect 9805 4928 10125 5952
rect 9805 4864 9813 4928
rect 9877 4864 9893 4928
rect 9957 4864 9973 4928
rect 10037 4864 10053 4928
rect 10117 4864 10125 4928
rect 9805 3840 10125 4864
rect 9805 3776 9813 3840
rect 9877 3776 9893 3840
rect 9957 3776 9973 3840
rect 10037 3776 10053 3840
rect 10117 3776 10125 3840
rect 9805 2752 10125 3776
rect 9805 2688 9813 2752
rect 9877 2688 9893 2752
rect 9957 2688 9973 2752
rect 10037 2688 10053 2752
rect 10117 2688 10125 2752
rect 9805 2128 10125 2688
rect 14472 25056 14792 25616
rect 14472 24992 14480 25056
rect 14544 24992 14560 25056
rect 14624 24992 14640 25056
rect 14704 24992 14720 25056
rect 14784 24992 14792 25056
rect 14472 23968 14792 24992
rect 14472 23904 14480 23968
rect 14544 23904 14560 23968
rect 14624 23904 14640 23968
rect 14704 23904 14720 23968
rect 14784 23904 14792 23968
rect 14472 22880 14792 23904
rect 14472 22816 14480 22880
rect 14544 22816 14560 22880
rect 14624 22816 14640 22880
rect 14704 22816 14720 22880
rect 14784 22816 14792 22880
rect 14472 21792 14792 22816
rect 14472 21728 14480 21792
rect 14544 21728 14560 21792
rect 14624 21728 14640 21792
rect 14704 21728 14720 21792
rect 14784 21728 14792 21792
rect 14472 20704 14792 21728
rect 14472 20640 14480 20704
rect 14544 20640 14560 20704
rect 14624 20640 14640 20704
rect 14704 20640 14720 20704
rect 14784 20640 14792 20704
rect 14472 19616 14792 20640
rect 14472 19552 14480 19616
rect 14544 19552 14560 19616
rect 14624 19552 14640 19616
rect 14704 19552 14720 19616
rect 14784 19552 14792 19616
rect 14472 18528 14792 19552
rect 14472 18464 14480 18528
rect 14544 18464 14560 18528
rect 14624 18464 14640 18528
rect 14704 18464 14720 18528
rect 14784 18464 14792 18528
rect 14472 17440 14792 18464
rect 14472 17376 14480 17440
rect 14544 17376 14560 17440
rect 14624 17376 14640 17440
rect 14704 17376 14720 17440
rect 14784 17376 14792 17440
rect 14472 16352 14792 17376
rect 14472 16288 14480 16352
rect 14544 16288 14560 16352
rect 14624 16288 14640 16352
rect 14704 16288 14720 16352
rect 14784 16288 14792 16352
rect 14472 15264 14792 16288
rect 14472 15200 14480 15264
rect 14544 15200 14560 15264
rect 14624 15200 14640 15264
rect 14704 15200 14720 15264
rect 14784 15200 14792 15264
rect 14472 14176 14792 15200
rect 14472 14112 14480 14176
rect 14544 14112 14560 14176
rect 14624 14112 14640 14176
rect 14704 14112 14720 14176
rect 14784 14112 14792 14176
rect 14472 13088 14792 14112
rect 14472 13024 14480 13088
rect 14544 13024 14560 13088
rect 14624 13024 14640 13088
rect 14704 13024 14720 13088
rect 14784 13024 14792 13088
rect 14472 12000 14792 13024
rect 14472 11936 14480 12000
rect 14544 11936 14560 12000
rect 14624 11936 14640 12000
rect 14704 11936 14720 12000
rect 14784 11936 14792 12000
rect 14472 10912 14792 11936
rect 14472 10848 14480 10912
rect 14544 10848 14560 10912
rect 14624 10848 14640 10912
rect 14704 10848 14720 10912
rect 14784 10848 14792 10912
rect 14472 9824 14792 10848
rect 14472 9760 14480 9824
rect 14544 9760 14560 9824
rect 14624 9760 14640 9824
rect 14704 9760 14720 9824
rect 14784 9760 14792 9824
rect 14472 8736 14792 9760
rect 14472 8672 14480 8736
rect 14544 8672 14560 8736
rect 14624 8672 14640 8736
rect 14704 8672 14720 8736
rect 14784 8672 14792 8736
rect 14472 7648 14792 8672
rect 14472 7584 14480 7648
rect 14544 7584 14560 7648
rect 14624 7584 14640 7648
rect 14704 7584 14720 7648
rect 14784 7584 14792 7648
rect 14472 6560 14792 7584
rect 14472 6496 14480 6560
rect 14544 6496 14560 6560
rect 14624 6496 14640 6560
rect 14704 6496 14720 6560
rect 14784 6496 14792 6560
rect 14472 5472 14792 6496
rect 14472 5408 14480 5472
rect 14544 5408 14560 5472
rect 14624 5408 14640 5472
rect 14704 5408 14720 5472
rect 14784 5408 14792 5472
rect 14472 4384 14792 5408
rect 14472 4320 14480 4384
rect 14544 4320 14560 4384
rect 14624 4320 14640 4384
rect 14704 4320 14720 4384
rect 14784 4320 14792 4384
rect 14472 3296 14792 4320
rect 14472 3232 14480 3296
rect 14544 3232 14560 3296
rect 14624 3232 14640 3296
rect 14704 3232 14720 3296
rect 14784 3232 14792 3296
rect 14472 2208 14792 3232
rect 14472 2144 14480 2208
rect 14544 2144 14560 2208
rect 14624 2144 14640 2208
rect 14704 2144 14720 2208
rect 14784 2144 14792 2208
rect 14472 2128 14792 2144
rect 19138 25600 19458 25616
rect 19138 25536 19146 25600
rect 19210 25536 19226 25600
rect 19290 25536 19306 25600
rect 19370 25536 19386 25600
rect 19450 25536 19458 25600
rect 19138 24512 19458 25536
rect 19138 24448 19146 24512
rect 19210 24448 19226 24512
rect 19290 24448 19306 24512
rect 19370 24448 19386 24512
rect 19450 24448 19458 24512
rect 19138 23424 19458 24448
rect 19138 23360 19146 23424
rect 19210 23360 19226 23424
rect 19290 23360 19306 23424
rect 19370 23360 19386 23424
rect 19450 23360 19458 23424
rect 19138 22336 19458 23360
rect 19138 22272 19146 22336
rect 19210 22272 19226 22336
rect 19290 22272 19306 22336
rect 19370 22272 19386 22336
rect 19450 22272 19458 22336
rect 19138 21248 19458 22272
rect 19138 21184 19146 21248
rect 19210 21184 19226 21248
rect 19290 21184 19306 21248
rect 19370 21184 19386 21248
rect 19450 21184 19458 21248
rect 19138 20160 19458 21184
rect 19138 20096 19146 20160
rect 19210 20096 19226 20160
rect 19290 20096 19306 20160
rect 19370 20096 19386 20160
rect 19450 20096 19458 20160
rect 19138 19072 19458 20096
rect 19138 19008 19146 19072
rect 19210 19008 19226 19072
rect 19290 19008 19306 19072
rect 19370 19008 19386 19072
rect 19450 19008 19458 19072
rect 19138 17984 19458 19008
rect 19138 17920 19146 17984
rect 19210 17920 19226 17984
rect 19290 17920 19306 17984
rect 19370 17920 19386 17984
rect 19450 17920 19458 17984
rect 19138 16896 19458 17920
rect 19138 16832 19146 16896
rect 19210 16832 19226 16896
rect 19290 16832 19306 16896
rect 19370 16832 19386 16896
rect 19450 16832 19458 16896
rect 19138 15808 19458 16832
rect 19138 15744 19146 15808
rect 19210 15744 19226 15808
rect 19290 15744 19306 15808
rect 19370 15744 19386 15808
rect 19450 15744 19458 15808
rect 19138 14720 19458 15744
rect 19138 14656 19146 14720
rect 19210 14656 19226 14720
rect 19290 14656 19306 14720
rect 19370 14656 19386 14720
rect 19450 14656 19458 14720
rect 19138 13632 19458 14656
rect 19138 13568 19146 13632
rect 19210 13568 19226 13632
rect 19290 13568 19306 13632
rect 19370 13568 19386 13632
rect 19450 13568 19458 13632
rect 19138 12544 19458 13568
rect 19138 12480 19146 12544
rect 19210 12480 19226 12544
rect 19290 12480 19306 12544
rect 19370 12480 19386 12544
rect 19450 12480 19458 12544
rect 19138 11456 19458 12480
rect 19138 11392 19146 11456
rect 19210 11392 19226 11456
rect 19290 11392 19306 11456
rect 19370 11392 19386 11456
rect 19450 11392 19458 11456
rect 19138 10368 19458 11392
rect 19138 10304 19146 10368
rect 19210 10304 19226 10368
rect 19290 10304 19306 10368
rect 19370 10304 19386 10368
rect 19450 10304 19458 10368
rect 19138 9280 19458 10304
rect 19138 9216 19146 9280
rect 19210 9216 19226 9280
rect 19290 9216 19306 9280
rect 19370 9216 19386 9280
rect 19450 9216 19458 9280
rect 19138 8192 19458 9216
rect 19138 8128 19146 8192
rect 19210 8128 19226 8192
rect 19290 8128 19306 8192
rect 19370 8128 19386 8192
rect 19450 8128 19458 8192
rect 19138 7104 19458 8128
rect 19138 7040 19146 7104
rect 19210 7040 19226 7104
rect 19290 7040 19306 7104
rect 19370 7040 19386 7104
rect 19450 7040 19458 7104
rect 19138 6016 19458 7040
rect 19138 5952 19146 6016
rect 19210 5952 19226 6016
rect 19290 5952 19306 6016
rect 19370 5952 19386 6016
rect 19450 5952 19458 6016
rect 19138 4928 19458 5952
rect 19138 4864 19146 4928
rect 19210 4864 19226 4928
rect 19290 4864 19306 4928
rect 19370 4864 19386 4928
rect 19450 4864 19458 4928
rect 19138 3840 19458 4864
rect 19138 3776 19146 3840
rect 19210 3776 19226 3840
rect 19290 3776 19306 3840
rect 19370 3776 19386 3840
rect 19450 3776 19458 3840
rect 19138 2752 19458 3776
rect 19138 2688 19146 2752
rect 19210 2688 19226 2752
rect 19290 2688 19306 2752
rect 19370 2688 19386 2752
rect 19450 2688 19458 2752
rect 19138 2128 19458 2688
rect 23805 25056 24125 25616
rect 23805 24992 23813 25056
rect 23877 24992 23893 25056
rect 23957 24992 23973 25056
rect 24037 24992 24053 25056
rect 24117 24992 24125 25056
rect 23805 23968 24125 24992
rect 23805 23904 23813 23968
rect 23877 23904 23893 23968
rect 23957 23904 23973 23968
rect 24037 23904 24053 23968
rect 24117 23904 24125 23968
rect 23805 22880 24125 23904
rect 23805 22816 23813 22880
rect 23877 22816 23893 22880
rect 23957 22816 23973 22880
rect 24037 22816 24053 22880
rect 24117 22816 24125 22880
rect 23805 21792 24125 22816
rect 23805 21728 23813 21792
rect 23877 21728 23893 21792
rect 23957 21728 23973 21792
rect 24037 21728 24053 21792
rect 24117 21728 24125 21792
rect 23805 20704 24125 21728
rect 23805 20640 23813 20704
rect 23877 20640 23893 20704
rect 23957 20640 23973 20704
rect 24037 20640 24053 20704
rect 24117 20640 24125 20704
rect 23805 19616 24125 20640
rect 23805 19552 23813 19616
rect 23877 19552 23893 19616
rect 23957 19552 23973 19616
rect 24037 19552 24053 19616
rect 24117 19552 24125 19616
rect 23805 18528 24125 19552
rect 23805 18464 23813 18528
rect 23877 18464 23893 18528
rect 23957 18464 23973 18528
rect 24037 18464 24053 18528
rect 24117 18464 24125 18528
rect 23805 17440 24125 18464
rect 23805 17376 23813 17440
rect 23877 17376 23893 17440
rect 23957 17376 23973 17440
rect 24037 17376 24053 17440
rect 24117 17376 24125 17440
rect 23805 16352 24125 17376
rect 23805 16288 23813 16352
rect 23877 16288 23893 16352
rect 23957 16288 23973 16352
rect 24037 16288 24053 16352
rect 24117 16288 24125 16352
rect 23805 15264 24125 16288
rect 23805 15200 23813 15264
rect 23877 15200 23893 15264
rect 23957 15200 23973 15264
rect 24037 15200 24053 15264
rect 24117 15200 24125 15264
rect 23805 14176 24125 15200
rect 23805 14112 23813 14176
rect 23877 14112 23893 14176
rect 23957 14112 23973 14176
rect 24037 14112 24053 14176
rect 24117 14112 24125 14176
rect 23805 13088 24125 14112
rect 24243 13972 24309 13973
rect 24243 13908 24244 13972
rect 24308 13908 24309 13972
rect 24243 13907 24309 13908
rect 23805 13024 23813 13088
rect 23877 13024 23893 13088
rect 23957 13024 23973 13088
rect 24037 13024 24053 13088
rect 24117 13024 24125 13088
rect 23805 12000 24125 13024
rect 23805 11936 23813 12000
rect 23877 11936 23893 12000
rect 23957 11936 23973 12000
rect 24037 11936 24053 12000
rect 24117 11936 24125 12000
rect 23805 10912 24125 11936
rect 23805 10848 23813 10912
rect 23877 10848 23893 10912
rect 23957 10848 23973 10912
rect 24037 10848 24053 10912
rect 24117 10848 24125 10912
rect 23805 9824 24125 10848
rect 23805 9760 23813 9824
rect 23877 9760 23893 9824
rect 23957 9760 23973 9824
rect 24037 9760 24053 9824
rect 24117 9760 24125 9824
rect 23805 8736 24125 9760
rect 24246 9757 24306 13907
rect 24243 9756 24309 9757
rect 24243 9692 24244 9756
rect 24308 9692 24309 9756
rect 24243 9691 24309 9692
rect 23805 8672 23813 8736
rect 23877 8672 23893 8736
rect 23957 8672 23973 8736
rect 24037 8672 24053 8736
rect 24117 8672 24125 8736
rect 23805 7648 24125 8672
rect 23805 7584 23813 7648
rect 23877 7584 23893 7648
rect 23957 7584 23973 7648
rect 24037 7584 24053 7648
rect 24117 7584 24125 7648
rect 23805 6560 24125 7584
rect 23805 6496 23813 6560
rect 23877 6496 23893 6560
rect 23957 6496 23973 6560
rect 24037 6496 24053 6560
rect 24117 6496 24125 6560
rect 23805 5472 24125 6496
rect 23805 5408 23813 5472
rect 23877 5408 23893 5472
rect 23957 5408 23973 5472
rect 24037 5408 24053 5472
rect 24117 5408 24125 5472
rect 23805 4384 24125 5408
rect 23805 4320 23813 4384
rect 23877 4320 23893 4384
rect 23957 4320 23973 4384
rect 24037 4320 24053 4384
rect 24117 4320 24125 4384
rect 23805 3296 24125 4320
rect 23805 3232 23813 3296
rect 23877 3232 23893 3296
rect 23957 3232 23973 3296
rect 24037 3232 24053 3296
rect 24117 3232 24125 3296
rect 23805 2208 24125 3232
rect 23805 2144 23813 2208
rect 23877 2144 23893 2208
rect 23957 2144 23973 2208
rect 24037 2144 24053 2208
rect 24117 2144 24125 2208
rect 23805 2128 24125 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 632 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 632 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 908 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 908 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3116 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2012 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3116 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3484 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 3576 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4220 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 4680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5324 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6336 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6244 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5784 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6428 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6060 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6336 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 7532 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7440 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9188 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 8636 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9280 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 8544 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 9648 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 10752 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12040 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 11856 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11488 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 11948 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12132 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13052 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14340 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14156 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 14892 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 14984 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_159
timestamp 1586364061
transform 1 0 15260 0 1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16180 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16088 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_167
timestamp 1586364061
transform 1 0 15996 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16364 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 17744 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17468 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17192 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 17836 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 17560 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 18940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 18664 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20596 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20044 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 20688 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 19768 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 20872 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 21792 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 21976 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23448 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23080 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 22896 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 23540 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23172 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24092 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24368 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 24736 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24276 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 25840 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25380 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26392 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26392 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 632 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 908 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2012 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3116 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3484 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 3576 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 4680 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 5784 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 6888 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 7992 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9096 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9188 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10292 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11396 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12500 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 13604 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 14708 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 14800 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_166
timestamp 1586364061
transform 1 0 15904 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16180 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_172
timestamp 1586364061
transform 1 0 16456 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_184
timestamp 1586364061
transform 1 0 17560 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_196
timestamp 1586364061
transform 1 0 18664 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20320 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_208
timestamp 1586364061
transform 1 0 19768 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20412 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21516 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 22620 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 23724 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 25932 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 24828 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26024 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26392 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 632 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 908 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2012 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3116 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4220 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5324 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6244 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6060 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6336 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7440 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 8544 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 9648 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 10752 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 11856 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 11948 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13052 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_147
timestamp 1586364061
transform 1 0 14156 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _197_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15076 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 14892 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_166
timestamp 1586364061
transform 1 0 15904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16088 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_170
timestamp 1586364061
transform 1 0 16272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_174
timestamp 1586364061
transform 1 0 16640 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17468 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17376 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 17560 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 18756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_196
timestamp 1586364061
transform 1 0 18664 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_199
timestamp 1586364061
transform 1 0 18940 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_211
timestamp 1586364061
transform 1 0 20044 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_223
timestamp 1586364061
transform 1 0 21148 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_235
timestamp 1586364061
transform 1 0 22252 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23080 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 22988 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23172 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 23908 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_262
timestamp 1586364061
transform 1 0 24736 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24920 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_266
timestamp 1586364061
transform 1 0 25104 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 25840 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26392 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 632 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 908 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2012 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3116 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3484 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 3576 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 4680 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 5784 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 6888 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 7992 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9096 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9188 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10292 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11396 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12500 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 13604 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15720 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 14708 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14984 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 14800 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_158
timestamp 1586364061
transform 1 0 15168 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_173
timestamp 1586364061
transform 1 0 16548 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17560 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_181
timestamp 1586364061
transform 1 0 17284 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_186
timestamp 1586364061
transform 1 0 17744 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 18756 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_194
timestamp 1586364061
transform 1 0 18480 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 19584 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20320 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20412 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21516 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 22620 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_251
timestamp 1586364061
transform 1 0 23724 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_258
timestamp 1586364061
transform 1 0 24368 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 25932 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25472 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 25840 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26024 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26392 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 632 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 908 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2012 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3116 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4220 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5324 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6244 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6060 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6336 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7440 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 8544 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 9648 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 10752 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 11856 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 11948 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13052 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 13788 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_147
timestamp 1586364061
transform 1 0 14156 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_151
timestamp 1586364061
transform 1 0 14524 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14892 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14708 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_164
timestamp 1586364061
transform 1 0 15720 0 1 4896
box -38 -48 590 592
use scs8hd_conb_1  _215_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16456 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16916 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 16732 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17100 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17468 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18388 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19492 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19308 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 18572 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18940 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 18756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_201
timestamp 1586364061
transform 1 0 19124 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20504 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20872 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20320 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 20688 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_222
timestamp 1586364061
transform 1 0 21056 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_234
timestamp 1586364061
transform 1 0 22160 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23080 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 22896 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_245
timestamp 1586364061
transform 1 0 23172 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_249
timestamp 1586364061
transform 1 0 23540 0 1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_262
timestamp 1586364061
transform 1 0 24736 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24920 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_266
timestamp 1586364061
transform 1 0 25104 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_274
timestamp 1586364061
transform 1 0 25840 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26392 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 632 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 632 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 908 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 908 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2012 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3116 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2012 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3116 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3484 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 3576 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4220 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 4680 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5324 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6244 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 5784 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 6888 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6060 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6336 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 7992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7440 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9096 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9188 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 8544 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10292 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 9648 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_110
timestamp 1586364061
transform 1 0 10752 0 1 5984
box -38 -48 406 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 11948 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 11856 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 11580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 11212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 11948 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_117
timestamp 1586364061
transform 1 0 11396 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_114
timestamp 1586364061
transform 1 0 11120 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_117
timestamp 1586364061
transform 1 0 11396 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 11764 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 13144 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_125
timestamp 1586364061
transform 1 0 12132 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_137
timestamp 1586364061
transform 1 0 13236 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 12776 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13328 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 14432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 13512 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_149
timestamp 1586364061
transform 1 0 14340 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_142
timestamp 1586364061
transform 1 0 13696 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 14616 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14800 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15352 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 14708 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15168 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 14800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_165
timestamp 1586364061
transform 1 0 15812 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 14984 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16548 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 16548 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 16916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_171
timestamp 1586364061
transform 1 0 16364 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 16732 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17100 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 18112 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17560 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17468 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17284 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17560 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17376 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_186
timestamp 1586364061
transform 1 0 17744 0 -1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19308 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19124 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19308 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_199
timestamp 1586364061
transform 1 0 18940 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_205
timestamp 1586364061
transform 1 0 19492 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 18572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 18940 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20412 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20320 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20872 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20504 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20228 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_214
timestamp 1586364061
transform 1 0 20320 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 20688 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21056 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 22068 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_224
timestamp 1586364061
transform 1 0 21240 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 21884 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_235
timestamp 1586364061
transform 1 0 22252 0 1 5984
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23080 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23172 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23080 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22896 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_236
timestamp 1586364061
transform 1 0 22344 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_247
timestamp 1586364061
transform 1 0 23356 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_241
timestamp 1586364061
transform 1 0 22804 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_248
timestamp 1586364061
transform 1 0 23448 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24184 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24644 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23816 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24368 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24000 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24460 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 25932 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25012 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25472 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 25840 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26024 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_263
timestamp 1586364061
transform 1 0 24828 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_267
timestamp 1586364061
transform 1 0 25196 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 25932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26392 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26392 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 632 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 908 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2012 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3116 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3484 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 3576 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 4680 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 5784 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 6888 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 7992 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9096 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9188 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10292 0 -1 7072
box -38 -48 1142 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11580 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_117
timestamp 1586364061
transform 1 0 11396 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _156_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13144 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_128
timestamp 1586364061
transform 1 0 12408 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 14156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 13972 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14340 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 14800 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 14708 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15812 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_163
timestamp 1586364061
transform 1 0 15628 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 16364 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_167
timestamp 1586364061
transform 1 0 15996 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_180
timestamp 1586364061
transform 1 0 17192 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_192
timestamp 1586364061
transform 1 0 18296 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18664 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18480 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19492 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 20412 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20320 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20228 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 21516 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_224
timestamp 1586364061
transform 1 0 21240 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_229
timestamp 1586364061
transform 1 0 21700 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 22804 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 23264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_244
timestamp 1586364061
transform 1 0 23080 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_248
timestamp 1586364061
transform 1 0 23448 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23816 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_255
timestamp 1586364061
transform 1 0 24092 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24828 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 25932 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_266
timestamp 1586364061
transform 1 0 25104 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 25840 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26024 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26392 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 632 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 908 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3116 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4220 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5324 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6244 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6060 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6336 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7440 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 8544 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 9648 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_110
timestamp 1586364061
transform 1 0 10752 0 1 7072
box -38 -48 774 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12040 0 1 7072
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 11856 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 11672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11488 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_123
timestamp 1586364061
transform 1 0 11948 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 12868 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 13236 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 12684 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_135
timestamp 1586364061
transform 1 0 13052 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _153_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13788 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 13604 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_139
timestamp 1586364061
transform 1 0 13420 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 14616 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 15352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 15168 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 14800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 14984 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 16364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 16732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_169
timestamp 1586364061
transform 1 0 16180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 16548 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_177
timestamp 1586364061
transform 1 0 16916 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 17744 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17468 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 17284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 17560 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19124 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_195
timestamp 1586364061
transform 1 0 18572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 18940 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_203
timestamp 1586364061
transform 1 0 19308 0 1 7072
box -38 -48 774 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 20136 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_211
timestamp 1586364061
transform 1 0 20044 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_215
timestamp 1586364061
transform 1 0 20412 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 21516 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21148 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 23172 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23080 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22344 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 22712 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _231_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24736 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 24552 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_254
timestamp 1586364061
transform 1 0 24000 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25288 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25104 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25472 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26024 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26392 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 632 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 908 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2012 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3116 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3484 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 3576 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 4680 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 5784 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 6888 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 7992 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9096 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9188 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10292 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11396 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 13144 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_129
timestamp 1586364061
transform 1 0 12500 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_135
timestamp 1586364061
transform 1 0 13052 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_138
timestamp 1586364061
transform 1 0 13328 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 13696 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 14064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_144
timestamp 1586364061
transform 1 0 13880 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_148
timestamp 1586364061
transform 1 0 14248 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 14616 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 15904 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 14708 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 15352 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 15720 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_154
timestamp 1586364061
transform 1 0 14800 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_162
timestamp 1586364061
transform 1 0 15536 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16916 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_175
timestamp 1586364061
transform 1 0 16732 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_179
timestamp 1586364061
transform 1 0 17100 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18388 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17560 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18204 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_183
timestamp 1586364061
transform 1 0 17468 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_186
timestamp 1586364061
transform 1 0 17744 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_190
timestamp 1586364061
transform 1 0 18112 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19216 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20320 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_215
timestamp 1586364061
transform 1 0 20412 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21424 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  FILLER_10_223
timestamp 1586364061
transform 1 0 21148 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_235
timestamp 1586364061
transform 1 0 22252 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22988 0 -1 8160
box -38 -48 866 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24552 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_252
timestamp 1586364061
transform 1 0 23816 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 25932 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_264
timestamp 1586364061
transform 1 0 24920 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 25656 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26024 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26392 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 632 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 908 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2012 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4220 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5324 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6244 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6060 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6336 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7440 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 8544 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 9648 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 10752 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 11856 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_123
timestamp 1586364061
transform 1 0 11948 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 13144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 12776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_131
timestamp 1586364061
transform 1 0 12684 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 12960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13328 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 13696 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 13512 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_151
timestamp 1586364061
transform 1 0 14524 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 15904 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 15720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 14984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 15352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_155
timestamp 1586364061
transform 1 0 14892 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 15536 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16916 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 16732 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17100 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17560 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17468 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17284 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19308 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19124 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 18572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 18940 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20688 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20320 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_212
timestamp 1586364061
transform 1 0 20136 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20504 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_220
timestamp 1586364061
transform 1 0 20872 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21332 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21148 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23080 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22344 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 22712 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 24736 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24184 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 24552 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25288 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_266
timestamp 1586364061
transform 1 0 25104 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_270
timestamp 1586364061
transform 1 0 25472 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26024 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26392 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 632 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 908 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2012 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3116 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3484 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 3576 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 4680 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 5784 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 6888 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 7992 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9096 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9188 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10292 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_117
timestamp 1586364061
transform 1 0 11396 0 -1 9248
box -38 -48 774 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 13144 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 12316 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12132 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_129
timestamp 1586364061
transform 1 0 12500 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_135
timestamp 1586364061
transform 1 0 13052 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 14524 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 14156 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 13972 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14340 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 14984 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 14708 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 14800 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 15812 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16548 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 15996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 16364 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_169
timestamp 1586364061
transform 1 0 16180 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18296 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_184
timestamp 1586364061
transform 1 0 17560 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19308 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19124 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19492 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20688 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20320 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20228 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_215
timestamp 1586364061
transform 1 0 20412 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21884 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_229
timestamp 1586364061
transform 1 0 21700 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_233
timestamp 1586364061
transform 1 0 22068 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22896 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22528 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_237
timestamp 1586364061
transform 1 0 22436 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_240
timestamp 1586364061
transform 1 0 22712 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 24460 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23908 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_251
timestamp 1586364061
transform 1 0 23724 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_255
timestamp 1586364061
transform 1 0 24092 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 25932 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 24828 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26024 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26392 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 632 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 632 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 908 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 908 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2012 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3116 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2012 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3116 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3484 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4220 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 3576 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5324 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 4680 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6244 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6060 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6336 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 5784 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 6888 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7440 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 7992 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9096 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 8544 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9188 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 9648 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 10752 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10292 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 11856 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 11948 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11396 0 -1 10336
box -38 -48 1142 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 12316 0 1 9248
box -38 -48 682 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 13144 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 13144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 12132 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 12960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13328 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_129
timestamp 1586364061
transform 1 0 12500 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_135
timestamp 1586364061
transform 1 0 13052 0 -1 10336
box -38 -48 130 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 13696 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 13512 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 14524 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 14156 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_151
timestamp 1586364061
transform 1 0 14524 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 13972 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14340 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 15260 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 14800 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 14708 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 15076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 14708 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 15812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_155
timestamp 1586364061
transform 1 0 14892 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 15628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 16272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 16640 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 16180 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_168
timestamp 1586364061
transform 1 0 16088 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16456 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_176
timestamp 1586364061
transform 1 0 16824 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_167
timestamp 1586364061
transform 1 0 15996 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_171
timestamp 1586364061
transform 1 0 16364 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17468 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 18296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17928 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17376 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_184
timestamp 1586364061
transform 1 0 17560 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_190
timestamp 1586364061
transform 1 0 18112 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_183
timestamp 1586364061
transform 1 0 17468 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 18664 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18848 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18664 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_194
timestamp 1586364061
transform 1 0 18480 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_207
timestamp 1586364061
transform 1 0 19676 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_195
timestamp 1586364061
transform 1 0 18572 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19492 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 20412 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 20412 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20320 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 20872 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_218
timestamp 1586364061
transform 1 0 20688 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20228 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22068 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 21240 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_222
timestamp 1586364061
transform 1 0 21056 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_226
timestamp 1586364061
transform 1 0 21424 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 21976 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_224
timestamp 1586364061
transform 1 0 21240 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_241
timestamp 1586364061
transform 1 0 22804 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_236
timestamp 1586364061
transform 1 0 22344 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 22712 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22344 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22528 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22896 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22528 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_247
timestamp 1586364061
transform 1 0 23356 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 23172 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23080 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23540 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 23172 0 1 9248
box -38 -48 866 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 24736 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24552 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24000 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_258
timestamp 1586364061
transform 1 0 24368 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_258
timestamp 1586364061
transform 1 0 24368 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_262
timestamp 1586364061
transform 1 0 24736 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 25932 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25288 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_266
timestamp 1586364061
transform 1 0 25104 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_270
timestamp 1586364061
transform 1 0 25472 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26024 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 25840 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26024 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26392 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26392 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 632 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 908 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2012 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3116 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4220 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5324 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6244 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6060 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6336 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7440 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 8544 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 9648 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 10752 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 11856 0 1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_15_123
timestamp 1586364061
transform 1 0 11948 0 1 10336
box -38 -48 590 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 13052 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 12868 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 12500 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_131
timestamp 1586364061
transform 1 0 12684 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _122_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14616 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 14064 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 14432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 13880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14248 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 15812 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 15076 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 15628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_155
timestamp 1586364061
transform 1 0 14892 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_159
timestamp 1586364061
transform 1 0 15260 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 16640 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_178
timestamp 1586364061
transform 1 0 17008 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17468 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18112 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17744 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17376 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 17560 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 17928 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_192
timestamp 1586364061
transform 1 0 18296 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 18664 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 19676 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 18480 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_205
timestamp 1586364061
transform 1 0 19492 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 20228 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 20044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_209
timestamp 1586364061
transform 1 0 19860 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 22068 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21792 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_222
timestamp 1586364061
transform 1 0 21056 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_232
timestamp 1586364061
transform 1 0 21976 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23356 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23080 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 22712 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_245
timestamp 1586364061
transform 1 0 23172 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24736 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_256
timestamp 1586364061
transform 1 0 24184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_260
timestamp 1586364061
transform 1 0 24552 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 24920 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 25472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25288 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_272
timestamp 1586364061
transform 1 0 25656 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26024 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26392 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 632 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 908 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2012 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3116 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3484 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 3576 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 4680 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 5784 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 6888 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 7992 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9096 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9188 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10292 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11396 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 12500 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_132
timestamp 1586364061
transform 1 0 12776 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 13512 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 13972 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 14340 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_143
timestamp 1586364061
transform 1 0 13788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_147
timestamp 1586364061
transform 1 0 14156 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14524 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 14800 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 14708 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 15812 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 15628 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16364 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_16_167
timestamp 1586364061
transform 1 0 15996 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18112 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17560 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17928 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17376 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 17744 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19308 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_199
timestamp 1586364061
transform 1 0 18940 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_205
timestamp 1586364061
transform 1 0 19492 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20320 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 20596 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20228 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20412 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_219
timestamp 1586364061
transform 1 0 20780 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21792 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21332 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_227
timestamp 1586364061
transform 1 0 21516 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23540 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23172 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_241
timestamp 1586364061
transform 1 0 22804 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_247
timestamp 1586364061
transform 1 0 23356 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_258
timestamp 1586364061
transform 1 0 24368 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 25932 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25472 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 25840 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26024 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26392 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 632 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 908 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2012 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5324 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6244 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6060 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6336 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7440 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 8544 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 9648 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 10752 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 11856 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_123
timestamp 1586364061
transform 1 0 11948 0 1 11424
box -38 -48 774 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 12868 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 13328 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 12684 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13144 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 13880 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 13696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13512 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 15444 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 15260 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 14892 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 14708 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15076 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 16456 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16916 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_170
timestamp 1586364061
transform 1 0 16272 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_174
timestamp 1586364061
transform 1 0 16640 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17100 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17560 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17468 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17284 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19308 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19124 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_195
timestamp 1586364061
transform 1 0 18572 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 20504 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_212
timestamp 1586364061
transform 1 0 20136 0 1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_17_218
timestamp 1586364061
transform 1 0 20688 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21332 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_222
timestamp 1586364061
transform 1 0 21056 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23080 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 22528 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22344 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 22712 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_254
timestamp 1586364061
transform 1 0 24000 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_266
timestamp 1586364061
transform 1 0 25104 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 25840 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26392 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 632 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 908 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2012 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3116 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3484 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 3576 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 4680 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 5784 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 6888 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 7992 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9096 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9188 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10292 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11396 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 12684 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 13144 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_129
timestamp 1586364061
transform 1 0 12500 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_134
timestamp 1586364061
transform 1 0 12960 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13328 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 13696 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 14156 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 14524 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 13512 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 13972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14340 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 14800 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 14708 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 15444 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 15812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_157
timestamp 1586364061
transform 1 0 15076 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 15628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 16180 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 15996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_171
timestamp 1586364061
transform 1 0 16364 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_179
timestamp 1586364061
transform 1 0 17100 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17284 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_18_190
timestamp 1586364061
transform 1 0 18112 0 -1 12512
box -38 -48 590 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 19124 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19584 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18664 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_198
timestamp 1586364061
transform 1 0 18848 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_204
timestamp 1586364061
transform 1 0 19400 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 20504 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20320 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_208
timestamp 1586364061
transform 1 0 19768 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_215
timestamp 1586364061
transform 1 0 20412 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 21516 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_225
timestamp 1586364061
transform 1 0 21332 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_229
timestamp 1586364061
transform 1 0 21700 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 22712 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_237
timestamp 1586364061
transform 1 0 22436 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_249
timestamp 1586364061
transform 1 0 23540 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_261
timestamp 1586364061
transform 1 0 24644 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 25932 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_273
timestamp 1586364061
transform 1 0 25748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26024 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26392 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 632 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 632 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 908 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 908 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2012 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3116 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3116 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3484 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4220 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 3576 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5324 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 4680 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6244 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6060 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6336 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 5784 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 6888 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7440 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 7992 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9096 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 8544 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9188 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 9648 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 10752 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10292 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 11856 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 11948 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_117
timestamp 1586364061
transform 1 0 11396 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_20_128
timestamp 1586364061
transform 1 0 12408 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_131
timestamp 1586364061
transform 1 0 12684 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_127
timestamp 1586364061
transform 1 0 12316 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 12132 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 12132 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13328 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 12960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 12960 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 12776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 13144 0 1 12512
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 13144 0 -1 13600
box -38 -48 866 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 13696 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 13512 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 14156 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 14524 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_151
timestamp 1586364061
transform 1 0 14524 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 13972 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14340 0 -1 13600
box -38 -48 222 592
use scs8hd_nor3_4  _168_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14800 0 -1 13600
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15628 0 1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 14708 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15444 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 14800 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_156
timestamp 1586364061
transform 1 0 14984 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_160
timestamp 1586364061
transform 1 0 15352 0 1 12512
box -38 -48 130 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 17100 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 16916 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16180 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_174
timestamp 1586364061
transform 1 0 16640 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17100 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_167
timestamp 1586364061
transform 1 0 15996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_171
timestamp 1586364061
transform 1 0 16364 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 17560 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17468 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 17284 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_193
timestamp 1586364061
transform 1 0 18388 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_188
timestamp 1586364061
transform 1 0 17928 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19216 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18664 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19032 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18664 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_198
timestamp 1586364061
transform 1 0 18848 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_205
timestamp 1586364061
transform 1 0 19492 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 20596 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 20780 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20320 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 20596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 20228 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_211
timestamp 1586364061
transform 1 0 20044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_215
timestamp 1586364061
transform 1 0 20412 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20228 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20412 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22160 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 21976 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 21792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22160 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_228
timestamp 1586364061
transform 1 0 21608 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_232
timestamp 1586364061
transform 1 0 21976 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_226
timestamp 1586364061
transform 1 0 21424 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23080 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23356 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22896 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_236
timestamp 1586364061
transform 1 0 22344 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23172 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_249
timestamp 1586364061
transform 1 0 23540 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_237
timestamp 1586364061
transform 1 0 22436 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 24736 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23632 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24092 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 24736 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 23908 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_257
timestamp 1586364061
transform 1 0 24276 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_261
timestamp 1586364061
transform 1 0 24644 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_254
timestamp 1586364061
transform 1 0 24000 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 25932 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_264
timestamp 1586364061
transform 1 0 24920 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26024 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25104 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 25840 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26024 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26392 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26392 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 632 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 908 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2012 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3116 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4220 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5324 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6244 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6060 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6336 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7440 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 8544 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 9648 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 10752 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 11856 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_123
timestamp 1586364061
transform 1 0 11948 0 1 13600
box -38 -48 774 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 12960 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_131
timestamp 1586364061
transform 1 0 12684 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13236 0 1 13600
box -38 -48 222 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 14340 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 14156 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13420 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 13788 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_141
timestamp 1586364061
transform 1 0 13604 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 13972 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 15720 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 15536 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_166
timestamp 1586364061
transform 1 0 15904 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 16088 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 16456 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16272 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_174
timestamp 1586364061
transform 1 0 16640 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17468 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17744 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18112 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17376 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_184
timestamp 1586364061
transform 1 0 17560 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_188
timestamp 1586364061
transform 1 0 17928 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_192
timestamp 1586364061
transform 1 0 18296 0 1 13600
box -38 -48 590 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 19032 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 18848 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20780 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_209
timestamp 1586364061
transform 1 0 19860 0 1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_21_217
timestamp 1586364061
transform 1 0 20596 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_221
timestamp 1586364061
transform 1 0 20964 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21332 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21148 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23080 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 22528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 22712 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 24736 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 24184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24000 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24368 0 1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_21_265
timestamp 1586364061
transform 1 0 25012 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26392 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 632 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 908 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2012 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3116 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3484 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 3576 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 4680 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 5784 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 6888 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 7992 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9096 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9188 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10292 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11396 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12500 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 14340 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 13972 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_141
timestamp 1586364061
transform 1 0 13604 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_147
timestamp 1586364061
transform 1 0 14156 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_151
timestamp 1586364061
transform 1 0 14524 0 -1 14688
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 14800 0 -1 14688
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 14708 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16640 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_167
timestamp 1586364061
transform 1 0 15996 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_173
timestamp 1586364061
transform 1 0 16548 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_176
timestamp 1586364061
transform 1 0 16824 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17744 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17560 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19124 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_197
timestamp 1586364061
transform 1 0 18756 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_203
timestamp 1586364061
transform 1 0 19308 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20412 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20320 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20044 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 21976 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21424 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21240 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_228
timestamp 1586364061
transform 1 0 21608 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 23540 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23172 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_241
timestamp 1586364061
transform 1 0 22804 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_247
timestamp 1586364061
transform 1 0 23356 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_258
timestamp 1586364061
transform 1 0 24368 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 25932 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_270
timestamp 1586364061
transform 1 0 25472 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 25840 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26024 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26392 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 632 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 908 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2012 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3116 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4220 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5324 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6244 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6060 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6336 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7440 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 8544 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 9648 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 10752 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 11856 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 11948 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13052 0 1 14688
box -38 -48 774 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 14340 0 1 14688
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 14156 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 13788 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 13972 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 15536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 15904 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 16272 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17100 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16088 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_173
timestamp 1586364061
transform 1 0 16548 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_177
timestamp 1586364061
transform 1 0 16916 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17468 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_181
timestamp 1586364061
transform 1 0 17284 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18388 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19124 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18572 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18940 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 18756 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20964 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20780 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_210
timestamp 1586364061
transform 1 0 19952 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_218
timestamp 1586364061
transform 1 0 20688 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22160 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_232
timestamp 1586364061
transform 1 0 21976 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23080 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 23356 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22344 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_240
timestamp 1586364061
transform 1 0 22712 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23172 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_249
timestamp 1586364061
transform 1 0 23540 0 1 14688
box -38 -48 406 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 24092 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 23908 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_259
timestamp 1586364061
transform 1 0 24460 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24828 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_265
timestamp 1586364061
transform 1 0 25012 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26392 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 632 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 908 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2012 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3116 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3484 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 3576 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 4680 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 5784 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 6888 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 7992 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9096 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9188 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10292 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11396 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 13144 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_129
timestamp 1586364061
transform 1 0 12500 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13052 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_138
timestamp 1586364061
transform 1 0 13328 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 14064 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 14432 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_148
timestamp 1586364061
transform 1 0 14248 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 14616 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14892 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 14708 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_154
timestamp 1586364061
transform 1 0 14800 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_166
timestamp 1586364061
transform 1 0 15904 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16640 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16088 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16456 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_170
timestamp 1586364061
transform 1 0 16272 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18388 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 17836 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18204 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_185
timestamp 1586364061
transform 1 0 17652 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_189
timestamp 1586364061
transform 1 0 18020 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19400 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_202
timestamp 1586364061
transform 1 0 19216 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 19584 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 20412 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20320 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20964 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_218
timestamp 1586364061
transform 1 0 20688 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21700 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_223
timestamp 1586364061
transform 1 0 21148 0 -1 15776
box -38 -48 590 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 23264 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_238
timestamp 1586364061
transform 1 0 22528 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_255
timestamp 1586364061
transform 1 0 24092 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24828 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 25932 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_266
timestamp 1586364061
transform 1 0 25104 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 25840 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26024 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26392 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 632 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 908 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2012 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3116 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4220 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5324 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6244 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6060 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6336 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7440 0 1 15776
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 9464 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_86
timestamp 1586364061
transform 1 0 8544 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_94
timestamp 1586364061
transform 1 0 9280 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 9924 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10292 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 10660 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_99
timestamp 1586364061
transform 1 0 9740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_103
timestamp 1586364061
transform 1 0 10108 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_107
timestamp 1586364061
transform 1 0 10476 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 11856 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 11488 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_111
timestamp 1586364061
transform 1 0 10844 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_117
timestamp 1586364061
transform 1 0 11396 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 11672 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 11948 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 13144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 12776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 12408 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_127
timestamp 1586364061
transform 1 0 12316 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 12592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 12960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13328 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 14064 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 13880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 13512 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_142
timestamp 1586364061
transform 1 0 13696 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 15904 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 15076 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 15444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_155
timestamp 1586364061
transform 1 0 14892 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_159
timestamp 1586364061
transform 1 0 15260 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_163
timestamp 1586364061
transform 1 0 15628 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 16916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 16732 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17100 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 17836 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17468 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 17284 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_184
timestamp 1586364061
transform 1 0 17560 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19400 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19216 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18848 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_196
timestamp 1586364061
transform 1 0 18664 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_200
timestamp 1586364061
transform 1 0 19032 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 20596 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 20964 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_213
timestamp 1586364061
transform 1 0 20228 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_219
timestamp 1586364061
transform 1 0 20780 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_223
timestamp 1586364061
transform 1 0 21148 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_235
timestamp 1586364061
transform 1 0 22252 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23080 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 22712 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 24736 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24000 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_258
timestamp 1586364061
transform 1 0 24368 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 25288 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25104 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_270
timestamp 1586364061
transform 1 0 25472 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26024 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26392 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 632 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 632 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 908 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 908 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2012 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3116 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2012 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3116 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3484 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 3576 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4220 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 4680 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5324 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6244 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 5784 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 6888 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6060 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6336 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_80
timestamp 1586364061
transform 1 0 7992 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_27_74
timestamp 1586364061
transform 1 0 7440 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_82
timestamp 1586364061
transform 1 0 8176 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 8544 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9096 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 8360 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 8544 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9464 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 8728 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9188 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_95
timestamp 1586364061
transform 1 0 9372 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 9924 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10108 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_98
timestamp 1586364061
transform 1 0 9648 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_110
timestamp 1586364061
transform 1 0 10752 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 9740 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 11488 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 11856 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11488 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11304 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_114
timestamp 1586364061
transform 1 0 11120 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 11672 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_123
timestamp 1586364061
transform 1 0 11948 0 1 16864
box -38 -48 314 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 13144 0 -1 16864
box -38 -48 866 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 12776 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 12592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 12224 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 12776 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_127
timestamp 1586364061
transform 1 0 12316 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_131
timestamp 1586364061
transform 1 0 12684 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_134
timestamp 1586364061
transform 1 0 12960 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_128
timestamp 1586364061
transform 1 0 12408 0 1 16864
box -38 -48 222 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 14340 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 13788 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 14156 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 14340 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_145
timestamp 1586364061
transform 1 0 13972 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14524 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_141
timestamp 1586364061
transform 1 0 13604 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_145
timestamp 1586364061
transform 1 0 13972 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15168 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_157
timestamp 1586364061
transform 1 0 15076 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 15260 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 14708 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 14800 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 15536 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_165
timestamp 1586364061
transform 1 0 15812 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_161
timestamp 1586364061
transform 1 0 15444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 15628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 15720 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 15352 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15904 0 -1 16864
box -38 -48 866 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 15904 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 16916 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_175
timestamp 1586364061
transform 1 0 16732 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 16732 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17100 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 17468 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17468 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_192
timestamp 1586364061
transform 1 0 18296 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_193
timestamp 1586364061
transform 1 0 18388 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 19124 0 1 16864
box -38 -48 314 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 19032 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 19584 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 18664 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 18664 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_198
timestamp 1586364061
transform 1 0 18848 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_203
timestamp 1586364061
transform 1 0 19308 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_198
timestamp 1586364061
transform 1 0 18848 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_204
timestamp 1586364061
transform 1 0 19400 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 20596 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 20596 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20320 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 20412 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 20044 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20044 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20412 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_208
timestamp 1586364061
transform 1 0 19768 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_213
timestamp 1586364061
transform 1 0 20228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21976 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 21608 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_226
timestamp 1586364061
transform 1 0 21424 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_226
timestamp 1586364061
transform 1 0 21424 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_230
timestamp 1586364061
transform 1 0 21792 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_234
timestamp 1586364061
transform 1 0 22160 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_238
timestamp 1586364061
transform 1 0 22528 0 1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_26_238
timestamp 1586364061
transform 1 0 22528 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22344 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 22896 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_245
timestamp 1586364061
transform 1 0 23172 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_248
timestamp 1586364061
transform 1 0 23448 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_244
timestamp 1586364061
transform 1 0 23080 0 -1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23080 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23172 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 23356 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24184 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23632 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24000 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_252
timestamp 1586364061
transform 1 0 23816 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_259
timestamp 1586364061
transform 1 0 24460 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_256
timestamp 1586364061
transform 1 0 24184 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_260
timestamp 1586364061
transform 1 0 24552 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24920 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 25932 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_271
timestamp 1586364061
transform 1 0 25564 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26024 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_267
timestamp 1586364061
transform 1 0 25196 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_271
timestamp 1586364061
transform 1 0 25564 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26392 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26392 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 632 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 908 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2012 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3116 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3484 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 3576 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 4680 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 5784 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 6888 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 7992 0 -1 17952
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9464 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9096 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_93
timestamp 1586364061
transform 1 0 9188 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_107
timestamp 1586364061
transform 1 0 10476 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11488 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_6  FILLER_28_111
timestamp 1586364061
transform 1 0 10844 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_117
timestamp 1586364061
transform 1 0 11396 0 -1 17952
box -38 -48 130 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 13144 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 12960 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 12592 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_127
timestamp 1586364061
transform 1 0 12316 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_132
timestamp 1586364061
transform 1 0 12776 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 14156 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 14524 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 13972 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_149
timestamp 1586364061
transform 1 0 14340 0 -1 17952
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 14800 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 14708 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 15904 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 15628 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 16364 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 16824 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_168
timestamp 1586364061
transform 1 0 16088 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_174
timestamp 1586364061
transform 1 0 16640 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_178
timestamp 1586364061
transform 1 0 17008 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17560 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_186
timestamp 1586364061
transform 1 0 17744 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 18664 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19676 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_194
timestamp 1586364061
transform 1 0 18480 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_205
timestamp 1586364061
transform 1 0 19492 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 20412 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20320 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 20136 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_209
timestamp 1586364061
transform 1 0 19860 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21976 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 21424 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21240 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 21608 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23448 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_243
timestamp 1586364061
transform 1 0 22988 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_247
timestamp 1586364061
transform 1 0 23356 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23724 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_28_250
timestamp 1586364061
transform 1 0 23632 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_260
timestamp 1586364061
transform 1 0 24552 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 25932 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_272
timestamp 1586364061
transform 1 0 25656 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26024 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26392 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 632 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 908 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2012 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5324 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6244 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6060 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6336 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7440 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 8728 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 8544 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10292 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10108 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9740 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 9556 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 9924 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11948 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 11856 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11672 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11304 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11488 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 13328 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 12960 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 12776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13144 0 1 17952
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 13512 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 14524 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_149
timestamp 1586364061
transform 1 0 14340 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 15812 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 14892 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 15260 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_153
timestamp 1586364061
transform 1 0 14708 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15076 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_161
timestamp 1586364061
transform 1 0 15444 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 16180 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 16548 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_167
timestamp 1586364061
transform 1 0 15996 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_171
timestamp 1586364061
transform 1 0 16364 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_175
timestamp 1586364061
transform 1 0 16732 0 1 17952
box -38 -48 774 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 18204 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17468 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 18020 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_184
timestamp 1586364061
transform 1 0 17560 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_188
timestamp 1586364061
transform 1 0 17928 0 1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19216 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19032 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 18664 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_194
timestamp 1586364061
transform 1 0 18480 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_198
timestamp 1586364061
transform 1 0 18848 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 20412 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 20780 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_213
timestamp 1586364061
transform 1 0 20228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_217
timestamp 1586364061
transform 1 0 20596 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_221
timestamp 1586364061
transform 1 0 20964 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21332 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21148 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23080 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22896 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22344 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 22712 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_245
timestamp 1586364061
transform 1 0 23172 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_249
timestamp 1586364061
transform 1 0 23540 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23816 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23632 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_261
timestamp 1586364061
transform 1 0 24644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_273
timestamp 1586364061
transform 1 0 25748 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26392 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 632 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 908 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2012 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3116 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3484 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 3576 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 4680 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 5784 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 6888 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 7992 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9096 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 9464 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_93
timestamp 1586364061
transform 1 0 9188 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9740 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10752 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_98
timestamp 1586364061
transform 1 0 9648 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_108
timestamp 1586364061
transform 1 0 10568 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 11304 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 11948 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_112
timestamp 1586364061
transform 1 0 10936 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_119
timestamp 1586364061
transform 1 0 11580 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 13144 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12316 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12132 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_129
timestamp 1586364061
transform 1 0 12500 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_135
timestamp 1586364061
transform 1 0 13052 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_138
timestamp 1586364061
transform 1 0 13328 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 13512 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 13880 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 14524 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_142
timestamp 1586364061
transform 1 0 13696 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_146
timestamp 1586364061
transform 1 0 14064 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_150
timestamp 1586364061
transform 1 0 14432 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 15812 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 14708 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 15260 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 15628 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_154
timestamp 1586364061
transform 1 0 14800 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_158
timestamp 1586364061
transform 1 0 15168 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_161
timestamp 1586364061
transform 1 0 15444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_174
timestamp 1586364061
transform 1 0 16640 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 17744 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17560 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_182
timestamp 1586364061
transform 1 0 17376 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_189
timestamp 1586364061
transform 1 0 18020 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 18756 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_30_206
timestamp 1586364061
transform 1 0 19584 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 20412 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20320 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19768 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_210
timestamp 1586364061
transform 1 0 19952 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21424 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21240 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_228
timestamp 1586364061
transform 1 0 21608 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23448 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23264 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_240
timestamp 1586364061
transform 1 0 22712 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_30_257
timestamp 1586364061
transform 1 0 24276 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 25932 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_269
timestamp 1586364061
transform 1 0 25380 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26024 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26392 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 632 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 908 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2012 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3116 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4220 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5324 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6244 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6060 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6336 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7440 0 1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9280 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 9096 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 8728 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_86
timestamp 1586364061
transform 1 0 8544 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_90
timestamp 1586364061
transform 1 0 8912 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 10292 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 10752 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_103
timestamp 1586364061
transform 1 0 10108 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_107
timestamp 1586364061
transform 1 0 10476 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 11948 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 11856 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11488 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 11120 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_112
timestamp 1586364061
transform 1 0 10936 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_116
timestamp 1586364061
transform 1 0 11304 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 11672 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 13144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_132
timestamp 1586364061
transform 1 0 12776 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13328 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 13512 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 14524 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_149
timestamp 1586364061
transform 1 0 14340 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 15260 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 14892 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_153
timestamp 1586364061
transform 1 0 14708 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_157
timestamp 1586364061
transform 1 0 15076 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16456 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16824 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_168
timestamp 1586364061
transform 1 0 16088 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_174
timestamp 1586364061
transform 1 0 16640 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_178
timestamp 1586364061
transform 1 0 17008 0 1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17560 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17468 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17284 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19584 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 18756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_195
timestamp 1586364061
transform 1 0 18572 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_199
timestamp 1586364061
transform 1 0 18940 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_205
timestamp 1586364061
transform 1 0 19492 0 1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19768 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20964 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_219
timestamp 1586364061
transform 1 0 20780 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 22068 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21516 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21884 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_223
timestamp 1586364061
transform 1 0 21148 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_229
timestamp 1586364061
transform 1 0 21700 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23264 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23080 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 22528 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22344 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 22712 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_245
timestamp 1586364061
transform 1 0 23172 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_255
timestamp 1586364061
transform 1 0 24092 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24828 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25288 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_266
timestamp 1586364061
transform 1 0 25104 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_270
timestamp 1586364061
transform 1 0 25472 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 25840 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26392 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 632 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 908 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2012 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3116 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3484 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 3576 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 4680 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 5784 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 6888 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 7992 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 9464 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9096 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_93
timestamp 1586364061
transform 1 0 9188 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10292 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 11488 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_117
timestamp 1586364061
transform 1 0 11396 0 -1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 13144 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12500 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_127
timestamp 1586364061
transform 1 0 12316 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_131
timestamp 1586364061
transform 1 0 12684 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_135
timestamp 1586364061
transform 1 0 13052 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 14524 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_145
timestamp 1586364061
transform 1 0 13972 0 -1 20128
box -38 -48 590 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 14892 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 14708 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_154
timestamp 1586364061
transform 1 0 14800 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_164
timestamp 1586364061
transform 1 0 15720 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16456 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17652 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_183
timestamp 1586364061
transform 1 0 17468 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_187
timestamp 1586364061
transform 1 0 17836 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_193
timestamp 1586364061
transform 1 0 18388 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 18664 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18480 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_205
timestamp 1586364061
transform 1 0 19492 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20412 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20320 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20228 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_218
timestamp 1586364061
transform 1 0 20688 0 -1 20128
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21516 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21240 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_226
timestamp 1586364061
transform 1 0 21424 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 23264 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_238
timestamp 1586364061
transform 1 0 22528 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_255
timestamp 1586364061
transform 1 0 24092 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24828 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 25932 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_266
timestamp 1586364061
transform 1 0 25104 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 25840 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26024 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26392 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 632 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 632 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 908 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 908 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2012 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2012 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3116 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3484 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4220 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 3576 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5324 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 4680 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6244 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6060 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6336 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 5784 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_68
timestamp 1586364061
transform 1 0 6888 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 7532 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 7532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8084 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7348 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_74
timestamp 1586364061
transform 1 0 7440 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_77
timestamp 1586364061
transform 1 0 7716 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_83
timestamp 1586364061
transform 1 0 8268 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_72
timestamp 1586364061
transform 1 0 7256 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9004 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9280 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9096 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8820 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8452 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8912 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_87
timestamp 1586364061
transform 1 0 8636 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_84
timestamp 1586364061
transform 1 0 8360 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_93
timestamp 1586364061
transform 1 0 9188 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10200 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_102
timestamp 1586364061
transform 1 0 10016 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_106
timestamp 1586364061
transform 1 0 10384 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_105
timestamp 1586364061
transform 1 0 10292 0 -1 21216
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11304 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11948 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 11856 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11672 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11304 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10936 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11120 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11488 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_113
timestamp 1586364061
transform 1 0 11028 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_134
timestamp 1586364061
transform 1 0 12960 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_127
timestamp 1586364061
transform 1 0 12316 0 -1 21216
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13972 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13788 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13512 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13972 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_142
timestamp 1586364061
transform 1 0 13696 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_139
timestamp 1586364061
transform 1 0 13420 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_142
timestamp 1586364061
transform 1 0 13696 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_147
timestamp 1586364061
transform 1 0 14156 0 -1 21216
box -38 -48 590 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 14800 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15720 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 14708 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15536 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 15168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15812 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 14984 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15352 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_163
timestamp 1586364061
transform 1 0 15628 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16364 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16916 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 16732 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17100 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_167
timestamp 1586364061
transform 1 0 15996 0 -1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17468 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17284 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17560 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_182
timestamp 1586364061
transform 1 0 17376 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_186
timestamp 1586364061
transform 1 0 17744 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18756 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19124 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18940 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18572 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_197
timestamp 1586364061
transform 1 0 18756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_194
timestamp 1586364061
transform 1 0 18480 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 19584 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 20412 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20320 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 20412 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_210
timestamp 1586364061
transform 1 0 19952 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_214
timestamp 1586364061
transform 1 0 20320 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_217
timestamp 1586364061
transform 1 0 20596 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_221
timestamp 1586364061
transform 1 0 20964 0 1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21240 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21056 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_235
timestamp 1586364061
transform 1 0 22252 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_224
timestamp 1586364061
transform 1 0 21240 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 22896 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23080 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 23356 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 22988 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23172 0 1 20128
box -38 -48 774 592
use scs8hd_decap_6  FILLER_34_236
timestamp 1586364061
transform 1 0 22344 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_245
timestamp 1586364061
transform 1 0 23172 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_249
timestamp 1586364061
transform 1 0 23540 0 -1 21216
box -38 -48 590 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 24092 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 23908 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24368 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_262
timestamp 1586364061
transform 1 0 24736 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_259
timestamp 1586364061
transform 1 0 24460 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25104 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 25932 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25564 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 24920 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_269
timestamp 1586364061
transform 1 0 25380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_273
timestamp 1586364061
transform 1 0 25748 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_271
timestamp 1586364061
transform 1 0 25564 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26024 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26392 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26392 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 632 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1092 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 908 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_7
timestamp 1586364061
transform 1 0 1276 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_19
timestamp 1586364061
transform 1 0 2380 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3760 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4220 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_31
timestamp 1586364061
transform 1 0 3484 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_37
timestamp 1586364061
transform 1 0 4036 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_41
timestamp 1586364061
transform 1 0 4404 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_53
timestamp 1586364061
transform 1 0 5508 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6244 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_62
timestamp 1586364061
transform 1 0 6336 0 1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7348 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_70
timestamp 1586364061
transform 1 0 7072 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_82
timestamp 1586364061
transform 1 0 8176 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8912 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8728 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9924 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10292 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_99
timestamp 1586364061
transform 1 0 9740 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_103
timestamp 1586364061
transform 1 0 10108 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_107
timestamp 1586364061
transform 1 0 10476 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12040 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 11856 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 11580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 11764 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_123
timestamp 1586364061
transform 1 0 11948 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12500 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13328 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 12960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_127
timestamp 1586364061
transform 1 0 12316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_131
timestamp 1586364061
transform 1 0 12684 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_136
timestamp 1586364061
transform 1 0 13144 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13512 0 1 21216
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_35_151
timestamp 1586364061
transform 1 0 14524 0 1 21216
box -38 -48 314 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 15260 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14800 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15720 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_156
timestamp 1586364061
transform 1 0 14984 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 15536 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_166
timestamp 1586364061
transform 1 0 15904 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_178
timestamp 1586364061
transform 1 0 17008 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18388 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17468 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18204 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 17744 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_182
timestamp 1586364061
transform 1 0 17376 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_184
timestamp 1586364061
transform 1 0 17560 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_188
timestamp 1586364061
transform 1 0 17928 0 1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_35_202
timestamp 1586364061
transform 1 0 19216 0 1 21216
box -38 -48 590 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 20320 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20136 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 19768 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_210
timestamp 1586364061
transform 1 0 19952 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 21884 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 21700 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_223
timestamp 1586364061
transform 1 0 21148 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_227
timestamp 1586364061
transform 1 0 21516 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_235
timestamp 1586364061
transform 1 0 22252 0 1 21216
box -38 -48 222 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 23172 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23080 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22804 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22436 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_239
timestamp 1586364061
transform 1 0 22620 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 22988 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24736 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24368 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_254
timestamp 1586364061
transform 1 0 24000 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_260
timestamp 1586364061
transform 1 0 24552 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25196 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_265
timestamp 1586364061
transform 1 0 25012 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25380 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26392 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 908 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 632 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_6
timestamp 1586364061
transform 1 0 1184 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_18
timestamp 1586364061
transform 1 0 2288 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3484 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_30
timestamp 1586364061
transform 1 0 3392 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 3576 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 4680 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 5784 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 6888 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 7992 0 -1 22304
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9372 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9096 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9188 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10752 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_104
timestamp 1586364061
transform 1 0 10200 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 11580 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_6  FILLER_36_112
timestamp 1586364061
transform 1 0 10936 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_118
timestamp 1586364061
transform 1 0 11488 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 13144 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12592 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_128
timestamp 1586364061
transform 1 0 12408 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_132
timestamp 1586364061
transform 1 0 12776 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14156 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 13972 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14340 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14800 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 14708 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15812 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_163
timestamp 1586364061
transform 1 0 15628 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_167
timestamp 1586364061
transform 1 0 15996 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_36_179
timestamp 1586364061
transform 1 0 17100 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 17376 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18388 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_191
timestamp 1586364061
transform 1 0 18204 0 -1 22304
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 19308 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_195
timestamp 1586364061
transform 1 0 18572 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_8  FILLER_36_206
timestamp 1586364061
transform 1 0 19584 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20412 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20320 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_224
timestamp 1586364061
transform 1 0 21240 0 -1 22304
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22804 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_236
timestamp 1586364061
transform 1 0 22344 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_240
timestamp 1586364061
transform 1 0 22712 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24368 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23816 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_250
timestamp 1586364061
transform 1 0 23632 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_254
timestamp 1586364061
transform 1 0 24000 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_261
timestamp 1586364061
transform 1 0 24644 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 25932 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_273
timestamp 1586364061
transform 1 0 25748 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26024 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26392 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 632 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 908 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2012 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4220 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5324 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6244 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6060 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6336 0 1 22304
box -38 -48 1142 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 8268 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_74
timestamp 1586364061
transform 1 0 7440 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_82
timestamp 1586364061
transform 1 0 8176 0 1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9280 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9096 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8728 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_86
timestamp 1586364061
transform 1 0 8544 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_90
timestamp 1586364061
transform 1 0 8912 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 10292 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10660 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_103
timestamp 1586364061
transform 1 0 10108 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_107
timestamp 1586364061
transform 1 0 10476 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10844 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11948 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 11856 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11672 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11304 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11488 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12960 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13328 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 12776 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_136
timestamp 1586364061
transform 1 0 13144 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13972 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13788 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_140
timestamp 1586364061
transform 1 0 13512 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15536 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14984 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15352 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_154
timestamp 1586364061
transform 1 0 14800 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_158
timestamp 1586364061
transform 1 0 15168 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16548 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16916 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_171
timestamp 1586364061
transform 1 0 16364 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 16732 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_179
timestamp 1586364061
transform 1 0 17100 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17468 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18388 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19124 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18572 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18940 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19584 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_197
timestamp 1586364061
transform 1 0 18756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_204
timestamp 1586364061
transform 1 0 19400 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20596 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20412 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_208
timestamp 1586364061
transform 1 0 19768 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_214
timestamp 1586364061
transform 1 0 20320 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21608 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21976 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_226
timestamp 1586364061
transform 1 0 21424 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_230
timestamp 1586364061
transform 1 0 21792 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_234
timestamp 1586364061
transform 1 0 22160 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23080 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22528 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 22712 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24184 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24368 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_262
timestamp 1586364061
transform 1 0 24736 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 25840 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26392 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 632 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 908 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2012 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3116 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3484 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 3576 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 4680 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 5784 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 6888 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 7992 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 9188 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9096 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10752 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_102
timestamp 1586364061
transform 1 0 10016 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_6  FILLER_38_119
timestamp 1586364061
transform 1 0 11580 0 -1 23392
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12316 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 12132 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_136
timestamp 1586364061
transform 1 0 13144 0 -1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13880 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_146
timestamp 1586364061
transform 1 0 14064 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 14616 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14984 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 14708 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 14800 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_165
timestamp 1586364061
transform 1 0 15812 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16548 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15996 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_169
timestamp 1586364061
transform 1 0 16180 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18112 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17560 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_182
timestamp 1586364061
transform 1 0 17376 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_186
timestamp 1586364061
transform 1 0 17744 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_199
timestamp 1586364061
transform 1 0 18940 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20320 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20596 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20964 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20044 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_215
timestamp 1586364061
transform 1 0 20412 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_219
timestamp 1586364061
transform 1 0 20780 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21332 0 -1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_38_223
timestamp 1586364061
transform 1 0 21148 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_234
timestamp 1586364061
transform 1 0 22160 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22896 0 -1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24460 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_251
timestamp 1586364061
transform 1 0 23724 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_262
timestamp 1586364061
transform 1 0 24736 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 25932 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 25840 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26024 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26392 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1736 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 632 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 632 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_3
timestamp 1586364061
transform 1 0 908 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_11
timestamp 1586364061
transform 1 0 1644 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 908 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2748 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2196 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_15
timestamp 1586364061
transform 1 0 2012 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_19
timestamp 1586364061
transform 1 0 2380 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_26
timestamp 1586364061
transform 1 0 3024 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2012 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3116 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3484 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3208 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_30
timestamp 1586364061
transform 1 0 3392 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 3576 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4864 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5324 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_42
timestamp 1586364061
transform 1 0 4496 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_49
timestamp 1586364061
transform 1 0 5140 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_53
timestamp 1586364061
transform 1 0 5508 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 4680 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5876 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6888 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6244 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5876 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6060 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_62
timestamp 1586364061
transform 1 0 6336 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_56
timestamp 1586364061
transform 1 0 5784 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_60
timestamp 1586364061
transform 1 0 6152 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7992 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7992 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7164 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_75
timestamp 1586364061
transform 1 0 7532 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_79
timestamp 1586364061
transform 1 0 7900 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_82
timestamp 1586364061
transform 1 0 8176 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_72
timestamp 1586364061
transform 1 0 7256 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_83
timestamp 1586364061
transform 1 0 8268 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9188 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8544 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9096 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9188 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8360 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_89
timestamp 1586364061
transform 1 0 8820 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_95
timestamp 1586364061
transform 1 0 9372 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9004 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_96
timestamp 1586364061
transform 1 0 9464 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 10752 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9740 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10200 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_102
timestamp 1586364061
transform 1 0 10016 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_106
timestamp 1586364061
transform 1 0 10384 0 1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_40_108
timestamp 1586364061
transform 1 0 10568 0 -1 24480
box -38 -48 590 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 11120 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 11856 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11672 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 11304 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11120 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11488 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 11948 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_117
timestamp 1586364061
transform 1 0 11396 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 12132 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12316 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12132 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_136
timestamp 1586364061
transform 1 0 13144 0 1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_40_134
timestamp 1586364061
transform 1 0 12960 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13696 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13880 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13696 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 14340 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_147
timestamp 1586364061
transform 1 0 14156 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_151
timestamp 1586364061
transform 1 0 14524 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 13972 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 14892 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 14800 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 14708 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 14708 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_164
timestamp 1586364061
transform 1 0 15720 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_158
timestamp 1586364061
transform 1 0 15168 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 16732 0 -1 24480
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16456 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 16916 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16272 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 16732 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17100 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_170
timestamp 1586364061
transform 1 0 16272 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_174
timestamp 1586364061
transform 1 0 16640 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 18296 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17652 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17468 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17744 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_184
timestamp 1586364061
transform 1 0 17560 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_184
timestamp 1586364061
transform 1 0 17560 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_188
timestamp 1586364061
transform 1 0 17928 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 19492 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 19308 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 18664 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_194
timestamp 1586364061
transform 1 0 18480 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_198
timestamp 1586364061
transform 1 0 18848 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_202
timestamp 1586364061
transform 1 0 19216 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_196
timestamp 1586364061
transform 1 0 18664 0 -1 24480
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20412 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20596 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20320 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20412 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20044 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_209
timestamp 1586364061
transform 1 0 19860 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_213
timestamp 1586364061
transform 1 0 20228 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_208
timestamp 1586364061
transform 1 0 19768 0 -1 24480
box -38 -48 590 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 22068 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21608 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 22068 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_226
timestamp 1586364061
transform 1 0 21424 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_230
timestamp 1586364061
transform 1 0 21792 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_235
timestamp 1586364061
transform 1 0 22252 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_224
timestamp 1586364061
transform 1 0 21240 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_232
timestamp 1586364061
transform 1 0 21976 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 23172 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 23356 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23080 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 22896 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 22528 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_240
timestamp 1586364061
transform 1 0 22712 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_237
timestamp 1586364061
transform 1 0 22436 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_245
timestamp 1586364061
transform 1 0 23172 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24736 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24460 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24460 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_254
timestamp 1586364061
transform 1 0 24000 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_258
timestamp 1586364061
transform 1 0 24368 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_261
timestamp 1586364061
transform 1 0 24644 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_251
timestamp 1586364061
transform 1 0 23724 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_262
timestamp 1586364061
transform 1 0 24736 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 25932 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25196 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_265
timestamp 1586364061
transform 1 0 25012 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25380 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 25840 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26024 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26392 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26392 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 632 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 908 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2012 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3116 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4220 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5324 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6244 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6060 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6336 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7440 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 8544 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 9648 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_41_110
timestamp 1586364061
transform 1 0 10752 0 1 24480
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10844 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 11856 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11304 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11120 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_118
timestamp 1586364061
transform 1 0 11488 0 1 24480
box -38 -48 406 592
use scs8hd_decap_6  FILLER_41_123
timestamp 1586364061
transform 1 0 11948 0 1 24480
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12592 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13052 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_129
timestamp 1586364061
transform 1 0 12500 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_133
timestamp 1586364061
transform 1 0 12868 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_137
timestamp 1586364061
transform 1 0 13236 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 14248 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13420 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_141
timestamp 1586364061
transform 1 0 13604 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_147
timestamp 1586364061
transform 1 0 14156 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_152
timestamp 1586364061
transform 1 0 14616 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15352 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15812 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 14800 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_156
timestamp 1586364061
transform 1 0 14984 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_163
timestamp 1586364061
transform 1 0 15628 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_167
timestamp 1586364061
transform 1 0 15996 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_41_179
timestamp 1586364061
transform 1 0 17100 0 1 24480
box -38 -48 406 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 17652 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17468 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_184
timestamp 1586364061
transform 1 0 17560 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_188
timestamp 1586364061
transform 1 0 17928 0 1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 19584 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_200
timestamp 1586364061
transform 1 0 19032 0 1 24480
box -38 -48 590 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 19768 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20780 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_217
timestamp 1586364061
transform 1 0 20596 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_221
timestamp 1586364061
transform 1 0 20964 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21424 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21884 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_225
timestamp 1586364061
transform 1 0 21332 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_229
timestamp 1586364061
transform 1 0 21700 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_233
timestamp 1586364061
transform 1 0 22068 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23080 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_241
timestamp 1586364061
transform 1 0 22804 0 1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_41_245
timestamp 1586364061
transform 1 0 23172 0 1 24480
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23816 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24276 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_251
timestamp 1586364061
transform 1 0 23724 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_255
timestamp 1586364061
transform 1 0 24092 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_259
timestamp 1586364061
transform 1 0 24460 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24828 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25288 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_266
timestamp 1586364061
transform 1 0 25104 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_270
timestamp 1586364061
transform 1 0 25472 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_276
timestamp 1586364061
transform 1 0 26024 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26392 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 632 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 908 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3116 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3484 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 3576 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 4680 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6336 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 5784 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6428 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 7532 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9188 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 8636 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9280 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10384 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12040 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11488 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13052 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_125
timestamp 1586364061
transform 1 0 12132 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_133
timestamp 1586364061
transform 1 0 12868 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_138
timestamp 1586364061
transform 1 0 13328 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_150
timestamp 1586364061
transform 1 0 14432 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 14892 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_154
timestamp 1586364061
transform 1 0 14800 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 14984 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16088 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 17744 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17192 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 17836 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 18940 0 -1 25568
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20688 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 20596 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20044 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_221
timestamp 1586364061
transform 1 0 20964 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_233
timestamp 1586364061
transform 1 0 22068 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23448 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_245
timestamp 1586364061
transform 1 0 23172 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 23540 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 24644 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 25748 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26392 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4790 0 4846 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8286 0 8342 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 11782 0 11838 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15278 0 15334 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 18774 0 18830 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 22270 0 22326 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 27048 17960 27528 18080 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal3 s 27048 19048 27528 19168 6 chanx_right_in[1]
port 7 nsew default input
rlabel metal3 s 27048 20000 27528 20120 6 chanx_right_in[2]
port 8 nsew default input
rlabel metal3 s 27048 21088 27528 21208 6 chanx_right_in[3]
port 9 nsew default input
rlabel metal3 s 27048 22176 27528 22296 6 chanx_right_in[4]
port 10 nsew default input
rlabel metal3 s 27048 23128 27528 23248 6 chanx_right_in[5]
port 11 nsew default input
rlabel metal3 s 27048 24216 27528 24336 6 chanx_right_in[6]
port 12 nsew default input
rlabel metal3 s 27048 25304 27528 25424 6 chanx_right_in[7]
port 13 nsew default input
rlabel metal3 s 27048 26256 27528 26376 6 chanx_right_in[8]
port 14 nsew default input
rlabel metal3 s 27048 8712 27528 8832 6 chanx_right_out[0]
port 15 nsew default tristate
rlabel metal3 s 27048 9664 27528 9784 6 chanx_right_out[1]
port 16 nsew default tristate
rlabel metal3 s 27048 10752 27528 10872 6 chanx_right_out[2]
port 17 nsew default tristate
rlabel metal3 s 27048 11704 27528 11824 6 chanx_right_out[3]
port 18 nsew default tristate
rlabel metal3 s 27048 12792 27528 12912 6 chanx_right_out[4]
port 19 nsew default tristate
rlabel metal3 s 27048 13880 27528 14000 6 chanx_right_out[5]
port 20 nsew default tristate
rlabel metal3 s 27048 14832 27528 14952 6 chanx_right_out[6]
port 21 nsew default tristate
rlabel metal3 s 27048 15920 27528 16040 6 chanx_right_out[7]
port 22 nsew default tristate
rlabel metal3 s 27048 17008 27528 17128 6 chanx_right_out[8]
port 23 nsew default tristate
rlabel metal2 s 8286 27520 8342 28000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 9298 27520 9354 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 10310 27520 10366 28000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 11322 27520 11378 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 12426 27520 12482 28000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 13438 27520 13494 28000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 14450 27520 14506 28000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 15462 27520 15518 28000 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 16566 27520 16622 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 17578 27520 17634 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 18590 27520 18646 28000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 19602 27520 19658 28000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 20706 27520 20762 28000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 21718 27520 21774 28000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 22730 27520 22786 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 23742 27520 23798 28000 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 24846 27520 24902 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 25858 27520 25914 28000 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 25766 0 25822 480 6 data_in
port 42 nsew default input
rlabel metal2 s 1294 0 1350 480 6 enable
port 43 nsew default input
rlabel metal3 s 27048 5584 27528 5704 6 right_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 27048 6536 27528 6656 6 right_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal3 s 27048 7624 27528 7744 6 right_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 27048 416 27528 536 6 right_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 27048 1368 27528 1488 6 right_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 27048 2456 27528 2576 6 right_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal3 s 27048 3408 27528 3528 6 right_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 27048 4496 27528 4616 6 right_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 27048 27344 27528 27464 6 right_top_grid_pin_10_
port 52 nsew default input
rlabel metal2 s 5158 27520 5214 28000 6 top_left_grid_pin_11_
port 53 nsew default input
rlabel metal2 s 6170 27520 6226 28000 6 top_left_grid_pin_13_
port 54 nsew default input
rlabel metal2 s 7182 27520 7238 28000 6 top_left_grid_pin_15_
port 55 nsew default input
rlabel metal2 s 6 27520 62 28000 6 top_left_grid_pin_1_
port 56 nsew default input
rlabel metal2 s 1018 27520 1074 28000 6 top_left_grid_pin_3_
port 57 nsew default input
rlabel metal2 s 2030 27520 2086 28000 6 top_left_grid_pin_5_
port 58 nsew default input
rlabel metal2 s 3042 27520 3098 28000 6 top_left_grid_pin_7_
port 59 nsew default input
rlabel metal2 s 4146 27520 4202 28000 6 top_left_grid_pin_9_
port 60 nsew default input
rlabel metal2 s 26870 27520 26926 28000 6 top_right_grid_pin_11_
port 61 nsew default input
rlabel metal4 s 5139 2128 5459 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 9805 2128 10125 25616 6 vgnd
port 63 nsew default input
<< properties >>
string FIXED_BBOX 1 0 27528 28000
<< end >>
