magic
tech sky130A
magscale 1 2
timestamp 1606474215
<< locali >>
rect 13645 4539 13679 4641
rect 19349 3383 19383 3553
rect 14381 2907 14415 3145
rect 17785 2839 17819 3145
<< viali >>
rect 20729 20009 20763 20043
rect 20545 19873 20579 19907
rect 20177 19465 20211 19499
rect 16405 19261 16439 19295
rect 18521 19261 18555 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 16589 19125 16623 19159
rect 18705 19125 18739 19159
rect 20729 19125 20763 19159
rect 10057 18853 10091 18887
rect 15945 18853 15979 18887
rect 17969 18853 18003 18887
rect 19901 18853 19935 18887
rect 9781 18785 9815 18819
rect 12173 18785 12207 18819
rect 15669 18785 15703 18819
rect 17693 18785 17727 18819
rect 19625 18785 19659 18819
rect 12449 18717 12483 18751
rect 20177 18377 20211 18411
rect 20729 18377 20763 18411
rect 7757 18173 7791 18207
rect 19999 18173 20033 18207
rect 20545 18173 20579 18207
rect 8033 18105 8067 18139
rect 15485 17833 15519 17867
rect 20453 17833 20487 17867
rect 11345 17697 11379 17731
rect 15301 17697 15335 17731
rect 20275 17697 20309 17731
rect 11621 17629 11655 17663
rect 20177 17289 20211 17323
rect 20729 17289 20763 17323
rect 14473 17153 14507 17187
rect 14197 17085 14231 17119
rect 19993 17085 20027 17119
rect 20545 17085 20579 17119
rect 17325 16677 17359 16711
rect 17049 16609 17083 16643
rect 20729 16201 20763 16235
rect 19809 16065 19843 16099
rect 19533 15997 19567 16031
rect 20545 15997 20579 16031
rect 20453 15657 20487 15691
rect 11897 15521 11931 15555
rect 13829 15521 13863 15555
rect 20269 15521 20303 15555
rect 12173 15453 12207 15487
rect 14105 15453 14139 15487
rect 20177 15113 20211 15147
rect 20729 15113 20763 15147
rect 9781 14909 9815 14943
rect 19993 14909 20027 14943
rect 20545 14909 20579 14943
rect 10057 14841 10091 14875
rect 19901 14569 19935 14603
rect 20453 14569 20487 14603
rect 8401 14433 8435 14467
rect 19717 14433 19751 14467
rect 20269 14433 20303 14467
rect 8677 14365 8711 14399
rect 19533 14025 19567 14059
rect 17509 13957 17543 13991
rect 11161 13889 11195 13923
rect 10885 13821 10919 13855
rect 16129 13821 16163 13855
rect 16396 13821 16430 13855
rect 19349 13821 19383 13855
rect 19901 13821 19935 13855
rect 20729 13753 20763 13787
rect 19257 13481 19291 13515
rect 19901 13413 19935 13447
rect 19073 13345 19107 13379
rect 19625 13345 19659 13379
rect 15117 12937 15151 12971
rect 18061 12937 18095 12971
rect 19257 12937 19291 12971
rect 15761 12801 15795 12835
rect 18613 12801 18647 12835
rect 19809 12801 19843 12835
rect 19073 12733 19107 12767
rect 19625 12733 19659 12767
rect 20361 12733 20395 12767
rect 18521 12665 18555 12699
rect 20637 12665 20671 12699
rect 15485 12597 15519 12631
rect 15577 12597 15611 12631
rect 17509 12597 17543 12631
rect 18429 12597 18463 12631
rect 15485 12393 15519 12427
rect 17325 12393 17359 12427
rect 20453 12393 20487 12427
rect 17868 12325 17902 12359
rect 19717 12325 19751 12359
rect 13625 12257 13659 12291
rect 16212 12257 16246 12291
rect 17601 12257 17635 12291
rect 19441 12257 19475 12291
rect 20269 12257 20303 12291
rect 13369 12189 13403 12223
rect 15945 12189 15979 12223
rect 14749 12053 14783 12087
rect 18981 12053 19015 12087
rect 15209 11849 15243 11883
rect 16865 11849 16899 11883
rect 13461 11713 13495 11747
rect 18613 11713 18647 11747
rect 20729 11713 20763 11747
rect 20821 11713 20855 11747
rect 13185 11645 13219 11679
rect 13829 11645 13863 11679
rect 15485 11645 15519 11679
rect 15752 11645 15786 11679
rect 18061 11645 18095 11679
rect 18880 11645 18914 11679
rect 14096 11577 14130 11611
rect 12817 11509 12851 11543
rect 13277 11509 13311 11543
rect 18245 11509 18279 11543
rect 19993 11509 20027 11543
rect 20269 11509 20303 11543
rect 20637 11509 20671 11543
rect 14105 11305 14139 11339
rect 15301 11305 15335 11339
rect 18705 11305 18739 11339
rect 20545 11305 20579 11339
rect 15669 11237 15703 11271
rect 16129 11237 16163 11271
rect 19432 11237 19466 11271
rect 12716 11169 12750 11203
rect 15761 11169 15795 11203
rect 16497 11169 16531 11203
rect 17132 11169 17166 11203
rect 12449 11101 12483 11135
rect 15853 11101 15887 11135
rect 16865 11101 16899 11135
rect 19165 11101 19199 11135
rect 13829 11033 13863 11067
rect 16313 10965 16347 10999
rect 18245 10965 18279 10999
rect 15393 10761 15427 10795
rect 16589 10761 16623 10795
rect 19073 10693 19107 10727
rect 16037 10625 16071 10659
rect 17141 10625 17175 10659
rect 18613 10625 18647 10659
rect 19717 10625 19751 10659
rect 20545 10625 20579 10659
rect 20637 10625 20671 10659
rect 12449 10557 12483 10591
rect 19441 10557 19475 10591
rect 19533 10557 19567 10591
rect 12725 10489 12759 10523
rect 15761 10489 15795 10523
rect 17049 10489 17083 10523
rect 18521 10489 18555 10523
rect 15853 10421 15887 10455
rect 16957 10421 16991 10455
rect 18061 10421 18095 10455
rect 18429 10421 18463 10455
rect 20085 10421 20119 10455
rect 20453 10421 20487 10455
rect 13277 10217 13311 10251
rect 14749 10217 14783 10251
rect 17141 10217 17175 10251
rect 17868 10149 17902 10183
rect 19625 10149 19659 10183
rect 13645 10081 13679 10115
rect 13737 10081 13771 10115
rect 15557 10081 15591 10115
rect 17601 10081 17635 10115
rect 19717 10081 19751 10115
rect 20269 10081 20303 10115
rect 13829 10013 13863 10047
rect 15301 10013 15335 10047
rect 19809 10013 19843 10047
rect 18981 9945 19015 9979
rect 16681 9877 16715 9911
rect 19257 9877 19291 9911
rect 20453 9877 20487 9911
rect 11161 9605 11195 9639
rect 11713 9537 11747 9571
rect 13093 9537 13127 9571
rect 18429 9537 18463 9571
rect 13553 9469 13587 9503
rect 15393 9469 15427 9503
rect 15660 9469 15694 9503
rect 18696 9469 18730 9503
rect 20545 9469 20579 9503
rect 11529 9401 11563 9435
rect 13820 9401 13854 9435
rect 11621 9333 11655 9367
rect 14933 9333 14967 9367
rect 16773 9333 16807 9367
rect 19809 9333 19843 9367
rect 20729 9333 20763 9367
rect 9689 9129 9723 9163
rect 13829 9129 13863 9163
rect 15301 9129 15335 9163
rect 16405 9129 16439 9163
rect 10057 8993 10091 9027
rect 11060 8993 11094 9027
rect 12449 8993 12483 9027
rect 12716 8993 12750 9027
rect 13921 8993 13955 9027
rect 15669 8993 15703 9027
rect 16773 8993 16807 9027
rect 17417 8993 17451 9027
rect 19073 8993 19107 9027
rect 19340 8993 19374 9027
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 10793 8925 10827 8959
rect 14197 8925 14231 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 16865 8925 16899 8959
rect 16957 8925 16991 8959
rect 18613 8925 18647 8959
rect 12173 8789 12207 8823
rect 20453 8789 20487 8823
rect 11621 8585 11655 8619
rect 14565 8585 14599 8619
rect 18613 8585 18647 8619
rect 21097 8585 21131 8619
rect 11897 8449 11931 8483
rect 15117 8449 15151 8483
rect 19073 8449 19107 8483
rect 19257 8449 19291 8483
rect 8585 8381 8619 8415
rect 10241 8381 10275 8415
rect 14933 8381 14967 8415
rect 15393 8381 15427 8415
rect 15945 8381 15979 8415
rect 16212 8381 16246 8415
rect 18981 8381 19015 8415
rect 19717 8381 19751 8415
rect 19984 8381 20018 8415
rect 8852 8313 8886 8347
rect 10486 8313 10520 8347
rect 12725 8313 12759 8347
rect 15669 8313 15703 8347
rect 9965 8245 9999 8279
rect 14013 8245 14047 8279
rect 15025 8245 15059 8279
rect 17325 8245 17359 8279
rect 9321 8041 9355 8075
rect 9689 8041 9723 8075
rect 10609 8041 10643 8075
rect 12541 8041 12575 8075
rect 16221 8041 16255 8075
rect 19257 8041 19291 8075
rect 19809 8041 19843 8075
rect 10977 7973 11011 8007
rect 13820 7973 13854 8007
rect 17509 7973 17543 8007
rect 20177 7973 20211 8007
rect 7941 7905 7975 7939
rect 8208 7905 8242 7939
rect 10333 7905 10367 7939
rect 11069 7905 11103 7939
rect 12909 7905 12943 7939
rect 13001 7905 13035 7939
rect 15669 7905 15703 7939
rect 16589 7905 16623 7939
rect 17233 7905 17267 7939
rect 19165 7905 19199 7939
rect 11161 7837 11195 7871
rect 13185 7837 13219 7871
rect 13553 7837 13587 7871
rect 16681 7837 16715 7871
rect 16773 7837 16807 7871
rect 19349 7837 19383 7871
rect 20269 7837 20303 7871
rect 20453 7837 20487 7871
rect 10149 7701 10183 7735
rect 14933 7701 14967 7735
rect 15485 7701 15519 7735
rect 18797 7701 18831 7735
rect 14473 7497 14507 7531
rect 16865 7497 16899 7531
rect 11345 7429 11379 7463
rect 11989 7361 12023 7395
rect 15117 7361 15151 7395
rect 19809 7361 19843 7395
rect 20269 7361 20303 7395
rect 11253 7293 11287 7327
rect 12449 7293 12483 7327
rect 12705 7293 12739 7327
rect 15485 7293 15519 7327
rect 17325 7293 17359 7327
rect 14841 7225 14875 7259
rect 15752 7225 15786 7259
rect 19717 7225 19751 7259
rect 11069 7157 11103 7191
rect 11713 7157 11747 7191
rect 11805 7157 11839 7191
rect 13829 7157 13863 7191
rect 14933 7157 14967 7191
rect 17141 7157 17175 7191
rect 19257 7157 19291 7191
rect 19625 7157 19659 7191
rect 12357 6953 12391 6987
rect 13461 6953 13495 6987
rect 15301 6953 15335 6987
rect 15669 6953 15703 6987
rect 19349 6953 19383 6987
rect 16580 6885 16614 6919
rect 10057 6817 10091 6851
rect 10968 6817 11002 6851
rect 13829 6817 13863 6851
rect 16313 6817 16347 6851
rect 18236 6817 18270 6851
rect 19993 6817 20027 6851
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10701 6749 10735 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 17969 6749 18003 6783
rect 20085 6749 20119 6783
rect 20177 6749 20211 6783
rect 9689 6681 9723 6715
rect 12081 6681 12115 6715
rect 17693 6681 17727 6715
rect 19625 6681 19659 6715
rect 6837 6409 6871 6443
rect 9229 6409 9263 6443
rect 10885 6409 10919 6443
rect 11161 6409 11195 6443
rect 13185 6409 13219 6443
rect 7481 6273 7515 6307
rect 11713 6273 11747 6307
rect 13737 6273 13771 6307
rect 14657 6273 14691 6307
rect 17049 6273 17083 6307
rect 17417 6273 17451 6307
rect 18797 6273 18831 6307
rect 7849 6205 7883 6239
rect 9505 6205 9539 6239
rect 9772 6205 9806 6239
rect 14924 6205 14958 6239
rect 19064 6205 19098 6239
rect 20545 6205 20579 6239
rect 8116 6137 8150 6171
rect 13645 6137 13679 6171
rect 16865 6137 16899 6171
rect 7205 6069 7239 6103
rect 7297 6069 7331 6103
rect 11529 6069 11563 6103
rect 11621 6069 11655 6103
rect 13553 6069 13587 6103
rect 16037 6069 16071 6103
rect 16405 6069 16439 6103
rect 16773 6069 16807 6103
rect 18337 6069 18371 6103
rect 20177 6069 20211 6103
rect 20729 6069 20763 6103
rect 9045 5865 9079 5899
rect 9689 5865 9723 5899
rect 10425 5865 10459 5899
rect 15669 5865 15703 5899
rect 16773 5865 16807 5899
rect 17877 5865 17911 5899
rect 19257 5865 19291 5899
rect 6000 5797 6034 5831
rect 11704 5797 11738 5831
rect 19349 5797 19383 5831
rect 5733 5729 5767 5763
rect 7656 5729 7690 5763
rect 10333 5729 10367 5763
rect 10793 5729 10827 5763
rect 13093 5729 13127 5763
rect 13360 5729 13394 5763
rect 15761 5729 15795 5763
rect 16681 5729 16715 5763
rect 18245 5729 18279 5763
rect 20269 5729 20303 5763
rect 7389 5661 7423 5695
rect 10885 5661 10919 5695
rect 10977 5661 11011 5695
rect 11437 5661 11471 5695
rect 15945 5661 15979 5695
rect 16957 5661 16991 5695
rect 18337 5661 18371 5695
rect 18521 5661 18555 5695
rect 19441 5661 19475 5695
rect 8769 5593 8803 5627
rect 14473 5593 14507 5627
rect 15301 5593 15335 5627
rect 18889 5593 18923 5627
rect 7113 5525 7147 5559
rect 10149 5525 10183 5559
rect 12817 5525 12851 5559
rect 16313 5525 16347 5559
rect 20453 5525 20487 5559
rect 8217 5321 8251 5355
rect 8677 5321 8711 5355
rect 11529 5321 11563 5355
rect 14013 5321 14047 5355
rect 15945 5321 15979 5355
rect 18061 5321 18095 5355
rect 19625 5321 19659 5355
rect 20821 5253 20855 5287
rect 9229 5185 9263 5219
rect 11805 5185 11839 5219
rect 13553 5185 13587 5219
rect 14565 5185 14599 5219
rect 16405 5185 16439 5219
rect 16497 5185 16531 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 10149 5117 10183 5151
rect 14381 5117 14415 5151
rect 19073 5117 19107 5151
rect 19993 5117 20027 5151
rect 20637 5117 20671 5151
rect 10416 5049 10450 5083
rect 16313 5049 16347 5083
rect 18429 5049 18463 5083
rect 18521 5049 18555 5083
rect 9045 4981 9079 5015
rect 9137 4981 9171 5015
rect 14473 4981 14507 5015
rect 19257 4981 19291 5015
rect 20085 4981 20119 5015
rect 7113 4777 7147 4811
rect 8585 4777 8619 4811
rect 10609 4777 10643 4811
rect 14197 4777 14231 4811
rect 8953 4709 8987 4743
rect 9045 4709 9079 4743
rect 17316 4709 17350 4743
rect 19432 4709 19466 4743
rect 7481 4641 7515 4675
rect 10977 4641 11011 4675
rect 11069 4641 11103 4675
rect 13645 4641 13679 4675
rect 14289 4641 14323 4675
rect 17049 4641 17083 4675
rect 19165 4641 19199 4675
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 9137 4573 9171 4607
rect 11253 4573 11287 4607
rect 14473 4573 14507 4607
rect 13645 4505 13679 4539
rect 13829 4437 13863 4471
rect 18429 4437 18463 4471
rect 20545 4437 20579 4471
rect 9229 4233 9263 4267
rect 19441 4233 19475 4267
rect 19717 4233 19751 4267
rect 10885 4097 10919 4131
rect 13093 4097 13127 4131
rect 14657 4097 14691 4131
rect 20269 4097 20303 4131
rect 7849 4029 7883 4063
rect 13001 4029 13035 4063
rect 15209 4029 15243 4063
rect 15476 4029 15510 4063
rect 18061 4029 18095 4063
rect 20729 4029 20763 4063
rect 8116 3961 8150 3995
rect 9781 3961 9815 3995
rect 10609 3961 10643 3995
rect 18306 3961 18340 3995
rect 10241 3893 10275 3927
rect 10701 3893 10735 3927
rect 11805 3893 11839 3927
rect 12541 3893 12575 3927
rect 12909 3893 12943 3927
rect 14105 3893 14139 3927
rect 14473 3893 14507 3927
rect 14565 3893 14599 3927
rect 16589 3893 16623 3927
rect 17509 3893 17543 3927
rect 20085 3893 20119 3927
rect 20177 3893 20211 3927
rect 20913 3893 20947 3927
rect 8585 3689 8619 3723
rect 12725 3689 12759 3723
rect 17877 3689 17911 3723
rect 19441 3689 19475 3723
rect 9956 3621 9990 3655
rect 7205 3553 7239 3587
rect 7472 3553 7506 3587
rect 9689 3553 9723 3587
rect 11345 3553 11379 3587
rect 11612 3553 11646 3587
rect 13544 3553 13578 3587
rect 15301 3553 15335 3587
rect 15568 3553 15602 3587
rect 18705 3553 18739 3587
rect 19349 3553 19383 3587
rect 19809 3553 19843 3587
rect 8861 3485 8895 3519
rect 13277 3485 13311 3519
rect 17969 3485 18003 3519
rect 18153 3485 18187 3519
rect 18889 3485 18923 3519
rect 14657 3417 14691 3451
rect 19901 3485 19935 3519
rect 20085 3485 20119 3519
rect 11069 3349 11103 3383
rect 16681 3349 16715 3383
rect 17509 3349 17543 3383
rect 19349 3349 19383 3383
rect 8217 3145 8251 3179
rect 8493 3145 8527 3179
rect 10977 3145 11011 3179
rect 11345 3145 11379 3179
rect 14289 3145 14323 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 15117 3145 15151 3179
rect 17785 3145 17819 3179
rect 18061 3145 18095 3179
rect 19441 3145 19475 3179
rect 6837 3009 6871 3043
rect 9045 3009 9079 3043
rect 11989 3009 12023 3043
rect 7104 2941 7138 2975
rect 8861 2941 8895 2975
rect 8953 2941 8987 2975
rect 9597 2941 9631 2975
rect 9864 2941 9898 2975
rect 11713 2941 11747 2975
rect 12909 2941 12943 2975
rect 13176 2941 13210 2975
rect 15761 3009 15795 3043
rect 16681 3009 16715 3043
rect 14565 2941 14599 2975
rect 17417 2941 17451 2975
rect 11805 2873 11839 2907
rect 14381 2873 14415 2907
rect 16497 2873 16531 2907
rect 20729 3077 20763 3111
rect 18521 3009 18555 3043
rect 18705 3009 18739 3043
rect 19901 3009 19935 3043
rect 20085 3009 20119 3043
rect 18429 2941 18463 2975
rect 20545 2941 20579 2975
rect 12449 2805 12483 2839
rect 15485 2805 15519 2839
rect 15577 2805 15611 2839
rect 16129 2805 16163 2839
rect 16589 2805 16623 2839
rect 17601 2805 17635 2839
rect 17785 2805 17819 2839
rect 19809 2805 19843 2839
rect 7481 2601 7515 2635
rect 10149 2601 10183 2635
rect 13369 2601 13403 2635
rect 15853 2601 15887 2635
rect 16221 2601 16255 2635
rect 17877 2601 17911 2635
rect 20729 2601 20763 2635
rect 10517 2533 10551 2567
rect 10609 2533 10643 2567
rect 7849 2465 7883 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 16313 2465 16347 2499
rect 16957 2465 16991 2499
rect 17693 2465 17727 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 7941 2397 7975 2431
rect 8125 2397 8159 2431
rect 10793 2397 10827 2431
rect 13461 2397 13495 2431
rect 13645 2397 13679 2431
rect 16497 2397 16531 2431
rect 13001 2329 13035 2363
rect 18521 2329 18555 2363
rect 19625 2329 19659 2363
rect 11621 2261 11655 2295
rect 12173 2261 12207 2295
rect 17141 2261 17175 2295
rect 19073 2261 19107 2295
rect 20177 2261 20211 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 19944 19876 20545 19904
rect 19944 19864 19950 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 20162 19496 20168 19508
rect 20123 19468 20168 19496
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 15856 19332 16528 19360
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 15856 19292 15884 19332
rect 5776 19264 15884 19292
rect 5776 19252 5782 19264
rect 15930 19252 15936 19304
rect 15988 19292 15994 19304
rect 16393 19295 16451 19301
rect 16393 19292 16405 19295
rect 15988 19264 16405 19292
rect 15988 19252 15994 19264
rect 16393 19261 16405 19264
rect 16439 19261 16451 19295
rect 16500 19292 16528 19332
rect 17880 19332 18644 19360
rect 17880 19292 17908 19332
rect 16500 19264 17908 19292
rect 16393 19255 16451 19261
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18012 19264 18521 19292
rect 18012 19252 18018 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18616 19292 18644 19332
rect 19812 19332 20116 19360
rect 19812 19292 19840 19332
rect 19978 19292 19984 19304
rect 18616 19264 19840 19292
rect 19939 19264 19984 19292
rect 18509 19255 18567 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20088 19292 20116 19332
rect 20533 19295 20591 19301
rect 20533 19292 20545 19295
rect 20088 19264 20545 19292
rect 20533 19261 20545 19264
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 16577 19159 16635 19165
rect 16577 19125 16589 19159
rect 16623 19156 16635 19159
rect 17862 19156 17868 19168
rect 16623 19128 17868 19156
rect 16623 19125 16635 19128
rect 16577 19119 16635 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18690 19156 18696 19168
rect 18651 19128 18696 19156
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 20898 19156 20904 19168
rect 20763 19128 20904 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 20530 18952 20536 18964
rect 10060 18924 20536 18952
rect 10060 18893 10088 18924
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18853 10103 18887
rect 15930 18884 15936 18896
rect 15891 18856 15936 18884
rect 10045 18847 10103 18853
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 17954 18884 17960 18896
rect 17915 18856 17960 18884
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 19886 18884 19892 18896
rect 19847 18856 19892 18884
rect 19886 18844 19892 18856
rect 19944 18844 19950 18896
rect 9769 18819 9827 18825
rect 9769 18785 9781 18819
rect 9815 18816 9827 18819
rect 9950 18816 9956 18828
rect 9815 18788 9956 18816
rect 9815 18785 9827 18788
rect 9769 18779 9827 18785
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11756 18788 12173 18816
rect 11756 18776 11762 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 12161 18779 12219 18785
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 19610 18816 19616 18828
rect 17727 18788 18000 18816
rect 19571 18788 19616 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 17972 18760 18000 18788
rect 19610 18776 19616 18788
rect 19668 18776 19674 18828
rect 12437 18751 12495 18757
rect 12437 18717 12449 18751
rect 12483 18717 12495 18751
rect 12437 18711 12495 18717
rect 12452 18612 12480 18711
rect 17954 18708 17960 18760
rect 18012 18708 18018 18760
rect 19978 18612 19984 18624
rect 12452 18584 19984 18612
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 20162 18408 20168 18420
rect 20123 18380 20168 18408
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 7558 18164 7564 18216
rect 7616 18204 7622 18216
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 7616 18176 7757 18204
rect 7616 18164 7622 18176
rect 7745 18173 7757 18176
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 19987 18207 20045 18213
rect 19987 18173 19999 18207
rect 20033 18173 20045 18207
rect 20530 18204 20536 18216
rect 20491 18176 20536 18204
rect 19987 18167 20045 18173
rect 8021 18139 8079 18145
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 19996 18136 20024 18167
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 8067 18108 20024 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 15473 17867 15531 17873
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 17862 17864 17868 17876
rect 15519 17836 17868 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 20438 17864 20444 17876
rect 20399 17836 20444 17864
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 10870 17688 10876 17740
rect 10928 17728 10934 17740
rect 11333 17731 11391 17737
rect 11333 17728 11345 17731
rect 10928 17700 11345 17728
rect 10928 17688 10934 17700
rect 11333 17697 11345 17700
rect 11379 17697 11391 17731
rect 11333 17691 11391 17697
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14516 17700 15301 17728
rect 14516 17688 14522 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 20263 17731 20321 17737
rect 20263 17697 20275 17731
rect 20309 17697 20321 17731
rect 20263 17691 20321 17697
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17660 11667 17663
rect 20272 17660 20300 17691
rect 11655 17632 20300 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 14056 17088 14197 17116
rect 14056 17076 14062 17088
rect 14185 17085 14197 17088
rect 14231 17085 14243 17119
rect 19978 17116 19984 17128
rect 19939 17088 19984 17116
rect 14185 17079 14243 17085
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 20530 17116 20536 17128
rect 20491 17088 20536 17116
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 17313 16711 17371 16717
rect 17313 16677 17325 16711
rect 17359 16708 17371 16711
rect 20530 16708 20536 16720
rect 17359 16680 20536 16708
rect 17359 16677 17371 16680
rect 17313 16671 17371 16677
rect 20530 16668 20536 16680
rect 20588 16668 20594 16720
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 17037 16643 17095 16649
rect 17037 16640 17049 16643
rect 16448 16612 17049 16640
rect 16448 16600 16454 16612
rect 17037 16609 17049 16612
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 19978 16096 19984 16108
rect 19843 16068 19984 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 15436 16000 19533 16028
rect 15436 15988 15442 16000
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 19521 15991 19579 15997
rect 19610 15988 19616 16040
rect 19668 16028 19674 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 19668 16000 20545 16028
rect 19668 15988 19674 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 11882 15552 11888 15564
rect 11843 15524 11888 15552
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 13814 15552 13820 15564
rect 13775 15524 13820 15552
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 20257 15555 20315 15561
rect 20257 15521 20269 15555
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 19610 15484 19616 15496
rect 14139 15456 19616 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 12176 15416 12204 15447
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 20272 15416 20300 15515
rect 12176 15388 20300 15416
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 20162 15144 20168 15156
rect 20123 15116 20168 15144
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20714 15144 20720 15156
rect 20675 15116 20720 15144
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 9766 14940 9772 14952
rect 9727 14912 9772 14940
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 10045 14875 10103 14881
rect 10045 14841 10057 14875
rect 10091 14872 10103 14875
rect 20548 14872 20576 14903
rect 10091 14844 20576 14872
rect 10091 14841 10103 14844
rect 10045 14835 10103 14841
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 20070 14600 20076 14612
rect 19935 14572 20076 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20438 14600 20444 14612
rect 20399 14572 20444 14600
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 8478 14464 8484 14476
rect 8435 14436 8484 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 20257 14467 20315 14473
rect 20257 14433 20269 14467
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 19978 14396 19984 14408
rect 8711 14368 19984 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 11146 14288 11152 14340
rect 11204 14328 11210 14340
rect 20272 14328 20300 14427
rect 11204 14300 20300 14328
rect 11204 14288 11210 14300
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19300 14028 19533 14056
rect 19300 14016 19306 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17497 13991 17555 13997
rect 17497 13988 17509 13991
rect 17368 13960 17509 13988
rect 17368 13948 17374 13960
rect 17497 13957 17509 13960
rect 17543 13957 17555 13991
rect 17497 13951 17555 13957
rect 11146 13920 11152 13932
rect 11107 13892 11152 13920
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10284 13824 10885 13852
rect 10284 13812 10290 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 16114 13852 16120 13864
rect 16075 13824 16120 13852
rect 10873 13815 10931 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16384 13855 16442 13861
rect 16384 13821 16396 13855
rect 16430 13852 16442 13855
rect 16666 13852 16672 13864
rect 16430 13824 16672 13852
rect 16430 13821 16442 13824
rect 16384 13815 16442 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 19337 13855 19395 13861
rect 19337 13821 19349 13855
rect 19383 13821 19395 13855
rect 19886 13852 19892 13864
rect 19847 13824 19892 13852
rect 19337 13815 19395 13821
rect 19352 13784 19380 13815
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 19794 13784 19800 13796
rect 19352 13756 19800 13784
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 20717 13787 20775 13793
rect 20717 13784 20729 13787
rect 19904 13756 20729 13784
rect 18782 13676 18788 13728
rect 18840 13716 18846 13728
rect 19904 13716 19932 13756
rect 20717 13753 20729 13756
rect 20763 13753 20775 13787
rect 20717 13747 20775 13753
rect 18840 13688 19932 13716
rect 18840 13676 18846 13688
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 19242 13512 19248 13524
rect 19203 13484 19248 13512
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19702 13404 19708 13456
rect 19760 13444 19766 13456
rect 19889 13447 19947 13453
rect 19889 13444 19901 13447
rect 19760 13416 19901 13444
rect 19760 13404 19766 13416
rect 19889 13413 19901 13416
rect 19935 13413 19947 13447
rect 19889 13407 19947 13413
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13376 19119 13379
rect 19334 13376 19340 13388
rect 19107 13348 19340 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13345 19671 13379
rect 19613 13339 19671 13345
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 19628 13308 19656 13339
rect 12676 13280 19656 13308
rect 12676 13268 12682 13280
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 15105 12971 15163 12977
rect 15105 12937 15117 12971
rect 15151 12968 15163 12971
rect 15654 12968 15660 12980
rect 15151 12940 15660 12968
rect 15151 12937 15163 12940
rect 15105 12931 15163 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18049 12971 18107 12977
rect 18049 12968 18061 12971
rect 18012 12940 18061 12968
rect 18012 12928 18018 12940
rect 18049 12937 18061 12940
rect 18095 12937 18107 12971
rect 19242 12968 19248 12980
rect 19203 12940 19248 12968
rect 18049 12931 18107 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 13906 12860 13912 12912
rect 13964 12900 13970 12912
rect 13964 12872 19656 12900
rect 13964 12860 13970 12872
rect 15746 12832 15752 12844
rect 15707 12804 15752 12832
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 19628 12773 19656 12872
rect 19794 12832 19800 12844
rect 19755 12804 19800 12832
rect 19794 12792 19800 12804
rect 19852 12792 19858 12844
rect 19061 12767 19119 12773
rect 19061 12764 19073 12767
rect 17552 12736 19073 12764
rect 17552 12724 17558 12736
rect 19061 12733 19073 12736
rect 19107 12733 19119 12767
rect 19061 12727 19119 12733
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 19613 12727 19671 12733
rect 19812 12736 20361 12764
rect 19812 12708 19840 12736
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 16574 12656 16580 12708
rect 16632 12696 16638 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 16632 12668 18521 12696
rect 16632 12656 16638 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 19794 12656 19800 12708
rect 19852 12656 19858 12708
rect 20254 12656 20260 12708
rect 20312 12696 20318 12708
rect 20625 12699 20683 12705
rect 20625 12696 20637 12699
rect 20312 12668 20637 12696
rect 20312 12656 20318 12668
rect 20625 12665 20637 12668
rect 20671 12665 20683 12699
rect 20625 12659 20683 12665
rect 15470 12628 15476 12640
rect 15431 12600 15476 12628
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 17497 12631 17555 12637
rect 15620 12600 15665 12628
rect 15620 12588 15626 12600
rect 17497 12597 17509 12631
rect 17543 12628 17555 12631
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 17543 12600 18429 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 18417 12597 18429 12600
rect 18463 12597 18475 12631
rect 18417 12591 18475 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 11054 12424 11060 12436
rect 10928 12396 11060 12424
rect 10928 12384 10934 12396
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 15470 12424 15476 12436
rect 15431 12396 15476 12424
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 17313 12427 17371 12433
rect 17313 12393 17325 12427
rect 17359 12393 17371 12427
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 17313 12387 17371 12393
rect 16114 12356 16120 12368
rect 15948 12328 16120 12356
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 13613 12291 13671 12297
rect 13613 12288 13625 12291
rect 13504 12260 13625 12288
rect 13504 12248 13510 12260
rect 13613 12257 13625 12260
rect 13659 12257 13671 12291
rect 13613 12251 13671 12257
rect 13354 12220 13360 12232
rect 13315 12192 13360 12220
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15948 12229 15976 12328
rect 16114 12316 16120 12328
rect 16172 12356 16178 12368
rect 17328 12356 17356 12387
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 17856 12359 17914 12365
rect 17856 12356 17868 12359
rect 16172 12328 16896 12356
rect 17328 12328 17868 12356
rect 16172 12316 16178 12328
rect 16200 12291 16258 12297
rect 16200 12257 16212 12291
rect 16246 12288 16258 12291
rect 16758 12288 16764 12300
rect 16246 12260 16764 12288
rect 16246 12257 16258 12260
rect 16200 12251 16258 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16868 12288 16896 12328
rect 17856 12325 17868 12328
rect 17902 12356 17914 12359
rect 18598 12356 18604 12368
rect 17902 12328 18604 12356
rect 17902 12325 17914 12328
rect 17856 12319 17914 12325
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19705 12359 19763 12365
rect 19705 12356 19717 12359
rect 19392 12328 19717 12356
rect 19392 12316 19398 12328
rect 19705 12325 19717 12328
rect 19751 12325 19763 12359
rect 19705 12319 19763 12325
rect 17586 12288 17592 12300
rect 16868 12260 17592 12288
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 18616 12260 19441 12288
rect 18616 12232 18644 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 20254 12288 20260 12300
rect 20215 12260 20260 12288
rect 19429 12251 19487 12257
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15344 12192 15945 12220
rect 15344 12180 15350 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 18598 12180 18604 12232
rect 18656 12180 18662 12232
rect 14737 12087 14795 12093
rect 14737 12053 14749 12087
rect 14783 12084 14795 12087
rect 15838 12084 15844 12096
rect 14783 12056 15844 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18932 12056 18981 12084
rect 18932 12044 18938 12056
rect 18969 12053 18981 12056
rect 19015 12053 19027 12087
rect 18969 12047 19027 12053
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 15197 11883 15255 11889
rect 15197 11849 15209 11883
rect 15243 11880 15255 11883
rect 15746 11880 15752 11892
rect 15243 11852 15752 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 16853 11883 16911 11889
rect 16853 11880 16865 11883
rect 16816 11852 16865 11880
rect 16816 11840 16822 11852
rect 16853 11849 16865 11852
rect 16899 11849 16911 11883
rect 16853 11843 16911 11849
rect 13446 11744 13452 11756
rect 13407 11716 13452 11744
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 17586 11704 17592 11756
rect 17644 11744 17650 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17644 11716 18613 11744
rect 17644 11704 17650 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 13170 11676 13176 11688
rect 13131 11648 13176 11676
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 13412 11648 13829 11676
rect 13412 11636 13418 11648
rect 13817 11645 13829 11648
rect 13863 11676 13875 11679
rect 15286 11676 15292 11688
rect 13863 11648 15292 11676
rect 13863 11645 13875 11648
rect 13817 11639 13875 11645
rect 15286 11636 15292 11648
rect 15344 11676 15350 11688
rect 15746 11685 15752 11688
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 15344 11648 15485 11676
rect 15344 11636 15350 11648
rect 15473 11645 15485 11648
rect 15519 11645 15531 11679
rect 15740 11676 15752 11685
rect 15707 11648 15752 11676
rect 15473 11639 15531 11645
rect 15740 11639 15752 11648
rect 15746 11636 15752 11639
rect 15804 11636 15810 11688
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11676 18107 11679
rect 18506 11676 18512 11688
rect 18095 11648 18512 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18616 11676 18644 11707
rect 20622 11704 20628 11756
rect 20680 11744 20686 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20680 11716 20729 11744
rect 20680 11704 20686 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 18690 11676 18696 11688
rect 18616 11648 18696 11676
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 18874 11685 18880 11688
rect 18868 11676 18880 11685
rect 18787 11648 18880 11676
rect 18868 11639 18880 11648
rect 18932 11676 18938 11688
rect 20824 11676 20852 11707
rect 18932 11648 20852 11676
rect 18874 11636 18880 11639
rect 18932 11636 18938 11648
rect 14084 11611 14142 11617
rect 12820 11580 14044 11608
rect 12820 11549 12848 11580
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11509 12863 11543
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 12805 11503 12863 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 14016 11540 14044 11580
rect 14084 11577 14096 11611
rect 14130 11608 14142 11611
rect 15838 11608 15844 11620
rect 14130 11580 15844 11608
rect 14130 11577 14142 11580
rect 14084 11571 14142 11577
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 19518 11608 19524 11620
rect 16132 11580 19524 11608
rect 16132 11540 16160 11580
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 21910 11608 21916 11620
rect 19812 11580 21916 11608
rect 14016 11512 16160 11540
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 19812 11540 19840 11580
rect 21910 11568 21916 11580
rect 21968 11568 21974 11620
rect 19978 11540 19984 11552
rect 18279 11512 19840 11540
rect 19939 11512 19984 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20254 11540 20260 11552
rect 20215 11512 20260 11540
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20625 11543 20683 11549
rect 20625 11540 20637 11543
rect 20496 11512 20637 11540
rect 20496 11500 20502 11512
rect 20625 11509 20637 11512
rect 20671 11509 20683 11543
rect 20625 11503 20683 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13228 11308 14105 11336
rect 13228 11296 13234 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15562 11336 15568 11348
rect 15335 11308 15568 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 19334 11336 19340 11348
rect 18739 11308 19340 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20533 11339 20591 11345
rect 20533 11305 20545 11339
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 9640 11240 15669 11268
rect 9640 11228 9646 11240
rect 15657 11237 15669 11240
rect 15703 11268 15715 11271
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 15703 11240 16129 11268
rect 15703 11237 15715 11240
rect 15657 11231 15715 11237
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 18874 11268 18880 11280
rect 16117 11231 16175 11237
rect 16224 11240 18880 11268
rect 12704 11203 12762 11209
rect 12704 11169 12716 11203
rect 12750 11200 12762 11203
rect 13170 11200 13176 11212
rect 12750 11172 13176 11200
rect 12750 11169 12762 11172
rect 12704 11163 12762 11169
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 15930 11200 15936 11212
rect 15795 11172 15936 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 12437 11135 12495 11141
rect 12437 11132 12449 11135
rect 10836 11104 12449 11132
rect 10836 11092 10842 11104
rect 12437 11101 12449 11104
rect 12483 11101 12495 11135
rect 15838 11132 15844 11144
rect 15799 11104 15844 11132
rect 12437 11095 12495 11101
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4120 11036 12480 11064
rect 4120 11024 4126 11036
rect 12452 10996 12480 11036
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13817 11067 13875 11073
rect 13817 11064 13829 11067
rect 13504 11036 13829 11064
rect 13504 11024 13510 11036
rect 13817 11033 13829 11036
rect 13863 11033 13875 11067
rect 16224 11064 16252 11240
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 19420 11271 19478 11277
rect 19420 11237 19432 11271
rect 19466 11268 19478 11271
rect 19978 11268 19984 11280
rect 19466 11240 19984 11268
rect 19466 11237 19478 11240
rect 19420 11231 19478 11237
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 16298 11160 16304 11212
rect 16356 11200 16362 11212
rect 16485 11203 16543 11209
rect 16485 11200 16497 11203
rect 16356 11172 16497 11200
rect 16356 11160 16362 11172
rect 16485 11169 16497 11172
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 17120 11203 17178 11209
rect 17120 11169 17132 11203
rect 17166 11200 17178 11203
rect 20548 11200 20576 11299
rect 20622 11200 20628 11212
rect 17166 11172 20628 11200
rect 17166 11169 17178 11172
rect 17120 11163 17178 11169
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 13817 11027 13875 11033
rect 13924 11036 16252 11064
rect 16316 11104 16865 11132
rect 13924 10996 13952 11036
rect 12452 10968 13952 10996
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 16316 11005 16344 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 18748 11104 19165 11132
rect 18748 11092 18754 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 15344 10968 16313 10996
rect 15344 10956 15350 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 16301 10959 16359 10965
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18233 10999 18291 11005
rect 18233 10996 18245 10999
rect 18012 10968 18245 10996
rect 18012 10956 18018 10968
rect 18233 10965 18245 10968
rect 18279 10965 18291 10999
rect 18233 10959 18291 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 16574 10792 16580 10804
rect 16535 10764 16580 10792
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 19061 10727 19119 10733
rect 19061 10693 19073 10727
rect 19107 10693 19119 10727
rect 19061 10687 19119 10693
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16482 10656 16488 10668
rect 16071 10628 16488 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 17129 10659 17187 10665
rect 17129 10656 17141 10659
rect 16816 10628 17141 10656
rect 16816 10616 16822 10628
rect 17129 10625 17141 10628
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18012 10628 18613 10656
rect 18012 10616 18018 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 19076 10588 19104 10687
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 19978 10656 19984 10668
rect 19751 10628 19984 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20530 10656 20536 10668
rect 20491 10628 20536 10656
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 20680 10628 20725 10656
rect 20680 10616 20686 10628
rect 12483 10560 19104 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19392 10560 19441 10588
rect 19392 10548 19398 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20254 10588 20260 10600
rect 19567 10560 20260 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12713 10523 12771 10529
rect 12713 10520 12725 10523
rect 12032 10492 12725 10520
rect 12032 10480 12038 10492
rect 12713 10489 12725 10492
rect 12759 10489 12771 10523
rect 15746 10520 15752 10532
rect 15707 10492 15752 10520
rect 12713 10483 12771 10489
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 16666 10480 16672 10532
rect 16724 10520 16730 10532
rect 17037 10523 17095 10529
rect 17037 10520 17049 10523
rect 16724 10492 17049 10520
rect 16724 10480 16730 10492
rect 17037 10489 17049 10492
rect 17083 10489 17095 10523
rect 17037 10483 17095 10489
rect 18509 10523 18567 10529
rect 18509 10489 18521 10523
rect 18555 10520 18567 10523
rect 18555 10492 20116 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 658 10412 664 10464
rect 716 10452 722 10464
rect 9582 10452 9588 10464
rect 716 10424 9588 10452
rect 716 10412 722 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 15838 10452 15844 10464
rect 15799 10424 15844 10452
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16942 10452 16948 10464
rect 16903 10424 16948 10452
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18414 10452 18420 10464
rect 18375 10424 18420 10452
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 20088 10461 20116 10492
rect 20073 10455 20131 10461
rect 20073 10421 20085 10455
rect 20119 10421 20131 10455
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 20073 10415 20131 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13814 10248 13820 10260
rect 13311 10220 13820 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 15746 10248 15752 10260
rect 14783 10220 15752 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 18414 10248 18420 10260
rect 17175 10220 18420 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 17856 10183 17914 10189
rect 15344 10152 17632 10180
rect 15344 10140 15350 10152
rect 17604 10124 17632 10152
rect 17856 10149 17868 10183
rect 17902 10180 17914 10183
rect 17954 10180 17960 10192
rect 17902 10152 17960 10180
rect 17902 10149 17914 10152
rect 17856 10143 17914 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 19613 10183 19671 10189
rect 19613 10149 19625 10183
rect 19659 10180 19671 10183
rect 19978 10180 19984 10192
rect 19659 10152 19984 10180
rect 19659 10149 19671 10152
rect 19613 10143 19671 10149
rect 19978 10140 19984 10152
rect 20036 10180 20042 10192
rect 20438 10180 20444 10192
rect 20036 10152 20444 10180
rect 20036 10140 20042 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13136 10084 13645 10112
rect 13136 10072 13142 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14550 10112 14556 10124
rect 13771 10084 14556 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 15545 10115 15603 10121
rect 15545 10112 15557 10115
rect 15252 10084 15557 10112
rect 15252 10072 15258 10084
rect 15545 10081 15557 10084
rect 15591 10081 15603 10115
rect 17586 10112 17592 10124
rect 17499 10084 17592 10112
rect 15545 10075 15603 10081
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20257 10115 20315 10121
rect 19760 10084 19805 10112
rect 19760 10072 19766 10084
rect 20257 10081 20269 10115
rect 20303 10112 20315 10115
rect 20346 10112 20352 10124
rect 20303 10084 20352 10112
rect 20303 10081 20315 10084
rect 20257 10075 20315 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 13814 10044 13820 10056
rect 13775 10016 13820 10044
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 18984 10016 19809 10044
rect 18984 9988 19012 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 18966 9976 18972 9988
rect 18879 9948 18972 9976
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 16540 9880 16681 9908
rect 16540 9868 16546 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 19058 9868 19064 9920
rect 19116 9908 19122 9920
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 19116 9880 19257 9908
rect 19116 9868 19122 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 20441 9911 20499 9917
rect 20441 9908 20453 9911
rect 19576 9880 20453 9908
rect 19576 9868 19582 9880
rect 20441 9877 20453 9880
rect 20487 9877 20499 9911
rect 20441 9871 20499 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 11882 9636 11888 9648
rect 11195 9608 11888 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11882 9596 11888 9608
rect 11940 9596 11946 9648
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11664 9540 11713 9568
rect 11664 9528 11670 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 11701 9531 11759 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18414 9568 18420 9580
rect 17644 9540 18420 9568
rect 17644 9528 17650 9540
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 12492 9472 13553 9500
rect 12492 9460 12498 9472
rect 13541 9469 13553 9472
rect 13587 9500 13599 9503
rect 15286 9500 15292 9512
rect 13587 9472 15292 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 15286 9460 15292 9472
rect 15344 9500 15350 9512
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15344 9472 15393 9500
rect 15344 9460 15350 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 15648 9503 15706 9509
rect 15648 9469 15660 9503
rect 15694 9500 15706 9503
rect 16482 9500 16488 9512
rect 15694 9472 16488 9500
rect 15694 9469 15706 9472
rect 15648 9463 15706 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 18684 9503 18742 9509
rect 18684 9469 18696 9503
rect 18730 9500 18742 9503
rect 18966 9500 18972 9512
rect 18730 9472 18972 9500
rect 18730 9469 18742 9472
rect 18684 9463 18742 9469
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 20533 9503 20591 9509
rect 20533 9500 20545 9503
rect 19300 9472 20545 9500
rect 19300 9460 19306 9472
rect 20533 9469 20545 9472
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 11517 9435 11575 9441
rect 11517 9401 11529 9435
rect 11563 9432 11575 9435
rect 11882 9432 11888 9444
rect 11563 9404 11888 9432
rect 11563 9401 11575 9404
rect 11517 9395 11575 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 13814 9441 13820 9444
rect 13808 9432 13820 9441
rect 13775 9404 13820 9432
rect 13808 9395 13820 9404
rect 13814 9392 13820 9395
rect 13872 9392 13878 9444
rect 13924 9404 20760 9432
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11112 9336 11621 9364
rect 11112 9324 11118 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 13924 9364 13952 9404
rect 12216 9336 13952 9364
rect 14921 9367 14979 9373
rect 12216 9324 12222 9336
rect 14921 9333 14933 9367
rect 14967 9364 14979 9367
rect 15194 9364 15200 9376
rect 14967 9336 15200 9364
rect 14967 9333 14979 9336
rect 14921 9327 14979 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 16758 9364 16764 9376
rect 16719 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 20732 9373 20760 9404
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 19484 9336 19809 9364
rect 19484 9324 19490 9336
rect 19797 9333 19809 9336
rect 19843 9333 19855 9367
rect 19797 9327 19855 9333
rect 20717 9367 20775 9373
rect 20717 9333 20729 9367
rect 20763 9333 20775 9367
rect 20717 9327 20775 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9766 9160 9772 9172
rect 9723 9132 9772 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 13814 9160 13820 9172
rect 13775 9132 13820 9160
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15838 9160 15844 9172
rect 15335 9132 15844 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 16390 9160 16396 9172
rect 16351 9132 16396 9160
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 15252 9064 15884 9092
rect 15252 9052 15258 9064
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9824 8996 10057 9024
rect 9824 8984 9830 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 11048 9027 11106 9033
rect 11048 8993 11060 9027
rect 11094 9024 11106 9027
rect 11606 9024 11612 9036
rect 11094 8996 11612 9024
rect 11094 8993 11106 8996
rect 11048 8987 11106 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12704 9027 12762 9033
rect 12492 8996 12537 9024
rect 12492 8984 12498 8996
rect 12704 8993 12716 9027
rect 12750 9024 12762 9027
rect 13909 9027 13967 9033
rect 12750 8996 13492 9024
rect 12750 8993 12762 8996
rect 12704 8987 12762 8993
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9916 8928 10149 8956
rect 9916 8916 9922 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10244 8888 10272 8919
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10744 8928 10793 8956
rect 10744 8916 10750 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 9364 8860 10272 8888
rect 9364 8848 9370 8860
rect 12161 8823 12219 8829
rect 12161 8789 12173 8823
rect 12207 8820 12219 8823
rect 13464 8820 13492 8996
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 13924 8888 13952 8987
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 14056 8996 15669 9024
rect 14056 8984 14062 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14366 8956 14372 8968
rect 14231 8928 14372 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 15746 8956 15752 8968
rect 15707 8928 15752 8956
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 15856 8965 15884 9064
rect 19168 9064 19371 9092
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 16807 8996 17417 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 18414 8984 18420 9036
rect 18472 9024 18478 9036
rect 19061 9027 19119 9033
rect 19061 9024 19073 9027
rect 18472 8996 19073 9024
rect 18472 8984 18478 8996
rect 19061 8993 19073 8996
rect 19107 8993 19119 9027
rect 19061 8987 19119 8993
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 16850 8956 16856 8968
rect 16811 8928 16856 8956
rect 15841 8919 15899 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 16942 8916 16948 8968
rect 17000 8956 17006 8968
rect 18601 8959 18659 8965
rect 17000 8928 17045 8956
rect 17000 8916 17006 8928
rect 18601 8925 18613 8959
rect 18647 8956 18659 8959
rect 18966 8956 18972 8968
rect 18647 8928 18972 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19168 8956 19196 9064
rect 19343 9036 19371 9064
rect 19325 8984 19331 9036
rect 19383 9024 19389 9036
rect 19383 8996 19428 9024
rect 19383 8984 19389 8996
rect 19076 8928 19196 8956
rect 17954 8888 17960 8900
rect 13924 8860 17960 8888
rect 17954 8848 17960 8860
rect 18012 8848 18018 8900
rect 15102 8820 15108 8832
rect 12207 8792 15108 8820
rect 12207 8789 12219 8792
rect 12161 8783 12219 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 18782 8820 18788 8832
rect 15252 8792 18788 8820
rect 15252 8780 15258 8792
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19076 8820 19104 8928
rect 19242 8820 19248 8832
rect 19076 8792 19248 8820
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 20438 8820 20444 8832
rect 20399 8792 20444 8820
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 11606 8616 11612 8628
rect 5132 8588 11192 8616
rect 11567 8588 11612 8616
rect 5132 8576 5138 8588
rect 11164 8548 11192 8588
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 14550 8616 14556 8628
rect 14511 8588 14556 8616
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 18601 8619 18659 8625
rect 18601 8616 18613 8619
rect 15396 8588 18613 8616
rect 13998 8548 14004 8560
rect 11164 8520 14004 8548
rect 13998 8508 14004 8520
rect 14056 8508 14062 8560
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 15102 8480 15108 8492
rect 15063 8452 15108 8480
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 10134 8412 10140 8424
rect 8619 8384 10140 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8588 8344 8616 8375
rect 10134 8372 10140 8384
rect 10192 8412 10198 8424
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 10192 8384 10241 8412
rect 10192 8372 10198 8384
rect 10229 8381 10241 8384
rect 10275 8381 10287 8415
rect 10229 8375 10287 8381
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8412 14979 8415
rect 15010 8412 15016 8424
rect 14967 8384 15016 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15396 8421 15424 8588
rect 18601 8585 18613 8588
rect 18647 8585 18659 8619
rect 18601 8579 18659 8585
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 21085 8619 21143 8625
rect 21085 8616 21097 8619
rect 18932 8588 21097 8616
rect 18932 8576 18938 8588
rect 21085 8585 21097 8588
rect 21131 8585 21143 8619
rect 21085 8579 21143 8585
rect 19058 8480 19064 8492
rect 19019 8452 19064 8480
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19242 8480 19248 8492
rect 19203 8452 19248 8480
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16022 8412 16028 8424
rect 15979 8384 16028 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 16200 8415 16258 8421
rect 16200 8381 16212 8415
rect 16246 8412 16258 8415
rect 16758 8412 16764 8424
rect 16246 8384 16764 8412
rect 16246 8381 16258 8384
rect 16200 8375 16258 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 18966 8412 18972 8424
rect 18927 8384 18972 8412
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 19972 8415 20030 8421
rect 19972 8381 19984 8415
rect 20018 8412 20030 8415
rect 20438 8412 20444 8424
rect 20018 8384 20444 8412
rect 20018 8381 20030 8384
rect 19972 8375 20030 8381
rect 8312 8316 8616 8344
rect 8840 8347 8898 8353
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 8312 8276 8340 8316
rect 8840 8313 8852 8347
rect 8886 8344 8898 8347
rect 9306 8344 9312 8356
rect 8886 8316 9312 8344
rect 8886 8313 8898 8316
rect 8840 8307 8898 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 10474 8347 10532 8353
rect 10474 8344 10486 8347
rect 9968 8316 10486 8344
rect 9968 8285 9996 8316
rect 10474 8313 10486 8316
rect 10520 8344 10532 8347
rect 10870 8344 10876 8356
rect 10520 8316 10876 8344
rect 10520 8313 10532 8316
rect 10474 8307 10532 8313
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 12713 8347 12771 8353
rect 12713 8313 12725 8347
rect 12759 8344 12771 8347
rect 15194 8344 15200 8356
rect 12759 8316 15200 8344
rect 12759 8313 12771 8316
rect 12713 8307 12771 8313
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 15654 8344 15660 8356
rect 15615 8316 15660 8344
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 16942 8344 16948 8356
rect 16172 8316 16948 8344
rect 16172 8304 16178 8316
rect 16942 8304 16948 8316
rect 17000 8344 17006 8356
rect 19720 8344 19748 8375
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 17000 8316 17356 8344
rect 17000 8304 17006 8316
rect 8260 8248 8340 8276
rect 9953 8279 10011 8285
rect 8260 8236 8266 8248
rect 9953 8245 9965 8279
rect 9999 8245 10011 8279
rect 9953 8239 10011 8245
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 13998 8276 14004 8288
rect 11020 8248 14004 8276
rect 11020 8236 11026 8248
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 14090 8236 14096 8288
rect 14148 8276 14154 8288
rect 15013 8279 15071 8285
rect 15013 8276 15025 8279
rect 14148 8248 15025 8276
rect 14148 8236 14154 8248
rect 15013 8245 15025 8248
rect 15059 8276 15071 8279
rect 17218 8276 17224 8288
rect 15059 8248 17224 8276
rect 15059 8245 15071 8248
rect 15013 8239 15071 8245
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 17328 8285 17356 8316
rect 19168 8316 19748 8344
rect 19168 8288 19196 8316
rect 17313 8279 17371 8285
rect 17313 8245 17325 8279
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 19150 8236 19156 8288
rect 19208 8236 19214 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 8202 8072 8208 8084
rect 7944 8044 8208 8072
rect 7944 7945 7972 8044
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 9306 8072 9312 8084
rect 9267 8044 9312 8072
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 9766 8072 9772 8084
rect 9723 8044 9772 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 11054 8072 11060 8084
rect 10643 8044 11060 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 13262 8072 13268 8084
rect 12575 8044 13268 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 16114 8072 16120 8084
rect 13924 8044 16120 8072
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 10965 8007 11023 8013
rect 10965 8004 10977 8007
rect 8444 7976 10977 8004
rect 8444 7964 8450 7976
rect 10965 7973 10977 7976
rect 11011 7973 11023 8007
rect 10965 7967 11023 7973
rect 13808 8007 13866 8013
rect 13808 7973 13820 8007
rect 13854 8004 13866 8007
rect 13924 8004 13952 8044
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16850 8072 16856 8084
rect 16255 8044 16856 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 19245 8075 19303 8081
rect 19245 8041 19257 8075
rect 19291 8072 19303 8075
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19291 8044 19809 8072
rect 19291 8041 19303 8044
rect 19245 8035 19303 8041
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 19797 8035 19855 8041
rect 13854 7976 13952 8004
rect 13854 7973 13866 7976
rect 13808 7967 13866 7973
rect 13998 7964 14004 8016
rect 14056 8004 14062 8016
rect 14056 7976 15700 8004
rect 14056 7964 14062 7976
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8196 7939 8254 7945
rect 8196 7905 8208 7939
rect 8242 7936 8254 7939
rect 9030 7936 9036 7948
rect 8242 7908 9036 7936
rect 8242 7905 8254 7908
rect 8196 7899 8254 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 10318 7936 10324 7948
rect 10279 7908 10324 7936
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7936 11115 7939
rect 11606 7936 11612 7948
rect 11103 7908 11612 7936
rect 11103 7905 11115 7908
rect 11057 7899 11115 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 12894 7936 12900 7948
rect 12855 7908 12900 7936
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 14090 7936 14096 7948
rect 13035 7908 14096 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 15672 7945 15700 7976
rect 15838 7964 15844 8016
rect 15896 8004 15902 8016
rect 17126 8004 17132 8016
rect 15896 7976 17132 8004
rect 15896 7964 15902 7976
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 17494 8004 17500 8016
rect 17455 7976 17500 8004
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 19978 7964 19984 8016
rect 20036 8004 20042 8016
rect 20165 8007 20223 8013
rect 20165 8004 20177 8007
rect 20036 7976 20177 8004
rect 20036 7964 20042 7976
rect 20165 7973 20177 7976
rect 20211 7973 20223 8007
rect 20165 7967 20223 7973
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 15804 7908 16589 7936
rect 15804 7896 15810 7908
rect 16577 7905 16589 7908
rect 16623 7905 16635 7939
rect 16577 7899 16635 7905
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7936 19211 7939
rect 20070 7936 20076 7948
rect 19199 7908 20076 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 13170 7868 13176 7880
rect 13131 7840 13176 7868
rect 11149 7831 11207 7837
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 11164 7800 11192 7831
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 16666 7868 16672 7880
rect 16627 7840 16672 7868
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 16758 7828 16764 7880
rect 16816 7868 16822 7880
rect 16816 7840 16861 7868
rect 16816 7828 16822 7840
rect 10928 7772 11192 7800
rect 10928 7760 10934 7772
rect 14550 7760 14556 7812
rect 14608 7800 14614 7812
rect 17236 7800 17264 7899
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 18932 7840 19349 7868
rect 18932 7828 18938 7840
rect 19337 7837 19349 7840
rect 19383 7837 19395 7871
rect 20254 7868 20260 7880
rect 20215 7840 20260 7868
rect 19337 7831 19395 7837
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 20438 7868 20444 7880
rect 20399 7840 20444 7868
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 14608 7772 17264 7800
rect 14608 7760 14614 7772
rect 10134 7732 10140 7744
rect 10047 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7732 10198 7744
rect 10686 7732 10692 7744
rect 10192 7704 10692 7732
rect 10192 7692 10198 7704
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14240 7704 14933 7732
rect 14240 7692 14246 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 14921 7695 14979 7701
rect 15473 7735 15531 7741
rect 15473 7701 15485 7735
rect 15519 7732 15531 7735
rect 16390 7732 16396 7744
rect 15519 7704 16396 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 18785 7735 18843 7741
rect 18785 7732 18797 7735
rect 18748 7704 18797 7732
rect 18748 7692 18754 7704
rect 18785 7701 18797 7704
rect 18831 7701 18843 7735
rect 18785 7695 18843 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 14461 7531 14519 7537
rect 14461 7497 14473 7531
rect 14507 7528 14519 7531
rect 14550 7528 14556 7540
rect 14507 7500 14556 7528
rect 14507 7497 14519 7500
rect 14461 7491 14519 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 16574 7528 16580 7540
rect 15120 7500 16580 7528
rect 11333 7463 11391 7469
rect 11333 7429 11345 7463
rect 11379 7460 11391 7463
rect 11698 7460 11704 7472
rect 11379 7432 11704 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 11977 7395 12035 7401
rect 10652 7364 11376 7392
rect 10652 7352 10658 7364
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 11020 7296 11253 7324
rect 11020 7284 11026 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11348 7324 11376 7364
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7392 12130 7404
rect 15120 7401 15148 7500
rect 16574 7488 16580 7500
rect 16632 7528 16638 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16632 7500 16865 7528
rect 16632 7488 16638 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 16853 7491 16911 7497
rect 15105 7395 15163 7401
rect 12124 7364 12572 7392
rect 12124 7352 12130 7364
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 11348 7296 12449 7324
rect 11241 7287 11299 7293
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12544 7324 12572 7364
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 19794 7392 19800 7404
rect 19755 7364 19800 7392
rect 15105 7355 15163 7361
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 20070 7352 20076 7404
rect 20128 7392 20134 7404
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20128 7364 20269 7392
rect 20128 7352 20134 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 12693 7327 12751 7333
rect 12693 7324 12705 7327
rect 12544 7296 12705 7324
rect 12437 7287 12495 7293
rect 12693 7293 12705 7296
rect 12739 7293 12751 7327
rect 12693 7287 12751 7293
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 13596 7296 15485 7324
rect 13596 7284 13602 7296
rect 15473 7293 15485 7296
rect 15519 7324 15531 7327
rect 16298 7324 16304 7336
rect 15519 7296 16304 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 1210 7216 1216 7268
rect 1268 7256 1274 7268
rect 12894 7256 12900 7268
rect 1268 7228 12900 7256
rect 1268 7216 1274 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 14829 7259 14887 7265
rect 14829 7225 14841 7259
rect 14875 7256 14887 7259
rect 15286 7256 15292 7268
rect 14875 7228 15292 7256
rect 14875 7225 14887 7228
rect 14829 7219 14887 7225
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 15740 7259 15798 7265
rect 15740 7225 15752 7259
rect 15786 7256 15798 7259
rect 16022 7256 16028 7268
rect 15786 7228 16028 7256
rect 15786 7225 15798 7228
rect 15740 7219 15798 7225
rect 16022 7216 16028 7228
rect 16080 7216 16086 7268
rect 16390 7216 16396 7268
rect 16448 7256 16454 7268
rect 17328 7256 17356 7287
rect 16448 7228 17356 7256
rect 16448 7216 16454 7228
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 19705 7259 19763 7265
rect 19705 7256 19717 7259
rect 18564 7228 19717 7256
rect 18564 7216 18570 7228
rect 19705 7225 19717 7228
rect 19751 7225 19763 7259
rect 19705 7219 19763 7225
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 10376 7160 11069 7188
rect 10376 7148 10382 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11698 7188 11704 7200
rect 11659 7160 11704 7188
rect 11057 7151 11115 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 11848 7160 11893 7188
rect 11848 7148 11854 7160
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13228 7160 13829 7188
rect 13228 7148 13234 7160
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 14921 7191 14979 7197
rect 14921 7157 14933 7191
rect 14967 7188 14979 7191
rect 15930 7188 15936 7200
rect 14967 7160 15936 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 16356 7160 17141 7188
rect 16356 7148 16362 7160
rect 17129 7157 17141 7160
rect 17175 7188 17187 7191
rect 17954 7188 17960 7200
rect 17175 7160 17960 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 19245 7191 19303 7197
rect 19245 7157 19257 7191
rect 19291 7188 19303 7191
rect 19426 7188 19432 7200
rect 19291 7160 19432 7188
rect 19291 7157 19303 7160
rect 19245 7151 19303 7157
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 19610 7188 19616 7200
rect 19571 7160 19616 7188
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 11756 6956 12357 6984
rect 11756 6944 11762 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 13449 6987 13507 6993
rect 13449 6953 13461 6987
rect 13495 6984 13507 6987
rect 14090 6984 14096 6996
rect 13495 6956 14096 6984
rect 13495 6953 13507 6956
rect 13449 6947 13507 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 15286 6984 15292 6996
rect 15247 6956 15292 6984
rect 15286 6944 15292 6956
rect 15344 6944 15350 6996
rect 15657 6987 15715 6993
rect 15657 6953 15669 6987
rect 15703 6984 15715 6987
rect 17402 6984 17408 6996
rect 15703 6956 17408 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 19334 6984 19340 6996
rect 19247 6956 19340 6984
rect 19334 6944 19340 6956
rect 19392 6984 19398 6996
rect 19794 6984 19800 6996
rect 19392 6956 19800 6984
rect 19392 6944 19398 6956
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 19978 6944 19984 6996
rect 20036 6944 20042 6996
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 15746 6916 15752 6928
rect 4764 6888 15752 6916
rect 4764 6876 4770 6888
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 16574 6925 16580 6928
rect 16568 6916 16580 6925
rect 16535 6888 16580 6916
rect 16568 6879 16580 6888
rect 16574 6876 16580 6879
rect 16632 6876 16638 6928
rect 16942 6876 16948 6928
rect 17000 6916 17006 6928
rect 19058 6916 19064 6928
rect 17000 6888 19064 6916
rect 17000 6876 17006 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 19996 6916 20024 6944
rect 19812 6888 20024 6916
rect 19812 6860 19840 6888
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10962 6857 10968 6860
rect 10956 6811 10968 6857
rect 11020 6848 11026 6860
rect 13814 6848 13820 6860
rect 11020 6820 11056 6848
rect 13775 6820 13820 6848
rect 10962 6808 10968 6811
rect 11020 6808 11026 6820
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 16298 6848 16304 6860
rect 16259 6820 16304 6848
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 18224 6851 18282 6857
rect 18224 6848 18236 6851
rect 17696 6820 18236 6848
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10686 6780 10692 6792
rect 10647 6752 10692 6780
rect 10229 6743 10287 6749
rect 9674 6712 9680 6724
rect 9635 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 9766 6672 9772 6724
rect 9824 6712 9830 6724
rect 10244 6712 10272 6743
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 13906 6780 13912 6792
rect 13867 6752 13912 6780
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15344 6752 15761 6780
rect 15344 6740 15350 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 12066 6712 12072 6724
rect 9824 6684 10272 6712
rect 12027 6684 12072 6712
rect 9824 6672 9830 6684
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 17696 6721 17724 6820
rect 18224 6817 18236 6820
rect 18270 6848 18282 6851
rect 18782 6848 18788 6860
rect 18270 6820 18788 6848
rect 18270 6817 18282 6820
rect 18224 6811 18282 6817
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 19794 6808 19800 6860
rect 19852 6808 19858 6860
rect 19978 6848 19984 6860
rect 19939 6820 19984 6848
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 17954 6780 17960 6792
rect 17915 6752 17960 6780
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 20073 6783 20131 6789
rect 20073 6780 20085 6783
rect 19484 6752 20085 6780
rect 19484 6740 19490 6752
rect 20073 6749 20085 6752
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 20220 6752 20265 6780
rect 20220 6740 20226 6752
rect 17681 6715 17739 6721
rect 17681 6681 17693 6715
rect 17727 6681 17739 6715
rect 17681 6675 17739 6681
rect 19613 6715 19671 6721
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 19702 6712 19708 6724
rect 19659 6684 19708 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 17494 6604 17500 6656
rect 17552 6644 17558 6656
rect 19242 6644 19248 6656
rect 17552 6616 19248 6644
rect 17552 6604 17558 6616
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7558 6440 7564 6452
rect 6871 6412 7564 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 9217 6443 9275 6449
rect 9217 6409 9229 6443
rect 9263 6440 9275 6443
rect 9766 6440 9772 6452
rect 9263 6412 9772 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 10873 6443 10931 6449
rect 10873 6409 10885 6443
rect 10919 6440 10931 6443
rect 10962 6440 10968 6452
rect 10919 6412 10968 6440
rect 10919 6409 10931 6412
rect 10873 6403 10931 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11790 6440 11796 6452
rect 11195 6412 11796 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13814 6440 13820 6452
rect 13219 6412 13820 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 16298 6440 16304 6452
rect 14660 6412 16304 6440
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 10980 6304 11008 6400
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 10980 6276 11713 6304
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13412 6276 13737 6304
rect 13412 6264 13418 6276
rect 13725 6273 13737 6276
rect 13771 6304 13783 6307
rect 14182 6304 14188 6316
rect 13771 6276 14188 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 14660 6313 14688 6412
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 19150 6440 19156 6452
rect 18012 6412 19156 6440
rect 18012 6400 18018 6412
rect 17310 6372 17316 6384
rect 17052 6344 17316 6372
rect 17052 6313 17080 6344
rect 17310 6332 17316 6344
rect 17368 6332 17374 6384
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6273 17095 6307
rect 17402 6304 17408 6316
rect 17363 6276 17408 6304
rect 17037 6267 17095 6273
rect 9766 6245 9772 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 7883 6208 9505 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 9493 6205 9505 6208
rect 9539 6205 9551 6239
rect 9760 6236 9772 6245
rect 9727 6208 9772 6236
rect 9493 6199 9551 6205
rect 9760 6199 9772 6208
rect 8104 6171 8162 6177
rect 8104 6137 8116 6171
rect 8150 6168 8162 6171
rect 8754 6168 8760 6180
rect 8150 6140 8760 6168
rect 8150 6137 8162 6140
rect 8104 6131 8162 6137
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 9508 6168 9536 6199
rect 9766 6196 9772 6199
rect 9824 6196 9830 6248
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 14912 6239 14970 6245
rect 12492 6208 14780 6236
rect 12492 6196 12498 6208
rect 10686 6168 10692 6180
rect 9508 6140 10692 6168
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 12894 6128 12900 6180
rect 12952 6168 12958 6180
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 12952 6140 13645 6168
rect 12952 6128 12958 6140
rect 13633 6137 13645 6140
rect 13679 6137 13691 6171
rect 14752 6168 14780 6208
rect 14912 6205 14924 6239
rect 14958 6236 14970 6239
rect 17052 6236 17080 6267
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 18800 6313 18828 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 19702 6440 19708 6452
rect 19576 6412 19708 6440
rect 19576 6400 19582 6412
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 14958 6208 17080 6236
rect 19052 6239 19110 6245
rect 14958 6205 14970 6208
rect 14912 6199 14970 6205
rect 19052 6205 19064 6239
rect 19098 6236 19110 6239
rect 19334 6236 19340 6248
rect 19098 6208 19340 6236
rect 19098 6205 19110 6208
rect 19052 6199 19110 6205
rect 19334 6196 19340 6208
rect 19392 6196 19398 6248
rect 20530 6236 20536 6248
rect 20491 6208 20536 6236
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 16853 6171 16911 6177
rect 16853 6168 16865 6171
rect 14752 6140 16865 6168
rect 13633 6131 13691 6137
rect 16853 6137 16865 6140
rect 16899 6168 16911 6171
rect 18874 6168 18880 6180
rect 16899 6140 18880 6168
rect 16899 6137 16911 6140
rect 16853 6131 16911 6137
rect 18874 6128 18880 6140
rect 18932 6128 18938 6180
rect 7190 6100 7196 6112
rect 7151 6072 7196 6100
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7340 6072 7385 6100
rect 7340 6060 7346 6072
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11112 6072 11529 6100
rect 11112 6060 11118 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 12342 6100 12348 6112
rect 11664 6072 12348 6100
rect 11664 6060 11670 6072
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13538 6100 13544 6112
rect 13499 6072 13544 6100
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 16022 6100 16028 6112
rect 15983 6072 16028 6100
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16761 6103 16819 6109
rect 16761 6069 16773 6103
rect 16807 6100 16819 6103
rect 17126 6100 17132 6112
rect 16807 6072 17132 6100
rect 16807 6069 16819 6072
rect 16761 6063 16819 6069
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 19150 6100 19156 6112
rect 18371 6072 19156 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 19150 6060 19156 6072
rect 19208 6060 19214 6112
rect 20162 6100 20168 6112
rect 20123 6072 20168 6100
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 20714 6100 20720 6112
rect 20675 6072 20720 6100
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 7248 5868 9045 5896
rect 7248 5856 7254 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 10042 5896 10048 5908
rect 9723 5868 10048 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 11146 5896 11152 5908
rect 10459 5868 11152 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 11256 5868 15669 5896
rect 5988 5831 6046 5837
rect 5988 5797 6000 5831
rect 6034 5828 6046 5831
rect 6034 5800 9536 5828
rect 6034 5797 6046 5800
rect 5988 5791 6046 5797
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 5767 5732 6868 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6840 5704 6868 5732
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7644 5763 7702 5769
rect 7644 5760 7656 5763
rect 7524 5732 7656 5760
rect 7524 5720 7530 5732
rect 7644 5729 7656 5732
rect 7690 5760 7702 5763
rect 8202 5760 8208 5772
rect 7690 5732 8208 5760
rect 7690 5729 7702 5732
rect 7644 5723 7702 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 6880 5664 7389 5692
rect 6880 5652 6886 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 8754 5624 8760 5636
rect 8715 5596 8760 5624
rect 8754 5584 8760 5596
rect 8812 5584 8818 5636
rect 9508 5624 9536 5800
rect 10502 5788 10508 5840
rect 10560 5828 10566 5840
rect 11256 5828 11284 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 16758 5896 16764 5908
rect 16671 5868 16764 5896
rect 15657 5859 15715 5865
rect 16758 5856 16764 5868
rect 16816 5896 16822 5908
rect 17494 5896 17500 5908
rect 16816 5868 17500 5896
rect 16816 5856 16822 5868
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 17865 5899 17923 5905
rect 17865 5865 17877 5899
rect 17911 5896 17923 5899
rect 18506 5896 18512 5908
rect 17911 5868 18512 5896
rect 17911 5865 17923 5868
rect 17865 5859 17923 5865
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19150 5856 19156 5908
rect 19208 5896 19214 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 19208 5868 19257 5896
rect 19208 5856 19214 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19245 5859 19303 5865
rect 10560 5800 11284 5828
rect 11692 5831 11750 5837
rect 10560 5788 10566 5800
rect 11692 5797 11704 5831
rect 11738 5828 11750 5831
rect 11738 5800 13676 5828
rect 11738 5797 11750 5800
rect 11692 5791 11750 5797
rect 10318 5760 10324 5772
rect 10279 5732 10324 5760
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11146 5760 11152 5772
rect 10827 5732 11152 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 13354 5769 13360 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 11440 5732 13093 5760
rect 10870 5692 10876 5704
rect 10831 5664 10876 5692
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11440 5701 11468 5732
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13348 5760 13360 5769
rect 13315 5732 13360 5760
rect 13081 5723 13139 5729
rect 13348 5723 13360 5732
rect 13354 5720 13360 5723
rect 13412 5720 13418 5772
rect 13648 5760 13676 5800
rect 15562 5788 15568 5840
rect 15620 5828 15626 5840
rect 19337 5831 19395 5837
rect 19337 5828 19349 5831
rect 15620 5800 19349 5828
rect 15620 5788 15626 5800
rect 19337 5797 19349 5800
rect 19383 5797 19395 5831
rect 19337 5791 19395 5797
rect 14090 5760 14096 5772
rect 13648 5732 14096 5760
rect 14090 5720 14096 5732
rect 14148 5760 14154 5772
rect 15749 5763 15807 5769
rect 14148 5732 14504 5760
rect 14148 5720 14154 5732
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 10778 5624 10784 5636
rect 9508 5596 10784 5624
rect 10778 5584 10784 5596
rect 10836 5624 10842 5636
rect 10980 5624 11008 5655
rect 10836 5596 11008 5624
rect 10836 5584 10842 5596
rect 7098 5556 7104 5568
rect 7059 5528 7104 5556
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10137 5559 10195 5565
rect 10137 5556 10149 5559
rect 10100 5528 10149 5556
rect 10100 5516 10106 5528
rect 10137 5525 10149 5528
rect 10183 5556 10195 5559
rect 11440 5556 11468 5655
rect 14476 5633 14504 5732
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 16482 5760 16488 5772
rect 15795 5732 16488 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 14461 5627 14519 5633
rect 14461 5593 14473 5627
rect 14507 5593 14519 5627
rect 15286 5624 15292 5636
rect 15247 5596 15292 5624
rect 14461 5587 14519 5593
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 15948 5624 15976 5655
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 16684 5692 16712 5723
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 16908 5732 18245 5760
rect 16908 5720 16914 5732
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 19242 5720 19248 5772
rect 19300 5760 19306 5772
rect 19518 5760 19524 5772
rect 19300 5732 19524 5760
rect 19300 5720 19306 5732
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 16172 5664 16712 5692
rect 16945 5695 17003 5701
rect 16172 5652 16178 5664
rect 16945 5661 16957 5695
rect 16991 5692 17003 5695
rect 17310 5692 17316 5704
rect 16991 5664 17316 5692
rect 16991 5661 17003 5664
rect 16945 5655 17003 5661
rect 16960 5624 16988 5655
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 18325 5695 18383 5701
rect 18325 5692 18337 5695
rect 17736 5664 18337 5692
rect 17736 5652 17742 5664
rect 18325 5661 18337 5664
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 18782 5692 18788 5704
rect 18555 5664 18788 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 19484 5664 19529 5692
rect 19484 5652 19490 5664
rect 15948 5596 16988 5624
rect 18877 5627 18935 5633
rect 18877 5593 18889 5627
rect 18923 5624 18935 5627
rect 19978 5624 19984 5636
rect 18923 5596 19984 5624
rect 18923 5593 18935 5596
rect 18877 5587 18935 5593
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 10183 5528 11468 5556
rect 10183 5525 10195 5528
rect 10137 5519 10195 5525
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 11664 5528 12817 5556
rect 11664 5516 11670 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 16298 5556 16304 5568
rect 16259 5528 16304 5556
rect 12805 5519 12863 5525
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 20441 5559 20499 5565
rect 20441 5556 20453 5559
rect 19484 5528 20453 5556
rect 19484 5516 19490 5528
rect 20441 5525 20453 5528
rect 20487 5525 20499 5559
rect 20441 5519 20499 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8665 5355 8723 5361
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 10134 5352 10140 5364
rect 8711 5324 10140 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 10836 5324 11529 5352
rect 10836 5312 10842 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13964 5324 14013 5352
rect 13964 5312 13970 5324
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 15930 5352 15936 5364
rect 15891 5324 15936 5352
rect 14001 5315 14059 5321
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18598 5352 18604 5364
rect 18095 5324 18604 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 19610 5352 19616 5364
rect 19571 5324 19616 5352
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 16022 5244 16028 5296
rect 16080 5284 16086 5296
rect 16080 5256 16528 5284
rect 16080 5244 16086 5256
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8812 5188 9229 5216
rect 8812 5176 8818 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 11204 5188 11805 5216
rect 11204 5176 11210 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 11793 5179 11851 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 14182 5176 14188 5228
rect 14240 5216 14246 5228
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 14240 5188 14565 5216
rect 14240 5176 14246 5188
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 16500 5225 16528 5256
rect 19150 5244 19156 5296
rect 19208 5284 19214 5296
rect 20809 5287 20867 5293
rect 20809 5284 20821 5287
rect 19208 5256 20821 5284
rect 19208 5244 19214 5256
rect 20809 5253 20821 5256
rect 20855 5253 20867 5287
rect 20809 5247 20867 5253
rect 16393 5219 16451 5225
rect 16393 5216 16405 5219
rect 16356 5188 16405 5216
rect 16356 5176 16362 5188
rect 16393 5185 16405 5188
rect 16439 5185 16451 5219
rect 16393 5179 16451 5185
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 17828 5188 18613 5216
rect 17828 5176 17834 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 18782 5176 18788 5228
rect 18840 5216 18846 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 18840 5188 20177 5216
rect 18840 5176 18846 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7098 5157 7104 5160
rect 7092 5148 7104 5157
rect 7059 5120 7104 5148
rect 7092 5111 7104 5120
rect 7098 5108 7104 5111
rect 7156 5108 7162 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10042 5148 10048 5160
rect 9732 5120 10048 5148
rect 9732 5108 9738 5120
rect 10042 5108 10048 5120
rect 10100 5148 10106 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10100 5120 10149 5148
rect 10100 5108 10106 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14332 5120 14381 5148
rect 14332 5108 14338 5120
rect 14369 5117 14381 5120
rect 14415 5148 14427 5151
rect 16574 5148 16580 5160
rect 14415 5120 16580 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 19058 5148 19064 5160
rect 19019 5120 19064 5148
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 19242 5108 19248 5160
rect 19300 5148 19306 5160
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19300 5120 19993 5148
rect 19300 5108 19306 5120
rect 19981 5117 19993 5120
rect 20027 5117 20039 5151
rect 20622 5148 20628 5160
rect 20583 5120 20628 5148
rect 19981 5111 20039 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 10404 5083 10462 5089
rect 10404 5049 10416 5083
rect 10450 5080 10462 5083
rect 11606 5080 11612 5092
rect 10450 5052 11612 5080
rect 10450 5049 10462 5052
rect 10404 5043 10462 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 16301 5083 16359 5089
rect 16301 5049 16313 5083
rect 16347 5080 16359 5083
rect 16390 5080 16396 5092
rect 16347 5052 16396 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 18012 5052 18429 5080
rect 18012 5040 18018 5052
rect 18417 5049 18429 5052
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 18509 5083 18567 5089
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 19702 5080 19708 5092
rect 18555 5052 19708 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 19702 5040 19708 5052
rect 19760 5040 19766 5092
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 8352 4984 9045 5012
rect 8352 4972 8358 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 9180 4984 9225 5012
rect 9180 4972 9186 4984
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 14240 4984 14473 5012
rect 14240 4972 14246 4984
rect 14461 4981 14473 4984
rect 14507 5012 14519 5015
rect 16758 5012 16764 5024
rect 14507 4984 16764 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 19245 5015 19303 5021
rect 19245 4981 19257 5015
rect 19291 5012 19303 5015
rect 19886 5012 19892 5024
rect 19291 4984 19892 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 19886 4972 19892 4984
rect 19944 4972 19950 5024
rect 20073 5015 20131 5021
rect 20073 4981 20085 5015
rect 20119 5012 20131 5015
rect 20990 5012 20996 5024
rect 20119 4984 20996 5012
rect 20119 4981 20131 4984
rect 20073 4975 20131 4981
rect 20990 4972 20996 4984
rect 21048 4972 21054 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 7282 4808 7288 4820
rect 7147 4780 7288 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 9858 4808 9864 4820
rect 8619 4780 9864 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4808 10655 4811
rect 10870 4808 10876 4820
rect 10643 4780 10876 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 14185 4811 14243 4817
rect 14185 4777 14197 4811
rect 14231 4808 14243 4811
rect 14274 4808 14280 4820
rect 14231 4780 14280 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 19334 4768 19340 4820
rect 19392 4768 19398 4820
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 8941 4743 8999 4749
rect 8941 4740 8953 4743
rect 7064 4712 8953 4740
rect 7064 4700 7070 4712
rect 8941 4709 8953 4712
rect 8987 4709 8999 4743
rect 8941 4703 8999 4709
rect 9033 4743 9091 4749
rect 9033 4709 9045 4743
rect 9079 4740 9091 4743
rect 9122 4740 9128 4752
rect 9079 4712 9128 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 9122 4700 9128 4712
rect 9180 4740 9186 4752
rect 16390 4740 16396 4752
rect 9180 4712 16396 4740
rect 9180 4700 9186 4712
rect 16390 4700 16396 4712
rect 16448 4740 16454 4752
rect 16850 4740 16856 4752
rect 16448 4712 16856 4740
rect 16448 4700 16454 4712
rect 16850 4700 16856 4712
rect 16908 4700 16914 4752
rect 17304 4743 17362 4749
rect 17304 4709 17316 4743
rect 17350 4740 17362 4743
rect 19352 4740 19380 4768
rect 17350 4712 19380 4740
rect 19420 4743 19478 4749
rect 17350 4709 17362 4712
rect 17304 4703 17362 4709
rect 19420 4709 19432 4743
rect 19466 4740 19478 4743
rect 20162 4740 20168 4752
rect 19466 4712 20168 4740
rect 19466 4709 19478 4712
rect 19420 4703 19478 4709
rect 20162 4700 20168 4712
rect 20220 4700 20226 4752
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 5224 4644 7481 4672
rect 5224 4632 5230 4644
rect 7469 4641 7481 4644
rect 7515 4641 7527 4675
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 7469 4635 7527 4641
rect 7760 4644 10977 4672
rect 7558 4604 7564 4616
rect 7519 4576 7564 4604
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7668 4536 7696 4567
rect 7156 4508 7696 4536
rect 7156 4496 7162 4508
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 7760 4468 7788 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 11103 4644 13645 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 9088 4576 9137 4604
rect 9088 4564 9094 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9582 4496 9588 4548
rect 9640 4496 9646 4548
rect 10962 4496 10968 4548
rect 11020 4536 11026 4548
rect 11072 4536 11100 4635
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 14240 4644 14289 4672
rect 14240 4632 14246 4644
rect 14277 4641 14289 4644
rect 14323 4641 14335 4675
rect 16114 4672 16120 4684
rect 14277 4635 14335 4641
rect 14384 4644 16120 4672
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 11606 4604 11612 4616
rect 11287 4576 11612 4604
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 14384 4604 14412 4644
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16264 4644 17049 4672
rect 16264 4632 16270 4644
rect 17037 4641 17049 4644
rect 17083 4672 17095 4675
rect 18598 4672 18604 4684
rect 17083 4644 18604 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 18598 4632 18604 4644
rect 18656 4672 18662 4684
rect 19153 4675 19211 4681
rect 19153 4672 19165 4675
rect 18656 4644 19165 4672
rect 18656 4632 18662 4644
rect 19153 4641 19165 4644
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 12268 4576 14412 4604
rect 14461 4607 14519 4613
rect 11020 4508 11100 4536
rect 11020 4496 11026 4508
rect 5500 4440 7788 4468
rect 9600 4468 9628 4496
rect 12268 4468 12296 4576
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 14550 4604 14556 4616
rect 14507 4576 14556 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 13633 4539 13691 4545
rect 13633 4505 13645 4539
rect 13679 4536 13691 4539
rect 13679 4508 13952 4536
rect 13679 4505 13691 4508
rect 13633 4499 13691 4505
rect 13814 4468 13820 4480
rect 9600 4440 12296 4468
rect 13775 4440 13820 4468
rect 5500 4428 5506 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 13924 4468 13952 4508
rect 17678 4468 17684 4480
rect 13924 4440 17684 4468
rect 17678 4428 17684 4440
rect 17736 4428 17742 4480
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 17828 4440 18429 4468
rect 17828 4428 17834 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 20530 4468 20536 4480
rect 20491 4440 20536 4468
rect 18417 4431 18475 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 9030 4224 9036 4276
rect 9088 4264 9094 4276
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 9088 4236 9229 4264
rect 9088 4224 9094 4236
rect 9217 4233 9229 4236
rect 9263 4233 9275 4267
rect 9217 4227 9275 4233
rect 15212 4236 16252 4264
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 10870 4128 10876 4140
rect 9456 4100 10732 4128
rect 10831 4100 10876 4128
rect 9456 4088 9462 4100
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 6880 4032 7849 4060
rect 6880 4020 6886 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 7852 3992 7880 4023
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 10410 4060 10416 4072
rect 8720 4032 10416 4060
rect 8720 4020 8726 4032
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 8104 3995 8162 4001
rect 7852 3964 8064 3992
rect 8036 3924 8064 3964
rect 8104 3961 8116 3995
rect 8150 3992 8162 3995
rect 8570 3992 8576 4004
rect 8150 3964 8576 3992
rect 8150 3961 8162 3964
rect 8104 3955 8162 3961
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 10597 3995 10655 4001
rect 10597 3992 10609 3995
rect 9815 3964 10609 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10597 3961 10609 3964
rect 10643 3961 10655 3995
rect 10704 3992 10732 4100
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12894 4128 12900 4140
rect 12400 4100 12900 4128
rect 12400 4088 12406 4100
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13170 4088 13176 4140
rect 13228 4128 13234 4140
rect 13228 4100 13952 4128
rect 13228 4088 13234 4100
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13814 4060 13820 4072
rect 13035 4032 13820 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 13924 4060 13952 4100
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14332 4100 14657 4128
rect 14332 4088 14338 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 15212 4128 15240 4236
rect 14645 4091 14703 4097
rect 14752 4100 15240 4128
rect 16224 4128 16252 4236
rect 18064 4236 19288 4264
rect 18064 4128 18092 4236
rect 19260 4196 19288 4236
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 19392 4236 19441 4264
rect 19392 4224 19398 4236
rect 19429 4233 19441 4236
rect 19475 4233 19487 4267
rect 19702 4264 19708 4276
rect 19663 4236 19708 4264
rect 19429 4227 19487 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 19610 4196 19616 4208
rect 19260 4168 19616 4196
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 16224 4100 18092 4128
rect 14752 4060 14780 4100
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 19392 4100 20269 4128
rect 19392 4088 19398 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 22462 4128 22468 4140
rect 20956 4100 22468 4128
rect 20956 4088 20962 4100
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 15194 4060 15200 4072
rect 13924 4032 14780 4060
rect 15155 4032 15200 4060
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15464 4063 15522 4069
rect 15464 4029 15476 4063
rect 15510 4060 15522 4063
rect 17770 4060 17776 4072
rect 15510 4032 17776 4060
rect 15510 4029 15522 4032
rect 15464 4023 15522 4029
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18598 4060 18604 4072
rect 18095 4032 18604 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 18782 4020 18788 4072
rect 18840 4060 18846 4072
rect 19426 4060 19432 4072
rect 18840 4032 19432 4060
rect 18840 4020 18846 4032
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20404 4032 20729 4060
rect 20404 4020 20410 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 13722 3992 13728 4004
rect 10704 3964 13728 3992
rect 10597 3955 10655 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 18294 3995 18352 4001
rect 18294 3992 18306 3995
rect 18064 3964 18306 3992
rect 18064 3936 18092 3964
rect 18294 3961 18306 3964
rect 18340 3961 18352 3995
rect 18294 3955 18352 3961
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 18472 3964 20944 3992
rect 18472 3952 18478 3964
rect 9674 3924 9680 3936
rect 8036 3896 9680 3924
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10686 3924 10692 3936
rect 10647 3896 10692 3924
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11756 3896 11805 3924
rect 11756 3884 11762 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11793 3887 11851 3893
rect 12529 3927 12587 3933
rect 12529 3893 12541 3927
rect 12575 3924 12587 3927
rect 12618 3924 12624 3936
rect 12575 3896 12624 3924
rect 12575 3893 12587 3896
rect 12529 3887 12587 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12768 3896 12909 3924
rect 12768 3884 12774 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 14093 3927 14151 3933
rect 14093 3924 14105 3927
rect 14056 3896 14105 3924
rect 14056 3884 14062 3896
rect 14093 3893 14105 3896
rect 14139 3893 14151 3927
rect 14458 3924 14464 3936
rect 14419 3896 14464 3924
rect 14093 3887 14151 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3924 14611 3927
rect 15102 3924 15108 3936
rect 14599 3896 15108 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 16206 3924 16212 3936
rect 15252 3896 16212 3924
rect 15252 3884 15258 3896
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 16482 3884 16488 3936
rect 16540 3924 16546 3936
rect 16577 3927 16635 3933
rect 16577 3924 16589 3927
rect 16540 3896 16589 3924
rect 16540 3884 16546 3896
rect 16577 3893 16589 3896
rect 16623 3893 16635 3927
rect 17494 3924 17500 3936
rect 17455 3896 17500 3924
rect 16577 3887 16635 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 18046 3884 18052 3936
rect 18104 3884 18110 3936
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20916 3933 20944 3964
rect 20901 3927 20959 3933
rect 20220 3896 20265 3924
rect 20220 3884 20226 3896
rect 20901 3893 20913 3927
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 8294 3720 8300 3732
rect 2372 3692 8300 3720
rect 2372 3680 2378 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8570 3720 8576 3732
rect 8531 3692 8576 3720
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 12250 3720 12256 3732
rect 8680 3692 12256 3720
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 5166 3652 5172 3664
rect 2924 3624 5172 3652
rect 2924 3612 2930 3624
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 8680 3652 8708 3692
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 12713 3723 12771 3729
rect 12713 3689 12725 3723
rect 12759 3720 12771 3723
rect 13078 3720 13084 3732
rect 12759 3692 13084 3720
rect 12759 3689 12771 3692
rect 12713 3683 12771 3689
rect 5552 3624 8708 3652
rect 9944 3655 10002 3661
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 5442 3584 5448 3596
rect 3476 3556 5448 3584
rect 3476 3544 3482 3556
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 5552 3516 5580 3624
rect 9944 3621 9956 3655
rect 9990 3652 10002 3655
rect 12728 3652 12756 3683
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 13780 3692 17877 3720
rect 13780 3680 13786 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 18230 3680 18236 3732
rect 18288 3720 18294 3732
rect 19429 3723 19487 3729
rect 18288 3692 19380 3720
rect 18288 3680 18294 3692
rect 9990 3624 12756 3652
rect 9990 3621 10002 3624
rect 9944 3615 10002 3621
rect 18046 3612 18052 3664
rect 18104 3652 18110 3664
rect 18104 3624 18184 3652
rect 18104 3612 18110 3624
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6880 3556 7205 3584
rect 6880 3544 6886 3556
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 7460 3587 7518 3593
rect 7460 3553 7472 3587
rect 7506 3584 7518 3587
rect 8202 3584 8208 3596
rect 7506 3556 8208 3584
rect 7506 3553 7518 3556
rect 7460 3547 7518 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9674 3584 9680 3596
rect 9587 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 9732 3556 11345 3584
rect 9732 3544 9738 3556
rect 11333 3553 11345 3556
rect 11379 3584 11391 3587
rect 11422 3584 11428 3596
rect 11379 3556 11428 3584
rect 11379 3553 11391 3556
rect 11333 3547 11391 3553
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 11600 3587 11658 3593
rect 11600 3553 11612 3587
rect 11646 3584 11658 3587
rect 11974 3584 11980 3596
rect 11646 3556 11980 3584
rect 11646 3553 11658 3556
rect 11600 3547 11658 3553
rect 11974 3544 11980 3556
rect 12032 3584 12038 3596
rect 13532 3587 13590 3593
rect 12032 3556 12388 3584
rect 12032 3544 12038 3556
rect 8846 3516 8852 3528
rect 4028 3488 5580 3516
rect 8807 3488 8852 3516
rect 4028 3476 4034 3488
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 12360 3516 12388 3556
rect 13532 3553 13544 3587
rect 13578 3584 13590 3587
rect 14274 3584 14280 3596
rect 13578 3556 14280 3584
rect 13578 3553 13590 3556
rect 13532 3547 13590 3553
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15252 3556 15301 3584
rect 15252 3544 15258 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15556 3587 15614 3593
rect 15556 3553 15568 3587
rect 15602 3584 15614 3587
rect 16482 3584 16488 3596
rect 15602 3556 16488 3584
rect 15602 3553 15614 3556
rect 15556 3547 15614 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 12360 3488 12480 3516
rect 12452 3448 12480 3488
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13044 3488 13277 3516
rect 13044 3476 13050 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 16632 3488 17969 3516
rect 16632 3476 16638 3488
rect 17957 3485 17969 3488
rect 18003 3516 18015 3519
rect 18046 3516 18052 3528
rect 18003 3488 18052 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18156 3525 18184 3624
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 18932 3624 19012 3652
rect 18932 3612 18938 3624
rect 18690 3584 18696 3596
rect 18651 3556 18696 3584
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18874 3516 18880 3528
rect 18835 3488 18880 3516
rect 18141 3479 18199 3485
rect 12452 3420 13207 3448
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 10594 3380 10600 3392
rect 5684 3352 10600 3380
rect 5684 3340 5690 3352
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10836 3352 11069 3380
rect 10836 3340 10842 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11057 3343 11115 3349
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 13078 3380 13084 3392
rect 11204 3352 13084 3380
rect 11204 3340 11210 3352
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 13179 3380 13207 3420
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 14645 3451 14703 3457
rect 14645 3448 14657 3451
rect 14608 3420 14657 3448
rect 14608 3408 14614 3420
rect 14645 3417 14657 3420
rect 14691 3417 14703 3451
rect 18156 3448 18184 3479
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 18984 3516 19012 3624
rect 19352 3593 19380 3692
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 20070 3720 20076 3732
rect 19475 3692 20076 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 19702 3612 19708 3664
rect 19760 3652 19766 3664
rect 20714 3652 20720 3664
rect 19760 3624 20720 3652
rect 19760 3612 19766 3624
rect 20714 3612 20720 3624
rect 20772 3612 20778 3664
rect 19337 3587 19395 3593
rect 19337 3553 19349 3587
rect 19383 3584 19395 3587
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19383 3556 19809 3584
rect 19383 3553 19395 3556
rect 19337 3547 19395 3553
rect 19797 3553 19809 3556
rect 19843 3553 19855 3587
rect 20622 3584 20628 3596
rect 19797 3547 19855 3553
rect 19904 3556 20628 3584
rect 19904 3525 19932 3556
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 19889 3519 19947 3525
rect 19889 3516 19901 3519
rect 18984 3488 19901 3516
rect 19889 3485 19901 3488
rect 19935 3485 19947 3519
rect 20070 3516 20076 3528
rect 19983 3488 20076 3516
rect 19889 3479 19947 3485
rect 20070 3476 20076 3488
rect 20128 3516 20134 3528
rect 20530 3516 20536 3528
rect 20128 3488 20536 3516
rect 20128 3476 20134 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20088 3448 20116 3476
rect 18156 3420 20116 3448
rect 14645 3411 14703 3417
rect 14568 3380 14596 3408
rect 13179 3352 14596 3380
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 15988 3352 16681 3380
rect 15988 3340 15994 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16669 3343 16727 3349
rect 17497 3383 17555 3389
rect 17497 3349 17509 3383
rect 17543 3380 17555 3383
rect 18506 3380 18512 3392
rect 17543 3352 18512 3380
rect 17543 3349 17555 3352
rect 17497 3343 17555 3349
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 18690 3340 18696 3392
rect 18748 3380 18754 3392
rect 18966 3380 18972 3392
rect 18748 3352 18972 3380
rect 18748 3340 18754 3352
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 19337 3383 19395 3389
rect 19337 3349 19349 3383
rect 19383 3380 19395 3383
rect 20530 3380 20536 3392
rect 19383 3352 20536 3380
rect 19383 3349 19395 3352
rect 19337 3343 19395 3349
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 8202 3176 8208 3188
rect 6144 3148 7788 3176
rect 8163 3148 8208 3176
rect 6144 3136 6150 3148
rect 7760 3108 7788 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8478 3176 8484 3188
rect 8439 3148 8484 3176
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 10870 3176 10876 3188
rect 9600 3148 10876 3176
rect 8386 3108 8392 3120
rect 7760 3080 8392 3108
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 9600 3108 9628 3148
rect 10870 3136 10876 3148
rect 10928 3176 10934 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10928 3148 10977 3176
rect 10928 3136 10934 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 12710 3176 12716 3188
rect 11379 3148 12716 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 14274 3176 14280 3188
rect 12912 3148 13860 3176
rect 14235 3148 14280 3176
rect 8496 3080 9628 3108
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 7092 2975 7150 2981
rect 1820 2944 6040 2972
rect 1820 2932 1826 2944
rect 6012 2836 6040 2944
rect 7092 2941 7104 2975
rect 7138 2972 7150 2975
rect 8496 2972 8524 3080
rect 10594 3068 10600 3120
rect 10652 3108 10658 3120
rect 12912 3108 12940 3148
rect 10652 3080 12940 3108
rect 13832 3108 13860 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14369 3179 14427 3185
rect 14369 3145 14381 3179
rect 14415 3176 14427 3179
rect 14737 3179 14795 3185
rect 14737 3176 14749 3179
rect 14415 3148 14749 3176
rect 14415 3145 14427 3148
rect 14369 3139 14427 3145
rect 14737 3145 14749 3148
rect 14783 3145 14795 3179
rect 15102 3176 15108 3188
rect 15063 3148 15108 3176
rect 14737 3139 14795 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 16172 3148 17785 3176
rect 16172 3136 16178 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 19429 3179 19487 3185
rect 19429 3145 19441 3179
rect 19475 3176 19487 3179
rect 20162 3176 20168 3188
rect 19475 3148 20168 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 15010 3108 15016 3120
rect 13832 3080 15016 3108
rect 10652 3068 10658 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 16022 3068 16028 3120
rect 16080 3108 16086 3120
rect 20717 3111 20775 3117
rect 20717 3108 20729 3111
rect 16080 3080 20729 3108
rect 16080 3068 16086 3080
rect 20717 3077 20729 3080
rect 20763 3077 20775 3111
rect 20717 3071 20775 3077
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8628 3012 9045 3040
rect 8628 3000 8634 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11974 3040 11980 3052
rect 11664 3012 11836 3040
rect 11935 3012 11980 3040
rect 11664 3000 11670 3012
rect 8846 2972 8852 2984
rect 7138 2944 8524 2972
rect 8807 2944 8852 2972
rect 7138 2941 7150 2944
rect 7092 2935 7150 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9585 2975 9643 2981
rect 8996 2944 9041 2972
rect 8996 2932 9002 2944
rect 9585 2941 9597 2975
rect 9631 2972 9643 2975
rect 9674 2972 9680 2984
rect 9631 2944 9680 2972
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9852 2975 9910 2981
rect 9852 2941 9864 2975
rect 9898 2972 9910 2975
rect 10778 2972 10784 2984
rect 9898 2944 10784 2972
rect 9898 2941 9910 2944
rect 9852 2935 9910 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11698 2972 11704 2984
rect 11659 2944 11704 2972
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 11808 2972 11836 3012
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 13924 3012 15761 3040
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 11808 2944 12909 2972
rect 12897 2941 12909 2944
rect 12943 2972 12955 2975
rect 12986 2972 12992 2984
rect 12943 2944 12992 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 12986 2932 12992 2944
rect 13044 2932 13050 2984
rect 13164 2975 13222 2981
rect 13164 2941 13176 2975
rect 13210 2972 13222 2975
rect 13630 2972 13636 2984
rect 13210 2944 13636 2972
rect 13210 2941 13222 2944
rect 13164 2935 13222 2941
rect 13630 2932 13636 2944
rect 13688 2972 13694 2984
rect 13924 2972 13952 3012
rect 15749 3009 15761 3012
rect 15795 3040 15807 3043
rect 15930 3040 15936 3052
rect 15795 3012 15936 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16540 3012 16681 3040
rect 16540 3000 16546 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 17862 3040 17868 3052
rect 16669 3003 16727 3009
rect 17420 3012 17868 3040
rect 13688 2944 13952 2972
rect 14553 2975 14611 2981
rect 13688 2932 13694 2944
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 15654 2972 15660 2984
rect 14599 2944 15660 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 17034 2972 17040 2984
rect 15764 2944 17040 2972
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 11793 2907 11851 2913
rect 11793 2904 11805 2907
rect 8352 2876 11805 2904
rect 8352 2864 8358 2876
rect 11793 2873 11805 2876
rect 11839 2873 11851 2907
rect 11793 2867 11851 2873
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 14369 2907 14427 2913
rect 14369 2904 14381 2907
rect 13780 2876 14381 2904
rect 13780 2864 13786 2876
rect 14369 2873 14381 2876
rect 14415 2873 14427 2907
rect 15764 2904 15792 2944
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17420 2981 17448 3012
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 19334 3040 19340 3052
rect 18739 3012 19340 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19576 3012 19901 3040
rect 19576 3000 19582 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 19889 3003 19947 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17552 2944 18429 2972
rect 17552 2932 17558 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 20438 2932 20444 2984
rect 20496 2972 20502 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20496 2944 20545 2972
rect 20496 2932 20502 2944
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 14369 2867 14427 2873
rect 14936 2876 15792 2904
rect 11054 2836 11060 2848
rect 6012 2808 11060 2836
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12492 2808 12537 2836
rect 12492 2796 12498 2808
rect 13078 2796 13084 2848
rect 13136 2836 13142 2848
rect 14936 2836 14964 2876
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 16448 2876 16497 2904
rect 16448 2864 16454 2876
rect 16485 2873 16497 2876
rect 16531 2873 16543 2907
rect 17678 2904 17684 2916
rect 16485 2867 16543 2873
rect 16592 2876 17684 2904
rect 16592 2848 16620 2876
rect 17678 2864 17684 2876
rect 17736 2864 17742 2916
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 21358 2904 21364 2916
rect 19300 2876 21364 2904
rect 19300 2864 19306 2876
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 15470 2836 15476 2848
rect 13136 2808 14964 2836
rect 15431 2808 15476 2836
rect 13136 2796 13142 2808
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 15565 2839 15623 2845
rect 15565 2805 15577 2839
rect 15611 2836 15623 2839
rect 16117 2839 16175 2845
rect 16117 2836 16129 2839
rect 15611 2808 16129 2836
rect 15611 2805 15623 2808
rect 15565 2799 15623 2805
rect 16117 2805 16129 2808
rect 16163 2805 16175 2839
rect 16574 2836 16580 2848
rect 16535 2808 16580 2836
rect 16117 2799 16175 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 17589 2839 17647 2845
rect 17589 2836 17601 2839
rect 17092 2808 17601 2836
rect 17092 2796 17098 2808
rect 17589 2805 17601 2808
rect 17635 2805 17647 2839
rect 17589 2799 17647 2805
rect 17773 2839 17831 2845
rect 17773 2805 17785 2839
rect 17819 2836 17831 2839
rect 18966 2836 18972 2848
rect 17819 2808 18972 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 18966 2796 18972 2808
rect 19024 2836 19030 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 19024 2808 19809 2836
rect 19024 2796 19030 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 7469 2635 7527 2641
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 8938 2632 8944 2644
rect 7515 2604 8944 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10686 2632 10692 2644
rect 10183 2604 10692 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 12492 2604 13369 2632
rect 12492 2592 12498 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 13357 2595 13415 2601
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 15841 2635 15899 2641
rect 15841 2632 15853 2635
rect 15528 2604 15853 2632
rect 15528 2592 15534 2604
rect 15841 2601 15853 2604
rect 15887 2601 15899 2635
rect 15841 2595 15899 2601
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 16666 2632 16672 2644
rect 16255 2604 16672 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 16666 2592 16672 2604
rect 16724 2632 16730 2644
rect 17770 2632 17776 2644
rect 16724 2604 17776 2632
rect 16724 2592 16730 2604
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 17865 2635 17923 2641
rect 17865 2601 17877 2635
rect 17911 2632 17923 2635
rect 19242 2632 19248 2644
rect 17911 2604 19248 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20717 2635 20775 2641
rect 20717 2601 20729 2635
rect 20763 2601 20775 2635
rect 20717 2595 20775 2601
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 10505 2567 10563 2573
rect 10505 2564 10517 2567
rect 7800 2536 10517 2564
rect 7800 2524 7806 2536
rect 10505 2533 10517 2536
rect 10551 2533 10563 2567
rect 10505 2527 10563 2533
rect 10597 2567 10655 2573
rect 10597 2533 10609 2567
rect 10643 2564 10655 2567
rect 10962 2564 10968 2576
rect 10643 2536 10968 2564
rect 10643 2533 10655 2536
rect 10597 2527 10655 2533
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 20732 2564 20760 2595
rect 15436 2536 20760 2564
rect 15436 2524 15442 2536
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7248 2468 7849 2496
rect 7248 2456 7254 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11882 2496 11888 2508
rect 11471 2468 11888 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 14366 2496 14372 2508
rect 12023 2468 14372 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2496 16359 2499
rect 16942 2496 16948 2508
rect 16347 2468 16804 2496
rect 16903 2468 16948 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7616 2400 7941 2428
rect 7616 2388 7622 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 8202 2428 8208 2440
rect 8159 2400 8208 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 10778 2428 10784 2440
rect 10739 2400 10784 2428
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 10888 2400 13461 2428
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 10888 2360 10916 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13630 2428 13636 2440
rect 13591 2400 13636 2428
rect 13449 2391 13507 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 16482 2428 16488 2440
rect 16443 2400 16488 2428
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 16776 2428 16804 2468
rect 16942 2456 16948 2468
rect 17000 2456 17006 2508
rect 17218 2496 17224 2508
rect 17052 2468 17224 2496
rect 17052 2428 17080 2468
rect 17218 2456 17224 2468
rect 17276 2496 17282 2508
rect 17586 2496 17592 2508
rect 17276 2468 17592 2496
rect 17276 2456 17282 2468
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2496 17739 2499
rect 18230 2496 18236 2508
rect 17727 2468 18236 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18690 2496 18696 2508
rect 18371 2468 18696 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 18874 2496 18880 2508
rect 18835 2468 18880 2496
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19116 2468 19441 2496
rect 19116 2456 19122 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 19996 2428 20024 2459
rect 20254 2456 20260 2508
rect 20312 2496 20318 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20312 2468 20545 2496
rect 20312 2456 20318 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 21082 2428 21088 2440
rect 16776 2400 17080 2428
rect 17420 2400 19196 2428
rect 19996 2400 21088 2428
rect 8904 2332 10916 2360
rect 12989 2363 13047 2369
rect 8904 2320 8910 2332
rect 12989 2329 13001 2363
rect 13035 2360 13047 2363
rect 14458 2360 14464 2372
rect 13035 2332 14464 2360
rect 13035 2329 13047 2332
rect 12989 2323 13047 2329
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 14826 2320 14832 2372
rect 14884 2360 14890 2372
rect 17420 2360 17448 2400
rect 14884 2332 17448 2360
rect 14884 2320 14890 2332
rect 17494 2320 17500 2372
rect 17552 2360 17558 2372
rect 18509 2363 18567 2369
rect 18509 2360 18521 2363
rect 17552 2332 18521 2360
rect 17552 2320 17558 2332
rect 18509 2329 18521 2332
rect 18555 2329 18567 2363
rect 18509 2323 18567 2329
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 12618 2292 12624 2304
rect 12207 2264 12624 2292
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 16482 2252 16488 2304
rect 16540 2292 16546 2304
rect 17129 2295 17187 2301
rect 17129 2292 17141 2295
rect 16540 2264 17141 2292
rect 16540 2252 16546 2264
rect 17129 2261 17141 2264
rect 17175 2261 17187 2295
rect 17129 2255 17187 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 19061 2295 19119 2301
rect 19061 2292 19073 2295
rect 18012 2264 19073 2292
rect 18012 2252 18018 2264
rect 19061 2261 19073 2264
rect 19107 2261 19119 2295
rect 19168 2292 19196 2400
rect 21082 2388 21088 2400
rect 21140 2388 21146 2440
rect 19613 2363 19671 2369
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 20806 2360 20812 2372
rect 19659 2332 20812 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 20806 2320 20812 2332
rect 20864 2320 20870 2372
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 19168 2264 20177 2292
rect 19061 2255 19119 2261
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 9950 1776 9956 1828
rect 10008 1816 10014 1828
rect 15562 1816 15568 1828
rect 10008 1788 15568 1816
rect 10008 1776 10014 1788
rect 15562 1776 15568 1788
rect 15620 1776 15626 1828
rect 198 824 204 876
rect 256 864 262 876
rect 8662 864 8668 876
rect 256 836 8668 864
rect 256 824 262 836
rect 8662 824 8668 836
rect 8720 824 8726 876
rect 6638 552 6644 604
rect 6696 592 6702 604
rect 7006 592 7012 604
rect 6696 564 7012 592
rect 6696 552 6702 564
rect 7006 552 7012 564
rect 7064 552 7070 604
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 20628 20000 20680 20052
rect 19892 19864 19944 19916
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 5724 19252 5776 19304
rect 15936 19252 15988 19304
rect 17960 19252 18012 19304
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 17868 19116 17920 19168
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 20904 19116 20956 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 20536 18912 20588 18964
rect 15936 18887 15988 18896
rect 15936 18853 15945 18887
rect 15945 18853 15979 18887
rect 15979 18853 15988 18887
rect 15936 18844 15988 18853
rect 17960 18887 18012 18896
rect 17960 18853 17969 18887
rect 17969 18853 18003 18887
rect 18003 18853 18012 18887
rect 17960 18844 18012 18853
rect 19892 18887 19944 18896
rect 19892 18853 19901 18887
rect 19901 18853 19935 18887
rect 19935 18853 19944 18887
rect 19892 18844 19944 18853
rect 9956 18776 10008 18828
rect 11704 18776 11756 18828
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 19616 18819 19668 18828
rect 19616 18785 19625 18819
rect 19625 18785 19659 18819
rect 19659 18785 19668 18819
rect 19616 18776 19668 18785
rect 17960 18708 18012 18760
rect 19984 18572 20036 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 20168 18411 20220 18420
rect 20168 18377 20177 18411
rect 20177 18377 20211 18411
rect 20211 18377 20220 18411
rect 20168 18368 20220 18377
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 7564 18164 7616 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 17868 17824 17920 17876
rect 20444 17867 20496 17876
rect 20444 17833 20453 17867
rect 20453 17833 20487 17867
rect 20487 17833 20496 17867
rect 20444 17824 20496 17833
rect 10876 17688 10928 17740
rect 14464 17688 14516 17740
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 14464 17187 14516 17196
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 14004 17076 14056 17128
rect 19984 17119 20036 17128
rect 19984 17085 19993 17119
rect 19993 17085 20027 17119
rect 20027 17085 20036 17119
rect 19984 17076 20036 17085
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 20536 16668 20588 16720
rect 16396 16600 16448 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 19984 16056 20036 16108
rect 15384 15988 15436 16040
rect 19616 15988 19668 16040
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 19616 15444 19668 15496
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 20168 15147 20220 15156
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 9772 14943 9824 14952
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 20076 14560 20128 14612
rect 20444 14603 20496 14612
rect 20444 14569 20453 14603
rect 20453 14569 20487 14603
rect 20487 14569 20496 14603
rect 20444 14560 20496 14569
rect 8484 14424 8536 14476
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 19984 14356 20036 14408
rect 11152 14288 11204 14340
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 19248 14016 19300 14068
rect 17316 13948 17368 14000
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 10232 13812 10284 13864
rect 16120 13855 16172 13864
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 16672 13812 16724 13864
rect 19892 13855 19944 13864
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 19800 13744 19852 13796
rect 18788 13676 18840 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 19248 13515 19300 13524
rect 19248 13481 19257 13515
rect 19257 13481 19291 13515
rect 19291 13481 19300 13515
rect 19248 13472 19300 13481
rect 19708 13404 19760 13456
rect 19340 13336 19392 13388
rect 12624 13268 12676 13320
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 15660 12928 15712 12980
rect 17960 12928 18012 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 13912 12860 13964 12912
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 17500 12724 17552 12776
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 16580 12656 16632 12708
rect 19800 12656 19852 12708
rect 20260 12656 20312 12708
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 10876 12384 10928 12436
rect 11060 12384 11112 12436
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 20444 12427 20496 12436
rect 13452 12248 13504 12300
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 15292 12180 15344 12232
rect 16120 12316 16172 12368
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 16764 12248 16816 12300
rect 18604 12316 18656 12368
rect 19340 12316 19392 12368
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 20260 12291 20312 12300
rect 20260 12257 20269 12291
rect 20269 12257 20303 12291
rect 20303 12257 20312 12291
rect 20260 12248 20312 12257
rect 18604 12180 18656 12232
rect 15844 12044 15896 12096
rect 18880 12044 18932 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 15752 11840 15804 11892
rect 16764 11840 16816 11892
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 17592 11704 17644 11756
rect 13176 11679 13228 11688
rect 13176 11645 13185 11679
rect 13185 11645 13219 11679
rect 13219 11645 13228 11679
rect 13176 11636 13228 11645
rect 13360 11636 13412 11688
rect 15292 11636 15344 11688
rect 15752 11679 15804 11688
rect 15752 11645 15786 11679
rect 15786 11645 15804 11679
rect 15752 11636 15804 11645
rect 18512 11636 18564 11688
rect 20628 11704 20680 11756
rect 18696 11636 18748 11688
rect 18880 11679 18932 11688
rect 18880 11645 18914 11679
rect 18914 11645 18932 11679
rect 18880 11636 18932 11645
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 15844 11568 15896 11620
rect 19524 11568 19576 11620
rect 21916 11568 21968 11620
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 20260 11543 20312 11552
rect 20260 11509 20269 11543
rect 20269 11509 20303 11543
rect 20303 11509 20312 11543
rect 20260 11500 20312 11509
rect 20444 11500 20496 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 13176 11296 13228 11348
rect 15568 11296 15620 11348
rect 19340 11296 19392 11348
rect 9588 11228 9640 11280
rect 13176 11160 13228 11212
rect 15936 11160 15988 11212
rect 10784 11092 10836 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 4068 11024 4120 11076
rect 13452 11024 13504 11076
rect 18880 11228 18932 11280
rect 19984 11228 20036 11280
rect 16304 11160 16356 11212
rect 20628 11160 20680 11212
rect 15292 10956 15344 11008
rect 18696 11092 18748 11144
rect 17960 10956 18012 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 16580 10795 16632 10804
rect 16580 10761 16589 10795
rect 16589 10761 16623 10795
rect 16623 10761 16632 10795
rect 16580 10752 16632 10761
rect 16488 10616 16540 10668
rect 16764 10616 16816 10668
rect 17960 10616 18012 10668
rect 19984 10616 20036 10668
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 20628 10659 20680 10668
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 19340 10548 19392 10600
rect 20260 10548 20312 10600
rect 11980 10480 12032 10532
rect 15752 10523 15804 10532
rect 15752 10489 15761 10523
rect 15761 10489 15795 10523
rect 15795 10489 15804 10523
rect 15752 10480 15804 10489
rect 16672 10480 16724 10532
rect 664 10412 716 10464
rect 9588 10412 9640 10464
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 13820 10208 13872 10260
rect 15752 10208 15804 10260
rect 18420 10208 18472 10260
rect 15292 10140 15344 10192
rect 17960 10140 18012 10192
rect 19984 10140 20036 10192
rect 20444 10140 20496 10192
rect 13084 10072 13136 10124
rect 14556 10072 14608 10124
rect 15200 10072 15252 10124
rect 17592 10115 17644 10124
rect 17592 10081 17601 10115
rect 17601 10081 17635 10115
rect 17635 10081 17644 10115
rect 17592 10072 17644 10081
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 20352 10072 20404 10124
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 18972 9979 19024 9988
rect 18972 9945 18981 9979
rect 18981 9945 19015 9979
rect 19015 9945 19024 9979
rect 18972 9936 19024 9945
rect 16488 9868 16540 9920
rect 19064 9868 19116 9920
rect 19524 9868 19576 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 11888 9596 11940 9648
rect 11612 9528 11664 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 17592 9528 17644 9580
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 12440 9460 12492 9512
rect 15292 9460 15344 9512
rect 16488 9460 16540 9512
rect 18972 9460 19024 9512
rect 19248 9460 19300 9512
rect 11888 9392 11940 9444
rect 13820 9435 13872 9444
rect 13820 9401 13854 9435
rect 13854 9401 13872 9435
rect 13820 9392 13872 9401
rect 11060 9324 11112 9376
rect 12164 9324 12216 9376
rect 15200 9324 15252 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 19432 9324 19484 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 9772 9120 9824 9172
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 15844 9120 15896 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 15200 9052 15252 9104
rect 9772 8984 9824 9036
rect 11612 8984 11664 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 9864 8916 9916 8968
rect 9312 8848 9364 8900
rect 10692 8916 10744 8968
rect 14004 8984 14056 9036
rect 14372 8916 14424 8968
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 18420 8984 18472 9036
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 18972 8916 19024 8968
rect 19331 9027 19383 9036
rect 19331 8993 19340 9027
rect 19340 8993 19374 9027
rect 19374 8993 19383 9027
rect 19331 8984 19383 8993
rect 17960 8848 18012 8900
rect 15108 8780 15160 8832
rect 15200 8780 15252 8832
rect 18788 8780 18840 8832
rect 19248 8780 19300 8832
rect 20444 8823 20496 8832
rect 20444 8789 20453 8823
rect 20453 8789 20487 8823
rect 20487 8789 20496 8823
rect 20444 8780 20496 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 5080 8576 5132 8628
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 14004 8508 14056 8560
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 10140 8372 10192 8424
rect 15016 8372 15068 8424
rect 18880 8576 18932 8628
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 16028 8372 16080 8424
rect 16764 8372 16816 8424
rect 18972 8415 19024 8424
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 8208 8236 8260 8288
rect 9312 8304 9364 8356
rect 10876 8304 10928 8356
rect 15200 8304 15252 8356
rect 15660 8347 15712 8356
rect 15660 8313 15669 8347
rect 15669 8313 15703 8347
rect 15703 8313 15712 8347
rect 15660 8304 15712 8313
rect 16120 8304 16172 8356
rect 16948 8304 17000 8356
rect 20444 8372 20496 8424
rect 10968 8236 11020 8288
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 14096 8236 14148 8288
rect 17224 8236 17276 8288
rect 19156 8236 19208 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 8208 8032 8260 8084
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 9772 8032 9824 8084
rect 11060 8032 11112 8084
rect 13268 8032 13320 8084
rect 8392 7964 8444 8016
rect 16120 8032 16172 8084
rect 16856 8032 16908 8084
rect 14004 7964 14056 8016
rect 9036 7896 9088 7948
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 11612 7896 11664 7948
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 14096 7896 14148 7948
rect 15844 7964 15896 8016
rect 17132 7964 17184 8016
rect 17500 8007 17552 8016
rect 17500 7973 17509 8007
rect 17509 7973 17543 8007
rect 17543 7973 17552 8007
rect 17500 7964 17552 7973
rect 19984 7964 20036 8016
rect 15752 7896 15804 7948
rect 13176 7871 13228 7880
rect 10876 7760 10928 7812
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 14556 7760 14608 7812
rect 20076 7896 20128 7948
rect 18880 7828 18932 7880
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 10692 7692 10744 7744
rect 14188 7692 14240 7744
rect 16396 7692 16448 7744
rect 18696 7692 18748 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 14556 7488 14608 7540
rect 11704 7420 11756 7472
rect 10600 7352 10652 7404
rect 10968 7284 11020 7336
rect 12072 7352 12124 7404
rect 16580 7488 16632 7540
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 20076 7352 20128 7404
rect 13544 7284 13596 7336
rect 16304 7284 16356 7336
rect 1216 7216 1268 7268
rect 12900 7216 12952 7268
rect 15292 7216 15344 7268
rect 16028 7216 16080 7268
rect 16396 7216 16448 7268
rect 18512 7216 18564 7268
rect 10324 7148 10376 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 13176 7148 13228 7200
rect 15936 7148 15988 7200
rect 16304 7148 16356 7200
rect 17960 7148 18012 7200
rect 19432 7148 19484 7200
rect 19616 7191 19668 7200
rect 19616 7157 19625 7191
rect 19625 7157 19659 7191
rect 19659 7157 19668 7191
rect 19616 7148 19668 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 11704 6944 11756 6996
rect 14096 6944 14148 6996
rect 15292 6987 15344 6996
rect 15292 6953 15301 6987
rect 15301 6953 15335 6987
rect 15335 6953 15344 6987
rect 15292 6944 15344 6953
rect 17408 6944 17460 6996
rect 19340 6987 19392 6996
rect 19340 6953 19349 6987
rect 19349 6953 19383 6987
rect 19383 6953 19392 6987
rect 19340 6944 19392 6953
rect 19800 6944 19852 6996
rect 19984 6944 20036 6996
rect 4712 6876 4764 6928
rect 15752 6876 15804 6928
rect 16580 6919 16632 6928
rect 16580 6885 16614 6919
rect 16614 6885 16632 6919
rect 16580 6876 16632 6885
rect 16948 6876 17000 6928
rect 19064 6876 19116 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10968 6851 11020 6860
rect 10968 6817 11002 6851
rect 11002 6817 11020 6851
rect 13820 6851 13872 6860
rect 10968 6808 11020 6817
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16304 6808 16356 6817
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10692 6783 10744 6792
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 9772 6672 9824 6724
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 15292 6740 15344 6792
rect 16028 6740 16080 6792
rect 12072 6715 12124 6724
rect 12072 6681 12081 6715
rect 12081 6681 12115 6715
rect 12115 6681 12124 6715
rect 12072 6672 12124 6681
rect 18788 6808 18840 6860
rect 19800 6808 19852 6860
rect 19984 6851 20036 6860
rect 19984 6817 19993 6851
rect 19993 6817 20027 6851
rect 20027 6817 20036 6851
rect 19984 6808 20036 6817
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 19432 6740 19484 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 19708 6672 19760 6724
rect 17500 6604 17552 6656
rect 19248 6604 19300 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 7564 6400 7616 6452
rect 9772 6400 9824 6452
rect 10968 6400 11020 6452
rect 11796 6400 11848 6452
rect 13820 6400 13872 6452
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 13360 6264 13412 6316
rect 14188 6264 14240 6316
rect 16304 6400 16356 6452
rect 17960 6400 18012 6452
rect 17316 6332 17368 6384
rect 17408 6307 17460 6316
rect 9772 6239 9824 6248
rect 9772 6205 9806 6239
rect 9806 6205 9824 6239
rect 8760 6128 8812 6180
rect 9772 6196 9824 6205
rect 12440 6196 12492 6248
rect 10692 6128 10744 6180
rect 12900 6128 12952 6180
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 19156 6400 19208 6452
rect 19524 6400 19576 6452
rect 19708 6400 19760 6452
rect 19340 6196 19392 6248
rect 20536 6239 20588 6248
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 18880 6128 18932 6180
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 11060 6060 11112 6112
rect 11612 6103 11664 6112
rect 11612 6069 11621 6103
rect 11621 6069 11655 6103
rect 11655 6069 11664 6103
rect 11612 6060 11664 6069
rect 12348 6060 12400 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 17132 6060 17184 6112
rect 19156 6060 19208 6112
rect 20168 6103 20220 6112
rect 20168 6069 20177 6103
rect 20177 6069 20211 6103
rect 20211 6069 20220 6103
rect 20168 6060 20220 6069
rect 20720 6103 20772 6112
rect 20720 6069 20729 6103
rect 20729 6069 20763 6103
rect 20763 6069 20772 6103
rect 20720 6060 20772 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 7196 5856 7248 5908
rect 10048 5856 10100 5908
rect 11152 5856 11204 5908
rect 7472 5720 7524 5772
rect 8208 5720 8260 5772
rect 6828 5652 6880 5704
rect 8760 5627 8812 5636
rect 8760 5593 8769 5627
rect 8769 5593 8803 5627
rect 8803 5593 8812 5627
rect 8760 5584 8812 5593
rect 10508 5788 10560 5840
rect 16764 5899 16816 5908
rect 16764 5865 16773 5899
rect 16773 5865 16807 5899
rect 16807 5865 16816 5899
rect 16764 5856 16816 5865
rect 17500 5856 17552 5908
rect 18512 5856 18564 5908
rect 19156 5856 19208 5908
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 11152 5720 11204 5772
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 13360 5763 13412 5772
rect 13360 5729 13394 5763
rect 13394 5729 13412 5763
rect 13360 5720 13412 5729
rect 15568 5788 15620 5840
rect 14096 5720 14148 5772
rect 10784 5584 10836 5636
rect 7104 5559 7156 5568
rect 7104 5525 7113 5559
rect 7113 5525 7147 5559
rect 7147 5525 7156 5559
rect 7104 5516 7156 5525
rect 10048 5516 10100 5568
rect 16488 5720 16540 5772
rect 15292 5627 15344 5636
rect 15292 5593 15301 5627
rect 15301 5593 15335 5627
rect 15335 5593 15344 5627
rect 15292 5584 15344 5593
rect 16120 5652 16172 5704
rect 16856 5720 16908 5772
rect 19248 5720 19300 5772
rect 19524 5720 19576 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 17316 5652 17368 5704
rect 17684 5652 17736 5704
rect 18788 5652 18840 5704
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 19984 5584 20036 5636
rect 11612 5516 11664 5568
rect 16304 5559 16356 5568
rect 16304 5525 16313 5559
rect 16313 5525 16347 5559
rect 16347 5525 16356 5559
rect 16304 5516 16356 5525
rect 19432 5516 19484 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 10140 5312 10192 5364
rect 10784 5312 10836 5364
rect 13912 5312 13964 5364
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 18604 5312 18656 5364
rect 19616 5355 19668 5364
rect 19616 5321 19625 5355
rect 19625 5321 19659 5355
rect 19659 5321 19668 5355
rect 19616 5312 19668 5321
rect 16028 5244 16080 5296
rect 8760 5176 8812 5228
rect 11152 5176 11204 5228
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 14188 5176 14240 5228
rect 16304 5176 16356 5228
rect 19156 5244 19208 5296
rect 17776 5176 17828 5228
rect 18788 5176 18840 5228
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7104 5151 7156 5160
rect 7104 5117 7138 5151
rect 7138 5117 7156 5151
rect 7104 5108 7156 5117
rect 9680 5108 9732 5160
rect 10048 5108 10100 5160
rect 14280 5108 14332 5160
rect 16580 5108 16632 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 19248 5108 19300 5160
rect 20628 5151 20680 5160
rect 20628 5117 20637 5151
rect 20637 5117 20671 5151
rect 20671 5117 20680 5151
rect 20628 5108 20680 5117
rect 11612 5040 11664 5092
rect 16396 5040 16448 5092
rect 17960 5040 18012 5092
rect 19708 5040 19760 5092
rect 8300 4972 8352 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 14188 4972 14240 5024
rect 16764 4972 16816 5024
rect 19892 4972 19944 5024
rect 20996 4972 21048 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 7288 4768 7340 4820
rect 9864 4768 9916 4820
rect 10876 4768 10928 4820
rect 14280 4768 14332 4820
rect 19340 4768 19392 4820
rect 7012 4700 7064 4752
rect 9128 4700 9180 4752
rect 16396 4700 16448 4752
rect 16856 4700 16908 4752
rect 20168 4700 20220 4752
rect 5172 4632 5224 4684
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 7104 4496 7156 4548
rect 5448 4428 5500 4480
rect 9036 4564 9088 4616
rect 9588 4496 9640 4548
rect 10968 4496 11020 4548
rect 14188 4632 14240 4684
rect 11612 4564 11664 4616
rect 16120 4632 16172 4684
rect 16212 4632 16264 4684
rect 18604 4632 18656 4684
rect 14556 4564 14608 4616
rect 13820 4471 13872 4480
rect 13820 4437 13829 4471
rect 13829 4437 13863 4471
rect 13863 4437 13872 4471
rect 13820 4428 13872 4437
rect 17684 4428 17736 4480
rect 17776 4428 17828 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 9036 4224 9088 4276
rect 9404 4088 9456 4140
rect 10876 4131 10928 4140
rect 6828 4020 6880 4072
rect 8668 4020 8720 4072
rect 10416 4020 10468 4072
rect 8576 3952 8628 4004
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 12348 4088 12400 4140
rect 12900 4088 12952 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13176 4088 13228 4140
rect 13820 4020 13872 4072
rect 14280 4088 14332 4140
rect 19340 4224 19392 4276
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 19616 4156 19668 4208
rect 19340 4088 19392 4140
rect 20904 4088 20956 4140
rect 22468 4088 22520 4140
rect 15200 4063 15252 4072
rect 15200 4029 15209 4063
rect 15209 4029 15243 4063
rect 15243 4029 15252 4063
rect 15200 4020 15252 4029
rect 17776 4020 17828 4072
rect 18604 4020 18656 4072
rect 18788 4020 18840 4072
rect 19432 4020 19484 4072
rect 20352 4020 20404 4072
rect 13728 3952 13780 4004
rect 18420 3952 18472 4004
rect 9680 3884 9732 3936
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 11704 3884 11756 3936
rect 12624 3884 12676 3936
rect 12716 3884 12768 3936
rect 14004 3884 14056 3936
rect 14464 3927 14516 3936
rect 14464 3893 14473 3927
rect 14473 3893 14507 3927
rect 14507 3893 14516 3927
rect 14464 3884 14516 3893
rect 15108 3884 15160 3936
rect 15200 3884 15252 3936
rect 16212 3884 16264 3936
rect 16488 3884 16540 3936
rect 17500 3927 17552 3936
rect 17500 3893 17509 3927
rect 17509 3893 17543 3927
rect 17543 3893 17552 3927
rect 17500 3884 17552 3893
rect 18052 3884 18104 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2320 3680 2372 3732
rect 8300 3680 8352 3732
rect 8576 3723 8628 3732
rect 8576 3689 8585 3723
rect 8585 3689 8619 3723
rect 8619 3689 8628 3723
rect 8576 3680 8628 3689
rect 2872 3612 2924 3664
rect 5172 3612 5224 3664
rect 12256 3680 12308 3732
rect 3424 3544 3476 3596
rect 5448 3544 5500 3596
rect 3976 3476 4028 3528
rect 13084 3680 13136 3732
rect 13728 3680 13780 3732
rect 18236 3680 18288 3732
rect 18052 3612 18104 3664
rect 6828 3544 6880 3596
rect 8208 3544 8260 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 11428 3544 11480 3596
rect 11980 3544 12032 3596
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 14280 3544 14332 3596
rect 15200 3544 15252 3596
rect 16488 3544 16540 3596
rect 12992 3476 13044 3528
rect 16580 3476 16632 3528
rect 18052 3476 18104 3528
rect 18880 3612 18932 3664
rect 18696 3587 18748 3596
rect 18696 3553 18705 3587
rect 18705 3553 18739 3587
rect 18739 3553 18748 3587
rect 18696 3544 18748 3553
rect 18880 3519 18932 3528
rect 5632 3340 5684 3392
rect 10600 3340 10652 3392
rect 10784 3340 10836 3392
rect 11152 3340 11204 3392
rect 13084 3340 13136 3392
rect 14556 3408 14608 3460
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 20076 3680 20128 3732
rect 19708 3612 19760 3664
rect 20720 3612 20772 3664
rect 20628 3544 20680 3596
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 20536 3476 20588 3528
rect 15936 3340 15988 3392
rect 18512 3340 18564 3392
rect 18696 3340 18748 3392
rect 18972 3340 19024 3392
rect 20536 3340 20588 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 6092 3136 6144 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 8392 3068 8444 3120
rect 10876 3136 10928 3188
rect 12716 3136 12768 3188
rect 14280 3179 14332 3188
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 1768 2932 1820 2984
rect 10600 3068 10652 3120
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 15108 3179 15160 3188
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 16120 3136 16172 3188
rect 17960 3136 18012 3188
rect 20168 3136 20220 3188
rect 15016 3068 15068 3120
rect 16028 3068 16080 3120
rect 8576 3000 8628 3052
rect 11612 3000 11664 3052
rect 11980 3043 12032 3052
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9680 2932 9732 2984
rect 10784 2932 10836 2984
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 12992 2932 13044 2984
rect 13636 2932 13688 2984
rect 15936 3000 15988 3052
rect 16488 3000 16540 3052
rect 15660 2932 15712 2984
rect 8300 2864 8352 2916
rect 13728 2864 13780 2916
rect 17040 2932 17092 2984
rect 17868 3000 17920 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 19340 3000 19392 3052
rect 19524 3000 19576 3052
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 17500 2932 17552 2984
rect 20444 2932 20496 2984
rect 11060 2796 11112 2848
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 13084 2796 13136 2848
rect 16396 2864 16448 2916
rect 17684 2864 17736 2916
rect 19248 2864 19300 2916
rect 21364 2864 21416 2916
rect 15476 2839 15528 2848
rect 15476 2805 15485 2839
rect 15485 2805 15519 2839
rect 15519 2805 15528 2839
rect 15476 2796 15528 2805
rect 16580 2839 16632 2848
rect 16580 2805 16589 2839
rect 16589 2805 16623 2839
rect 16623 2805 16632 2839
rect 16580 2796 16632 2805
rect 17040 2796 17092 2848
rect 18972 2796 19024 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 8944 2592 8996 2644
rect 10692 2592 10744 2644
rect 12440 2592 12492 2644
rect 15476 2592 15528 2644
rect 16672 2592 16724 2644
rect 17776 2592 17828 2644
rect 19248 2592 19300 2644
rect 7748 2524 7800 2576
rect 10968 2524 11020 2576
rect 15384 2524 15436 2576
rect 7196 2456 7248 2508
rect 11888 2456 11940 2508
rect 14372 2456 14424 2508
rect 16948 2499 17000 2508
rect 7564 2388 7616 2440
rect 8208 2388 8260 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 8852 2320 8904 2372
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 16948 2465 16957 2499
rect 16957 2465 16991 2499
rect 16991 2465 17000 2499
rect 16948 2456 17000 2465
rect 17224 2456 17276 2508
rect 17592 2456 17644 2508
rect 18236 2456 18288 2508
rect 18696 2456 18748 2508
rect 18880 2499 18932 2508
rect 18880 2465 18889 2499
rect 18889 2465 18923 2499
rect 18923 2465 18932 2499
rect 18880 2456 18932 2465
rect 19064 2456 19116 2508
rect 20260 2456 20312 2508
rect 14464 2320 14516 2372
rect 14832 2320 14884 2372
rect 17500 2320 17552 2372
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12624 2252 12676 2304
rect 16488 2252 16540 2304
rect 17960 2252 18012 2304
rect 21088 2388 21140 2440
rect 20812 2320 20864 2372
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 9956 1776 10008 1828
rect 15568 1776 15620 1828
rect 204 824 256 876
rect 8668 824 8720 876
rect 6644 552 6696 604
rect 7012 552 7064 604
<< metal2 >>
rect 5722 22320 5778 22800
rect 17130 22320 17186 22800
rect 18878 22536 18934 22545
rect 18878 22471 18934 22480
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 5736 19310 5764 22320
rect 17144 22250 17172 22320
rect 16684 22222 17172 22250
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15948 18902 15976 19246
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4066 11520 4122 11529
rect 4066 11455 4122 11464
rect 4080 11082 4108 11455
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 664 10464 716 10470
rect 664 10406 716 10412
rect 204 876 256 882
rect 204 818 256 824
rect 216 480 244 818
rect 676 480 704 10406
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 1216 7268 1268 7274
rect 1216 7210 1268 7216
rect 1228 480 1256 7210
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 480 1808 2926
rect 2332 480 2360 3674
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2884 480 2912 3606
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3436 480 3464 3538
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 480 4016 3470
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 1986 4752 6870
rect 4540 1958 4752 1986
rect 4540 480 4568 1958
rect 5092 480 5120 8570
rect 7576 6458 7604 18158
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8220 8090 8248 8230
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7208 5914 7236 6054
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5166 6868 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5166 7144 5510
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 3670 5212 4626
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5460 3602 5488 4422
rect 6840 4078 6868 5102
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6840 3602 6868 4014
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5644 480 5672 3334
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6104 480 6132 3130
rect 6840 3058 6868 3538
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 7024 610 7052 4694
rect 7116 4554 7144 5102
rect 7300 4826 7328 6054
rect 7484 5778 7512 6258
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5370 8248 5714
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7564 4616 7616 4622
rect 7562 4584 7564 4593
rect 7616 4584 7618 4593
rect 7104 4548 7156 4554
rect 7562 4519 7618 4528
rect 7104 4490 7156 4496
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 6644 604 6696 610
rect 6644 546 6696 552
rect 7012 604 7064 610
rect 7012 546 7064 552
rect 6656 480 6684 546
rect 7208 480 7236 2450
rect 7576 2446 7604 4519
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8312 3738 8340 4966
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8220 3194 8248 3538
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7760 480 7788 2518
rect 8220 2446 8248 3130
rect 8404 3126 8432 7958
rect 8496 3194 8524 14418
rect 9678 12472 9734 12481
rect 9678 12407 9734 12416
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9600 10470 9628 11222
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9324 8362 9352 8842
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 8090 9352 8298
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5642 8800 6122
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8772 5234 8800 5578
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 9048 4622 9076 7890
rect 9692 6730 9720 12407
rect 9784 9178 9812 14894
rect 9968 12481 9996 18770
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 9954 12472 10010 12481
rect 9954 12407 10010 12416
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8090 9812 8978
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9784 6458 9812 6666
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9784 6254 9812 6394
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4758 9168 4966
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9586 4584 9642 4593
rect 9048 4282 9076 4558
rect 9586 4519 9588 4528
rect 9640 4519 9642 4528
rect 9588 4490 9640 4496
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8588 3738 8616 3946
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8588 3058 8616 3674
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8312 480 8340 2858
rect 8680 882 8708 4014
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 2990 8892 3470
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8956 2650 8984 2926
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8668 876 8720 882
rect 8668 818 8720 824
rect 8864 480 8892 2314
rect 9416 480 9444 4082
rect 9692 3942 9720 5102
rect 9876 4826 9904 8910
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10152 7750 10180 8366
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 5914 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 5166 10088 5510
rect 10152 5370 10180 6734
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 10244 3942 10272 13806
rect 10888 12442 10916 17682
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11164 13938 11192 14282
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10692 8968 10744 8974
rect 10796 8956 10824 11086
rect 11072 9738 11100 12378
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11072 9710 11192 9738
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10744 8928 10824 8956
rect 10692 8910 10744 8916
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10336 7206 10364 7890
rect 10704 7750 10732 8910
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10888 7818 10916 8298
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10600 7404 10652 7410
rect 10704 7392 10732 7686
rect 10652 7364 10732 7392
rect 10600 7346 10652 7352
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 5778 10364 7142
rect 10704 6798 10732 7364
rect 10980 7342 11008 8230
rect 11072 8090 11100 9318
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6186 10732 6734
rect 10980 6458 11008 6802
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10414 5264 10470 5273
rect 10414 5199 10470 5208
rect 10428 4078 10456 5199
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9692 3602 9720 3878
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9692 2990 9720 3538
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 9968 480 9996 1770
rect 10520 480 10548 5782
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5370 10824 5578
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10888 4826 10916 5646
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 3126 10640 3334
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10704 2650 10732 3878
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 2990 10824 3334
rect 10888 3194 10916 4082
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10796 2446 10824 2926
rect 10980 2582 11008 4490
rect 11072 2854 11100 6054
rect 11164 5914 11192 9710
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11624 9042 11652 9522
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8634 11652 8978
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11624 6118 11652 7890
rect 11716 7478 11744 18770
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14476 17202 14504 17682
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 11900 9654 11928 15506
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11900 8498 11928 9386
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11716 7002 11744 7142
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11808 6458 11836 7142
rect 11992 6610 12020 10474
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 6730 12112 7346
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11900 6582 12020 6610
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11164 5234 11192 5714
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11624 5098 11652 5510
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11624 4622 11652 5034
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11440 3482 11468 3538
rect 11440 3454 11652 3482
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11164 1850 11192 3334
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11624 3058 11652 3454
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11716 2990 11744 3878
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11900 2514 11928 6582
rect 12176 4706 12204 9318
rect 12452 9042 12480 9454
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12348 6112 12400 6118
rect 12452 6100 12480 6190
rect 12400 6072 12480 6100
rect 12348 6054 12400 6060
rect 12084 4678 12204 4706
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11992 3058 12020 3538
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11072 1822 11192 1850
rect 11072 480 11100 1822
rect 11624 480 11652 2246
rect 12084 480 12112 4678
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12360 3754 12388 4082
rect 12636 3942 12664 13262
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 11694 13400 12174
rect 13464 11762 13492 12242
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13188 11354 13216 11630
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9586 13124 10066
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12912 7274 12940 7890
rect 13188 7886 13216 11154
rect 13280 8090 13308 11494
rect 13464 11082 13492 11698
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13832 10266 13860 15506
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13832 9450 13860 9998
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13832 9178 13860 9386
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 13188 7206 13216 7822
rect 13556 7342 13584 7822
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13924 6882 13952 12854
rect 14016 12424 14044 17070
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14016 12396 14228 12424
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14016 8566 14044 8978
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14016 8022 14044 8230
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 14108 7954 14136 8230
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14200 7834 14228 12396
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 11694 15332 12174
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15304 11014 15332 11630
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15304 10198 15332 10950
rect 15396 10810 15424 15982
rect 15672 12986 15700 18770
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15580 11354 15608 12582
rect 15764 11898 15792 12786
rect 16132 12374 16160 13806
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15764 11694 15792 11834
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15856 11626 15884 12038
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15856 11150 15884 11562
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15764 10266 15792 10474
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14108 7806 14228 7834
rect 14108 7002 14136 7806
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 13820 6860 13872 6866
rect 13924 6854 14044 6882
rect 13820 6802 13872 6808
rect 13832 6458 13860 6802
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12912 4146 12940 6122
rect 13372 5778 13400 6258
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13556 5234 13584 6054
rect 13924 5370 13952 6734
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12268 3738 12388 3754
rect 12256 3732 12388 3738
rect 12308 3726 12388 3732
rect 12256 3674 12308 3680
rect 12728 3194 12756 3878
rect 13096 3738 13124 4082
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 13004 2990 13032 3470
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 13096 2854 13124 3334
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12452 2650 12480 2790
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12636 480 12664 2246
rect 13188 480 13216 4082
rect 13832 4078 13860 4422
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13740 3738 13768 3946
rect 14016 3942 14044 6854
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 5778 14136 6734
rect 14200 6322 14228 7686
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14200 5234 14228 6258
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4690 14228 4966
rect 14292 4826 14320 5102
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13648 2446 13676 2926
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13740 480 13768 2858
rect 14108 2020 14136 3975
rect 14292 3602 14320 4082
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3194 14320 3538
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14384 2514 14412 8910
rect 14568 8634 14596 10066
rect 15212 9382 15240 10066
rect 15304 10062 15332 10134
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15304 9518 15332 9998
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15212 9110 15240 9318
rect 15856 9178 15884 10406
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15752 8968 15804 8974
rect 15948 8956 15976 11154
rect 15804 8928 15976 8956
rect 15752 8910 15804 8916
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 15120 8498 15148 8774
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 7546 14596 7754
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14476 2378 14504 3878
rect 14568 3466 14596 4558
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 15028 3126 15056 8366
rect 15212 8362 15240 8774
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15304 7002 15332 7210
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 5642 15332 6734
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15212 3942 15240 4014
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15120 3194 15148 3878
rect 15212 3602 15240 3878
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15488 2650 15516 2790
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 14108 1992 14320 2020
rect 14292 480 14320 1992
rect 14844 480 14872 2314
rect 15396 480 15424 2518
rect 15580 1834 15608 5782
rect 15672 2990 15700 8298
rect 15856 8022 15884 8928
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 16040 7970 16068 8366
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16132 8090 16160 8298
rect 16316 8106 16344 11154
rect 16408 9178 16436 16594
rect 16684 13870 16712 22222
rect 18694 21584 18750 21593
rect 18694 21519 18750 21528
rect 17866 21176 17922 21185
rect 17866 21111 17922 21120
rect 17880 19174 17908 21111
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17972 18902 18000 19246
rect 18708 19174 18736 21519
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17866 18320 17922 18329
rect 17866 18255 17922 18264
rect 17880 17882 17908 18255
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16592 10810 16620 12650
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11898 16804 12242
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16776 10674 16804 11834
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16500 9926 16528 10610
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9518 16528 9862
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16120 8084 16172 8090
rect 16316 8078 16436 8106
rect 16120 8026 16172 8032
rect 15752 7948 15804 7954
rect 16040 7942 16344 7970
rect 15752 7890 15804 7896
rect 15764 6934 15792 7890
rect 16316 7342 16344 7942
rect 16408 7750 16436 8078
rect 16684 7886 16712 10474
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 8430 16804 9318
rect 16960 9058 16988 10406
rect 16960 9030 17080 9058
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16776 7886 16804 8366
rect 16868 8090 16896 8910
rect 16960 8362 16988 8910
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15948 5370 15976 7142
rect 16040 6798 16068 7210
rect 16316 7206 16344 7278
rect 16408 7274 16436 7686
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 6866 16344 7142
rect 16592 6934 16620 7482
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6118 16068 6734
rect 16316 6458 16344 6802
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16040 5302 16068 6054
rect 16120 5704 16172 5710
rect 16316 5658 16344 6394
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16120 5646 16172 5652
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 16132 4690 16160 5646
rect 16224 5630 16344 5658
rect 16224 4690 16252 5630
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16316 5234 16344 5510
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16408 5098 16436 6054
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 5522 16528 5714
rect 16500 5494 16620 5522
rect 16592 5166 16620 5494
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 3058 15976 3334
rect 16132 3194 16160 4626
rect 16224 3942 16252 4626
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15568 1828 15620 1834
rect 15568 1770 15620 1776
rect 16040 1578 16068 3062
rect 16408 2922 16436 4694
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 3602 16528 3878
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16500 3058 16528 3538
rect 16592 3534 16620 5102
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 15948 1550 16068 1578
rect 15948 480 15976 1550
rect 16408 1057 16436 2858
rect 16500 2446 16528 2994
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16394 1048 16450 1057
rect 16394 983 16450 992
rect 16500 480 16528 2246
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6090 0 6146 480
rect 6642 0 6698 480
rect 7194 0 7250 480
rect 7746 0 7802 480
rect 8298 0 8354 480
rect 8850 0 8906 480
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12622 0 12678 480
rect 13174 0 13230 480
rect 13726 0 13782 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 16592 241 16620 2790
rect 16684 2650 16712 7822
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16776 5030 16804 5850
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16868 4758 16896 5714
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16960 2514 16988 6870
rect 17052 2990 17080 9030
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17144 6118 17172 7958
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17144 3777 17172 6054
rect 17130 3768 17186 3777
rect 17130 3703 17186 3712
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 17052 480 17080 2790
rect 17236 2514 17264 8230
rect 17328 6390 17356 13942
rect 17972 12986 18000 18702
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 8022 17540 12718
rect 18510 12472 18566 12481
rect 18510 12407 18566 12416
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17604 11762 17632 12242
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 18524 11694 18552 12407
rect 18616 12374 18644 12786
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10674 18000 10950
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17972 10198 18000 10610
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9586 17632 10066
rect 18064 10010 18092 10406
rect 18432 10266 18460 10406
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 17972 9982 18092 10010
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17972 8906 18000 9982
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 9042 18460 9522
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17866 7440 17922 7449
rect 17866 7375 17922 7384
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17328 5710 17356 6326
rect 17420 6322 17448 6938
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17512 5914 17540 6598
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17696 4486 17724 5646
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4486 17816 5170
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17512 2990 17540 3878
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17696 2922 17724 4422
rect 17788 4078 17816 4422
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17880 3058 17908 7375
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17972 6798 18000 7142
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17972 6458 18000 6734
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18524 5914 18552 7210
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18616 5370 18644 12174
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18708 11150 18736 11630
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18800 8838 18828 13670
rect 18892 12730 18920 22471
rect 19798 22128 19854 22137
rect 19798 22063 19854 22072
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19628 16130 19656 18770
rect 19812 17490 19840 22063
rect 20626 20768 20682 20777
rect 20626 20703 20682 20712
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19904 18902 19932 19858
rect 20180 19514 20208 20159
rect 20640 20058 20668 20703
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20166 19408 20222 19417
rect 20166 19343 20222 19352
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19996 18630 20024 19246
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 20180 18426 20208 19343
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20442 18864 20498 18873
rect 20442 18799 20498 18808
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20456 17882 20484 18799
rect 20548 18222 20576 18906
rect 20732 18426 20760 19751
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20718 18048 20774 18057
rect 20718 17983 20774 17992
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20166 17504 20222 17513
rect 19812 17462 19932 17490
rect 19536 16102 19656 16130
rect 19246 14376 19302 14385
rect 19246 14311 19302 14320
rect 19260 14074 19288 14311
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19246 13832 19302 13841
rect 19246 13767 19302 13776
rect 19260 13530 19288 13767
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19246 13016 19302 13025
rect 19246 12951 19248 12960
rect 19300 12951 19302 12960
rect 19248 12922 19300 12928
rect 18892 12702 19196 12730
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11694 18920 12038
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18892 8634 18920 11222
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 18984 9518 19012 9930
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18892 7886 18920 8570
rect 18984 8430 19012 8910
rect 19076 8498 19104 9862
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 19168 8378 19196 12702
rect 19352 12374 19380 13330
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19246 11656 19302 11665
rect 19536 11626 19564 16102
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19628 15502 19656 15982
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 13462 19748 14418
rect 19904 13870 19932 17462
rect 20166 17439 20222 17448
rect 20180 17338 20208 17439
rect 20732 17338 20760 17983
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20718 17096 20774 17105
rect 19996 16114 20024 17070
rect 20548 16726 20576 17070
rect 20718 17031 20774 17040
rect 20536 16720 20588 16726
rect 20536 16662 20588 16668
rect 20442 16552 20498 16561
rect 20442 16487 20498 16496
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 20166 15736 20222 15745
rect 20456 15706 20484 16487
rect 20732 16250 20760 17031
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20718 16144 20774 16153
rect 20718 16079 20774 16088
rect 20166 15671 20222 15680
rect 20444 15700 20496 15706
rect 20180 15162 20208 15671
rect 20444 15642 20496 15648
rect 20442 15192 20498 15201
rect 20168 15156 20220 15162
rect 20732 15162 20760 16079
rect 20442 15127 20498 15136
rect 20720 15156 20772 15162
rect 20168 15098 20220 15104
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19996 14414 20024 14894
rect 20074 14784 20130 14793
rect 20074 14719 20130 14728
rect 20088 14618 20116 14719
rect 20456 14618 20484 15127
rect 20720 15098 20772 15104
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19708 13456 19760 13462
rect 19708 13398 19760 13404
rect 19812 12850 19840 13738
rect 20442 13424 20498 13433
rect 20442 13359 20498 13368
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 19246 11591 19302 11600
rect 19524 11620 19576 11626
rect 19260 9518 19288 11591
rect 19524 11562 19576 11568
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19352 10606 19380 11290
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19706 10160 19762 10169
rect 19706 10095 19708 10104
rect 19760 10095 19762 10104
rect 19708 10066 19760 10072
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9058 19472 9318
rect 19343 9042 19472 9058
rect 19331 9036 19472 9042
rect 19383 9030 19472 9036
rect 19331 8978 19383 8984
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8498 19288 8774
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19168 8350 19288 8378
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19062 7984 19118 7993
rect 19062 7919 19118 7928
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 3194 18000 5034
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18616 4078 18644 4626
rect 18604 4072 18656 4078
rect 18418 4040 18474 4049
rect 18604 4014 18656 4020
rect 18418 3975 18420 3984
rect 18472 3975 18474 3984
rect 18420 3946 18472 3952
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3670 18092 3878
rect 18234 3768 18290 3777
rect 18234 3703 18236 3712
rect 18288 3703 18290 3712
rect 18602 3768 18658 3777
rect 18602 3703 18658 3712
rect 18236 3674 18288 3680
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 18052 3528 18104 3534
rect 18050 3496 18052 3505
rect 18104 3496 18106 3505
rect 18050 3431 18106 3440
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18524 3058 18552 3334
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 17774 2952 17830 2961
rect 17684 2916 17736 2922
rect 17774 2887 17830 2896
rect 17684 2858 17736 2864
rect 17788 2650 17816 2887
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18616 2530 18644 3703
rect 18708 3602 18736 7686
rect 18970 7032 19026 7041
rect 18970 6967 19026 6976
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18800 5710 18828 6802
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18800 5234 18828 5646
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18248 2514 18644 2530
rect 18708 2514 18736 3334
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 18236 2508 18644 2514
rect 18288 2502 18644 2508
rect 18696 2508 18748 2514
rect 18236 2450 18288 2456
rect 18696 2450 18748 2456
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 17512 480 17540 2314
rect 17604 2009 17632 2450
rect 18800 2394 18828 4014
rect 18892 3670 18920 6122
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18892 2514 18920 3470
rect 18984 3398 19012 6967
rect 19076 6934 19104 7919
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19168 6458 19196 8230
rect 19260 6662 19288 8350
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19168 5914 19196 6054
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19260 5778 19288 6598
rect 19352 6254 19380 6938
rect 19444 6798 19472 7142
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19536 6458 19564 9862
rect 19812 9466 19840 12650
rect 20272 12306 20300 12650
rect 20456 12442 20484 13359
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20626 12064 20682 12073
rect 20626 11999 20682 12008
rect 20640 11762 20668 11999
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 19996 11286 20024 11494
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19996 10674 20024 11222
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 20272 10606 20300 11494
rect 20350 10704 20406 10713
rect 20350 10639 20406 10648
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19720 9438 19840 9466
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19340 6248 19392 6254
rect 19392 6196 19472 6202
rect 19340 6190 19472 6196
rect 19352 6174 19472 6190
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19444 5710 19472 6174
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19156 5296 19208 5302
rect 19156 5238 19208 5244
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4729 19104 5102
rect 19062 4720 19118 4729
rect 19062 4655 19118 4664
rect 19062 4312 19118 4321
rect 19062 4247 19118 4256
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18616 2366 18828 2394
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17590 2000 17646 2009
rect 17590 1935 17646 1944
rect 17972 1170 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18092 1170
rect 18064 480 18092 1142
rect 18616 480 18644 2366
rect 18984 649 19012 2790
rect 19076 2514 19104 4247
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 18970 640 19026 649
rect 18970 575 19026 584
rect 19168 480 19196 5238
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19260 3097 19288 5102
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19352 4282 19380 4762
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19352 4146 19380 4218
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19246 3088 19302 3097
rect 19352 3058 19380 4082
rect 19444 4078 19472 5510
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19536 3058 19564 5714
rect 19628 5370 19656 7142
rect 19720 6730 19748 9438
rect 19996 8022 20024 10134
rect 20364 10130 20392 10639
rect 20456 10470 20484 11494
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20534 11112 20590 11121
rect 20534 11047 20590 11056
rect 20548 10674 20576 11047
rect 20640 10674 20668 11154
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 10198 20484 10406
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20350 9752 20406 9761
rect 20350 9687 20406 9696
rect 20166 8800 20222 8809
rect 20166 8735 20222 8744
rect 19984 8016 20036 8022
rect 19984 7958 20036 7964
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19812 7002 19840 7346
rect 19996 7002 20024 7958
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 20088 7410 20116 7890
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 20180 6882 20208 8735
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 20088 6854 20208 6882
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19720 5250 19748 6394
rect 19812 5273 19840 6802
rect 19996 5642 20024 6802
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19628 5222 19748 5250
rect 19798 5264 19854 5273
rect 19628 4214 19656 5222
rect 19798 5199 19854 5208
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19720 4282 19748 5034
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19904 3890 19932 4966
rect 20088 4570 20116 6854
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20180 6118 20208 6734
rect 20272 6633 20300 7822
rect 20258 6624 20314 6633
rect 20258 6559 20314 6568
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20258 6080 20314 6089
rect 20180 4758 20208 6054
rect 20258 6015 20314 6024
rect 20272 5778 20300 6015
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20168 4752 20220 4758
rect 20168 4694 20220 4700
rect 20088 4542 20300 4570
rect 20076 3936 20128 3942
rect 19904 3862 20024 3890
rect 20076 3878 20128 3884
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 19246 3023 19302 3032
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19260 2650 19288 2858
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19720 480 19748 3606
rect 19996 2122 20024 3862
rect 20088 3738 20116 3878
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 3058 20116 3470
rect 20180 3194 20208 3878
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20272 2514 20300 4542
rect 20364 4078 20392 9687
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20456 8430 20484 8774
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20534 8392 20590 8401
rect 20456 7886 20484 8366
rect 20534 8327 20590 8336
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20548 6338 20576 8327
rect 20456 6310 20576 6338
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20456 2990 20484 6310
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20548 5137 20576 6190
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20626 5672 20682 5681
rect 20626 5607 20682 5616
rect 20640 5166 20668 5607
rect 20628 5160 20680 5166
rect 20534 5128 20590 5137
rect 20628 5102 20680 5108
rect 20534 5063 20590 5072
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 3534 20576 4422
rect 20732 3670 20760 6054
rect 20916 4146 20944 19110
rect 21916 11620 21968 11626
rect 21916 11562 21968 11568
rect 21086 9344 21142 9353
rect 21086 9279 21142 9288
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20548 2417 20576 3334
rect 20534 2408 20590 2417
rect 20534 2343 20590 2352
rect 19996 2094 20300 2122
rect 20272 480 20300 2094
rect 20640 1601 20668 3538
rect 20812 2372 20864 2378
rect 20812 2314 20864 2320
rect 20626 1592 20682 1601
rect 20626 1527 20682 1536
rect 20824 480 20852 2314
rect 21008 2009 21036 4966
rect 21100 2446 21128 9279
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 20994 2000 21050 2009
rect 20994 1935 21050 1944
rect 21376 480 21404 2858
rect 21928 480 21956 11562
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22480 480 22508 4082
rect 16578 232 16634 241
rect 16578 167 16634 176
rect 17038 0 17094 480
rect 17498 0 17554 480
rect 18050 0 18106 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19706 0 19762 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
<< via2 >>
rect 18878 22480 18934 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11464 4122 11520
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7562 4564 7564 4584
rect 7564 4564 7616 4584
rect 7616 4564 7618 4584
rect 7562 4528 7618 4564
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9678 12416 9734 12472
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 9954 12416 10010 12472
rect 9586 4548 9642 4584
rect 9586 4528 9588 4548
rect 9588 4528 9640 4548
rect 9640 4528 9642 4548
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 10414 5208 10470 5264
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14094 3984 14150 4040
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18694 21528 18750 21584
rect 17866 21120 17922 21176
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17866 18264 17922 18320
rect 16394 992 16450 1048
rect 17130 3712 17186 3768
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18510 12416 18566 12472
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 17866 7384 17922 7440
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 19798 22072 19854 22128
rect 20626 20712 20682 20768
rect 20166 20168 20222 20224
rect 20718 19760 20774 19816
rect 20166 19352 20222 19408
rect 20442 18808 20498 18864
rect 20718 17992 20774 18048
rect 19246 14320 19302 14376
rect 19246 13776 19302 13832
rect 19246 12980 19302 13016
rect 19246 12960 19248 12980
rect 19248 12960 19300 12980
rect 19300 12960 19302 12980
rect 19246 11600 19302 11656
rect 20166 17448 20222 17504
rect 20718 17040 20774 17096
rect 20442 16496 20498 16552
rect 20166 15680 20222 15736
rect 20718 16088 20774 16144
rect 20442 15136 20498 15192
rect 20074 14728 20130 14784
rect 20442 13368 20498 13424
rect 19706 10124 19762 10160
rect 19706 10104 19708 10124
rect 19708 10104 19760 10124
rect 19760 10104 19762 10124
rect 19062 7928 19118 7984
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18418 4004 18474 4040
rect 18418 3984 18420 4004
rect 18420 3984 18472 4004
rect 18472 3984 18474 4004
rect 18234 3732 18290 3768
rect 18234 3712 18236 3732
rect 18236 3712 18288 3732
rect 18288 3712 18290 3732
rect 18602 3712 18658 3768
rect 18050 3476 18052 3496
rect 18052 3476 18104 3496
rect 18104 3476 18106 3496
rect 18050 3440 18106 3476
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 17774 2896 17830 2952
rect 18970 6976 19026 7032
rect 20626 12008 20682 12064
rect 20350 10648 20406 10704
rect 19062 4664 19118 4720
rect 19062 4256 19118 4312
rect 17590 1944 17646 2000
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18970 584 19026 640
rect 19246 3032 19302 3088
rect 20534 11056 20590 11112
rect 20350 9696 20406 9752
rect 20166 8744 20222 8800
rect 19798 5208 19854 5264
rect 20258 6568 20314 6624
rect 20258 6024 20314 6080
rect 20534 8336 20590 8392
rect 20626 5616 20682 5672
rect 20534 5072 20590 5128
rect 21086 9288 21142 9344
rect 20534 2352 20590 2408
rect 20626 1536 20682 1592
rect 20994 1944 21050 2000
rect 16578 176 16634 232
<< metal3 >>
rect 18873 22538 18939 22541
rect 22320 22538 22800 22568
rect 18873 22536 22800 22538
rect 18873 22480 18878 22536
rect 18934 22480 22800 22536
rect 18873 22478 22800 22480
rect 18873 22475 18939 22478
rect 22320 22448 22800 22478
rect 19793 22130 19859 22133
rect 22320 22130 22800 22160
rect 19793 22128 22800 22130
rect 19793 22072 19798 22128
rect 19854 22072 22800 22128
rect 19793 22070 22800 22072
rect 19793 22067 19859 22070
rect 22320 22040 22800 22070
rect 18689 21586 18755 21589
rect 22320 21586 22800 21616
rect 18689 21584 22800 21586
rect 18689 21528 18694 21584
rect 18750 21528 22800 21584
rect 18689 21526 22800 21528
rect 18689 21523 18755 21526
rect 22320 21496 22800 21526
rect 17861 21178 17927 21181
rect 22320 21178 22800 21208
rect 17861 21176 22800 21178
rect 17861 21120 17866 21176
rect 17922 21120 22800 21176
rect 17861 21118 22800 21120
rect 17861 21115 17927 21118
rect 22320 21088 22800 21118
rect 20621 20770 20687 20773
rect 22320 20770 22800 20800
rect 20621 20768 22800 20770
rect 20621 20712 20626 20768
rect 20682 20712 22800 20768
rect 20621 20710 22800 20712
rect 20621 20707 20687 20710
rect 22320 20680 22800 20710
rect 20161 20226 20227 20229
rect 22320 20226 22800 20256
rect 20161 20224 22800 20226
rect 20161 20168 20166 20224
rect 20222 20168 22800 20224
rect 20161 20166 22800 20168
rect 20161 20163 20227 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 20713 19818 20779 19821
rect 22320 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 20161 19410 20227 19413
rect 22320 19410 22800 19440
rect 20161 19408 22800 19410
rect 20161 19352 20166 19408
rect 20222 19352 22800 19408
rect 20161 19350 22800 19352
rect 20161 19347 20227 19350
rect 22320 19320 22800 19350
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 20437 18866 20503 18869
rect 22320 18866 22800 18896
rect 20437 18864 22800 18866
rect 20437 18808 20442 18864
rect 20498 18808 22800 18864
rect 20437 18806 22800 18808
rect 20437 18803 20503 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 22320 18458 22800 18488
rect 18646 18398 22800 18458
rect 17861 18322 17927 18325
rect 18646 18322 18706 18398
rect 22320 18368 22800 18398
rect 17861 18320 18706 18322
rect 17861 18264 17866 18320
rect 17922 18264 18706 18320
rect 17861 18262 18706 18264
rect 17861 18259 17927 18262
rect 20713 18050 20779 18053
rect 22320 18050 22800 18080
rect 20713 18048 22800 18050
rect 20713 17992 20718 18048
rect 20774 17992 22800 18048
rect 20713 17990 22800 17992
rect 20713 17987 20779 17990
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 22320 17960 22800 17990
rect 14672 17919 14992 17920
rect 20161 17506 20227 17509
rect 22320 17506 22800 17536
rect 20161 17504 22800 17506
rect 20161 17448 20166 17504
rect 20222 17448 22800 17504
rect 20161 17446 22800 17448
rect 20161 17443 20227 17446
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 22320 17416 22800 17446
rect 18104 17375 18424 17376
rect 20713 17098 20779 17101
rect 22320 17098 22800 17128
rect 20713 17096 22800 17098
rect 20713 17040 20718 17096
rect 20774 17040 22800 17096
rect 20713 17038 22800 17040
rect 20713 17035 20779 17038
rect 22320 17008 22800 17038
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 20437 16554 20503 16557
rect 22320 16554 22800 16584
rect 20437 16552 22800 16554
rect 20437 16496 20442 16552
rect 20498 16496 22800 16552
rect 20437 16494 22800 16496
rect 20437 16491 20503 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 20713 16146 20779 16149
rect 22320 16146 22800 16176
rect 20713 16144 22800 16146
rect 20713 16088 20718 16144
rect 20774 16088 22800 16144
rect 20713 16086 22800 16088
rect 20713 16083 20779 16086
rect 22320 16056 22800 16086
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 20161 15738 20227 15741
rect 22320 15738 22800 15768
rect 20161 15736 22800 15738
rect 20161 15680 20166 15736
rect 20222 15680 22800 15736
rect 20161 15678 22800 15680
rect 20161 15675 20227 15678
rect 22320 15648 22800 15678
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 20437 15194 20503 15197
rect 22320 15194 22800 15224
rect 20437 15192 22800 15194
rect 20437 15136 20442 15192
rect 20498 15136 22800 15192
rect 20437 15134 22800 15136
rect 20437 15131 20503 15134
rect 22320 15104 22800 15134
rect 20069 14786 20135 14789
rect 22320 14786 22800 14816
rect 20069 14784 22800 14786
rect 20069 14728 20074 14784
rect 20130 14728 22800 14784
rect 20069 14726 22800 14728
rect 20069 14723 20135 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 22320 14696 22800 14726
rect 14672 14655 14992 14656
rect 19241 14378 19307 14381
rect 22320 14378 22800 14408
rect 19241 14376 22800 14378
rect 19241 14320 19246 14376
rect 19302 14320 22800 14376
rect 19241 14318 22800 14320
rect 19241 14315 19307 14318
rect 22320 14288 22800 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19241 13834 19307 13837
rect 22320 13834 22800 13864
rect 19241 13832 22800 13834
rect 19241 13776 19246 13832
rect 19302 13776 22800 13832
rect 19241 13774 22800 13776
rect 19241 13771 19307 13774
rect 22320 13744 22800 13774
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 20437 13426 20503 13429
rect 22320 13426 22800 13456
rect 20437 13424 22800 13426
rect 20437 13368 20442 13424
rect 20498 13368 22800 13424
rect 20437 13366 22800 13368
rect 20437 13363 20503 13366
rect 22320 13336 22800 13366
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 19241 13018 19307 13021
rect 22320 13018 22800 13048
rect 19241 13016 22800 13018
rect 19241 12960 19246 13016
rect 19302 12960 22800 13016
rect 19241 12958 22800 12960
rect 19241 12955 19307 12958
rect 22320 12928 22800 12958
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 9673 12474 9739 12477
rect 9949 12474 10015 12477
rect 9673 12472 10015 12474
rect 9673 12416 9678 12472
rect 9734 12416 9954 12472
rect 10010 12416 10015 12472
rect 9673 12414 10015 12416
rect 9673 12411 9739 12414
rect 9949 12411 10015 12414
rect 18505 12474 18571 12477
rect 22320 12474 22800 12504
rect 18505 12472 22800 12474
rect 18505 12416 18510 12472
rect 18566 12416 22800 12472
rect 18505 12414 22800 12416
rect 18505 12411 18571 12414
rect 22320 12384 22800 12414
rect 20621 12066 20687 12069
rect 22320 12066 22800 12096
rect 20621 12064 22800 12066
rect 20621 12008 20626 12064
rect 20682 12008 22800 12064
rect 20621 12006 22800 12008
rect 20621 12003 20687 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 22320 11976 22800 12006
rect 18104 11935 18424 11936
rect 19241 11658 19307 11661
rect 22320 11658 22800 11688
rect 19241 11656 22800 11658
rect 19241 11600 19246 11656
rect 19302 11600 22800 11656
rect 19241 11598 22800 11600
rect 19241 11595 19307 11598
rect 22320 11568 22800 11598
rect 0 11522 480 11552
rect 4061 11522 4127 11525
rect 0 11520 4127 11522
rect 0 11464 4066 11520
rect 4122 11464 4127 11520
rect 0 11462 4127 11464
rect 0 11432 480 11462
rect 4061 11459 4127 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 20529 11114 20595 11117
rect 22320 11114 22800 11144
rect 20529 11112 22800 11114
rect 20529 11056 20534 11112
rect 20590 11056 22800 11112
rect 20529 11054 22800 11056
rect 20529 11051 20595 11054
rect 22320 11024 22800 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 20345 10706 20411 10709
rect 22320 10706 22800 10736
rect 20345 10704 22800 10706
rect 20345 10648 20350 10704
rect 20406 10648 22800 10704
rect 20345 10646 22800 10648
rect 20345 10643 20411 10646
rect 22320 10616 22800 10646
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 19701 10162 19767 10165
rect 22320 10162 22800 10192
rect 19701 10160 22800 10162
rect 19701 10104 19706 10160
rect 19762 10104 22800 10160
rect 19701 10102 22800 10104
rect 19701 10099 19767 10102
rect 22320 10072 22800 10102
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 20345 9754 20411 9757
rect 22320 9754 22800 9784
rect 20345 9752 22800 9754
rect 20345 9696 20350 9752
rect 20406 9696 22800 9752
rect 20345 9694 22800 9696
rect 20345 9691 20411 9694
rect 22320 9664 22800 9694
rect 21081 9346 21147 9349
rect 22320 9346 22800 9376
rect 21081 9344 22800 9346
rect 21081 9288 21086 9344
rect 21142 9288 22800 9344
rect 21081 9286 22800 9288
rect 21081 9283 21147 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 22320 9256 22800 9286
rect 14672 9215 14992 9216
rect 20161 8802 20227 8805
rect 22320 8802 22800 8832
rect 20161 8800 22800 8802
rect 20161 8744 20166 8800
rect 20222 8744 22800 8800
rect 20161 8742 22800 8744
rect 20161 8739 20227 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22320 8712 22800 8742
rect 18104 8671 18424 8672
rect 20529 8394 20595 8397
rect 22320 8394 22800 8424
rect 20529 8392 22800 8394
rect 20529 8336 20534 8392
rect 20590 8336 22800 8392
rect 20529 8334 22800 8336
rect 20529 8331 20595 8334
rect 22320 8304 22800 8334
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 19057 7986 19123 7989
rect 22320 7986 22800 8016
rect 19057 7984 22800 7986
rect 19057 7928 19062 7984
rect 19118 7928 22800 7984
rect 19057 7926 22800 7928
rect 19057 7923 19123 7926
rect 22320 7896 22800 7926
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 17861 7442 17927 7445
rect 22320 7442 22800 7472
rect 17861 7440 22800 7442
rect 17861 7384 17866 7440
rect 17922 7384 22800 7440
rect 17861 7382 22800 7384
rect 17861 7379 17927 7382
rect 22320 7352 22800 7382
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 18965 7034 19031 7037
rect 22320 7034 22800 7064
rect 18965 7032 22800 7034
rect 18965 6976 18970 7032
rect 19026 6976 22800 7032
rect 18965 6974 22800 6976
rect 18965 6971 19031 6974
rect 22320 6944 22800 6974
rect 20253 6626 20319 6629
rect 22320 6626 22800 6656
rect 20253 6624 22800 6626
rect 20253 6568 20258 6624
rect 20314 6568 22800 6624
rect 20253 6566 22800 6568
rect 20253 6563 20319 6566
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 22320 6536 22800 6566
rect 18104 6495 18424 6496
rect 20253 6082 20319 6085
rect 22320 6082 22800 6112
rect 20253 6080 22800 6082
rect 20253 6024 20258 6080
rect 20314 6024 22800 6080
rect 20253 6022 22800 6024
rect 20253 6019 20319 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 22320 5992 22800 6022
rect 14672 5951 14992 5952
rect 20621 5674 20687 5677
rect 22320 5674 22800 5704
rect 20621 5672 22800 5674
rect 20621 5616 20626 5672
rect 20682 5616 22800 5672
rect 20621 5614 22800 5616
rect 20621 5611 20687 5614
rect 22320 5584 22800 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 10409 5266 10475 5269
rect 19793 5266 19859 5269
rect 10409 5264 19859 5266
rect 10409 5208 10414 5264
rect 10470 5208 19798 5264
rect 19854 5208 19859 5264
rect 10409 5206 19859 5208
rect 10409 5203 10475 5206
rect 19793 5203 19859 5206
rect 20529 5130 20595 5133
rect 22320 5130 22800 5160
rect 20529 5128 22800 5130
rect 20529 5072 20534 5128
rect 20590 5072 22800 5128
rect 20529 5070 22800 5072
rect 20529 5067 20595 5070
rect 22320 5040 22800 5070
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 19057 4722 19123 4725
rect 22320 4722 22800 4752
rect 19057 4720 22800 4722
rect 19057 4664 19062 4720
rect 19118 4664 22800 4720
rect 19057 4662 22800 4664
rect 19057 4659 19123 4662
rect 22320 4632 22800 4662
rect 7557 4586 7623 4589
rect 9581 4586 9647 4589
rect 7557 4584 9647 4586
rect 7557 4528 7562 4584
rect 7618 4528 9586 4584
rect 9642 4528 9647 4584
rect 7557 4526 9647 4528
rect 7557 4523 7623 4526
rect 9581 4523 9647 4526
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 19057 4314 19123 4317
rect 22320 4314 22800 4344
rect 19057 4312 22800 4314
rect 19057 4256 19062 4312
rect 19118 4256 22800 4312
rect 19057 4254 22800 4256
rect 19057 4251 19123 4254
rect 22320 4224 22800 4254
rect 14089 4042 14155 4045
rect 18413 4042 18479 4045
rect 14089 4040 18479 4042
rect 14089 3984 14094 4040
rect 14150 3984 18418 4040
rect 18474 3984 18479 4040
rect 14089 3982 18479 3984
rect 14089 3979 14155 3982
rect 18413 3979 18479 3982
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 17125 3770 17191 3773
rect 18229 3770 18295 3773
rect 17125 3768 18295 3770
rect 17125 3712 17130 3768
rect 17186 3712 18234 3768
rect 18290 3712 18295 3768
rect 17125 3710 18295 3712
rect 17125 3707 17191 3710
rect 18229 3707 18295 3710
rect 18597 3770 18663 3773
rect 22320 3770 22800 3800
rect 18597 3768 22800 3770
rect 18597 3712 18602 3768
rect 18658 3712 22800 3768
rect 18597 3710 22800 3712
rect 18597 3707 18663 3710
rect 22320 3680 22800 3710
rect 18045 3498 18111 3501
rect 18045 3496 18568 3498
rect 18045 3440 18050 3496
rect 18106 3440 18568 3496
rect 18045 3438 18568 3440
rect 18045 3435 18111 3438
rect 18508 3362 18568 3438
rect 22320 3362 22800 3392
rect 18508 3302 22800 3362
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 22320 3272 22800 3302
rect 18104 3231 18424 3232
rect 19241 3090 19307 3093
rect 19198 3088 19307 3090
rect 19198 3032 19246 3088
rect 19302 3032 19307 3088
rect 19198 3027 19307 3032
rect 17769 2954 17835 2957
rect 19198 2954 19258 3027
rect 22320 2954 22800 2984
rect 17769 2952 22800 2954
rect 17769 2896 17774 2952
rect 17830 2896 22800 2952
rect 17769 2894 22800 2896
rect 17769 2891 17835 2894
rect 22320 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 20529 2410 20595 2413
rect 22320 2410 22800 2440
rect 20529 2408 22800 2410
rect 20529 2352 20534 2408
rect 20590 2352 22800 2408
rect 20529 2350 22800 2352
rect 20529 2347 20595 2350
rect 22320 2320 22800 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 17585 2002 17651 2005
rect 20989 2002 21055 2005
rect 22320 2002 22800 2032
rect 17585 2000 22800 2002
rect 17585 1944 17590 2000
rect 17646 1944 20994 2000
rect 21050 1944 22800 2000
rect 17585 1942 22800 1944
rect 17585 1939 17651 1942
rect 20989 1939 21055 1942
rect 22320 1912 22800 1942
rect 20621 1594 20687 1597
rect 22320 1594 22800 1624
rect 20621 1592 22800 1594
rect 20621 1536 20626 1592
rect 20682 1536 22800 1592
rect 20621 1534 22800 1536
rect 20621 1531 20687 1534
rect 22320 1504 22800 1534
rect 16389 1050 16455 1053
rect 22320 1050 22800 1080
rect 16389 1048 22800 1050
rect 16389 992 16394 1048
rect 16450 992 22800 1048
rect 16389 990 22800 992
rect 16389 987 16455 990
rect 22320 960 22800 990
rect 18965 642 19031 645
rect 22320 642 22800 672
rect 18965 640 22800 642
rect 18965 584 18970 640
rect 19026 584 22800 640
rect 18965 582 22800 584
rect 18965 579 19031 582
rect 22320 552 22800 582
rect 16573 234 16639 237
rect 22320 234 22800 264
rect 16573 232 22800 234
rect 16573 176 16578 232
rect 16634 176 22800 232
rect 16573 174 22800 176
rect 16573 171 16639 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7452 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_78
timestamp 1606256979
transform 1 0 8280 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1606256979
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9568 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10120 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1606256979
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_89
timestamp 1606256979
transform 1 0 9292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp 1606256979
transform 1 0 11040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1606256979
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _88_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606256979
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606256979
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12880 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12972 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_0_138
timestamp 1606256979
transform 1 0 13800 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1606256979
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1606256979
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1606256979
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1606256979
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1606256979
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15088 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606256979
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1606256979
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15824 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16100 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1606256979
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1606256979
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1606256979
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1606256979
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606256979
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606256979
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606256979
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606256979
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606256979
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19412 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1606256979
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1606256979
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1606256979
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1606256979
transform 1 0 18860 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1606256979
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1606256979
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606256979
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606256979
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606256979
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606256979
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1606256979
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606256979
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7176 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp 1606256979
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1606256979
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1606256979
transform 1 0 8832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1606256979
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1606256979
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11316 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_109
timestamp 1606256979
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13248 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1606256979
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_131
timestamp 1606256979
transform 1 0 13156 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1606256979
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1606256979
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 17480 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_170
timestamp 1606256979
transform 1 0 16744 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1606256979
transform 1 0 18308 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 18676 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19412 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1606256979
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_208
timestamp 1606256979
transform 1 0 20240 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_70
timestamp 1606256979
transform 1 0 7544 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1606256979
transform 1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10212 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1606256979
transform 1 0 9292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1606256979
transform 1 0 9660 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_97
timestamp 1606256979
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1606256979
transform 1 0 11776 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_108
timestamp 1606256979
transform 1 0 11040 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606256979
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_133
timestamp 1606256979
transform 1 0 13340 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15180 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_150
timestamp 1606256979
transform 1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606256979
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1606256979
transform 1 0 16652 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_177
timestamp 1606256979
transform 1 0 17388 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606256979
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1606256979
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606256979
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1606256979
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606256979
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606256979
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 1606256979
transform 1 0 6256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1606256979
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_74
timestamp 1606256979
transform 1 0 7912 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_80
timestamp 1606256979
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606256979
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1606256979
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_112
timestamp 1606256979
transform 1 0 11408 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1606256979
transform 1 0 12512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13800 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_136
timestamp 1606256979
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_147
timestamp 1606256979
transform 1 0 14628 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_166
timestamp 1606256979
transform 1 0 16376 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 17020 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_172
timestamp 1606256979
transform 1 0 16928 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1606256979
transform 1 0 18492 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1606256979
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606256979
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606256979
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_91
timestamp 1606256979
transform 1 0 9476 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1606256979
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606256979
transform 1 0 11776 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1606256979
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1606256979
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606256979
transform 1 0 13524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1606256979
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15916 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1606256979
transform 1 0 14812 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_170
timestamp 1606256979
transform 1 0 16744 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606256979
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 19044 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1606256979
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1606256979
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1606256979
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1606256979
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606256979
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5704 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_44
timestamp 1606256979
transform 1 0 5152 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606256979
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7820 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1606256979
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1606256979
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1606256979
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1606256979
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606256979
transform 1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_96
timestamp 1606256979
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10120 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10396 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9476 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11408 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1606256979
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1606256979
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606256979
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13064 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13156 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1606256979
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_140
timestamp 1606256979
transform 1 0 13984 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_146
timestamp 1606256979
transform 1 0 14536 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1606256979
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_146
timestamp 1606256979
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_163
timestamp 1606256979
transform 1 0 16100 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1606256979
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16284 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14628 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1606256979
transform 1 0 17388 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1606256979
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17848 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_174
timestamp 1606256979
transform 1 0 17112 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1606256979
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp 1606256979
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18768 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1606256979
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_202
timestamp 1606256979
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1606256979
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp 1606256979
transform 1 0 20240 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606256979
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1606256979
transform 1 0 20884 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1606256979
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606256979
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606256979
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606256979
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606256979
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1606256979
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10672 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1606256979
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606256979
transform 1 0 12328 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1606256979
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_125
timestamp 1606256979
transform 1 0 12604 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13432 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_133
timestamp 1606256979
transform 1 0 13340 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_143
timestamp 1606256979
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606256979
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17940 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1606256979
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19596 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1606256979
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1606256979
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606256979
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606256979
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606256979
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606256979
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1606256979
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1606256979
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_98
timestamp 1606256979
transform 1 0 10120 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1606256979
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606256979
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_139
timestamp 1606256979
transform 1 0 13892 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15456 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1606256979
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 17112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1606256979
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1606256979
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1606256979
transform 1 0 20240 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19228 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_196
timestamp 1606256979
transform 1 0 19136 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1606256979
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_211
timestamp 1606256979
transform 1 0 20516 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606256979
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606256979
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606256979
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606256979
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_68
timestamp 1606256979
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10580 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10120 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1606256979
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1606256979
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_112
timestamp 1606256979
transform 1 0 11408 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1606256979
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16192 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1606256979
transform 1 0 15732 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1606256979
transform 1 0 16100 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17204 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1606256979
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_181
timestamp 1606256979
transform 1 0 17756 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18768 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp 1606256979
transform 1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_201
timestamp 1606256979
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1606256979
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606256979
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606256979
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606256979
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606256979
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8556 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1606256979
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_80
timestamp 1606256979
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10212 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1606256979
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1606256979
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1606256979
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606256979
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12696 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15916 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15364 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_177
timestamp 1606256979
transform 1 0 17388 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19688 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18584 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_199
timestamp 1606256979
transform 1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_218
timestamp 1606256979
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606256979
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606256979
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606256979
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606256979
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606256979
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1606256979
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10764 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1606256979
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1606256979
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16376 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1606256979
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1606256979
transform 1 0 17388 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1606256979
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_180
timestamp 1606256979
transform 1 0 17664 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1606256979
transform 1 0 18584 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19044 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1606256979
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1606256979
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1606256979
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606256979
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606256979
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606256979
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606256979
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606256979
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606256979
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1606256979
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1606256979
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1606256979
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1606256979
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1606256979
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_98
timestamp 1606256979
transform 1 0 10120 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11132 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_106
timestamp 1606256979
transform 1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1606256979
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1606256979
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1606256979
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1606256979
transform 1 0 13064 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1606256979
transform 1 0 12972 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 1606256979
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_129
timestamp 1606256979
transform 1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1606256979
transform 1 0 14076 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1606256979
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15364 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1606256979
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1606256979
transform 1 0 14628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606256979
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1606256979
transform 1 0 17112 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17572 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1606256979
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1606256979
transform 1 0 16744 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_177
timestamp 1606256979
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606256979
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18400 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_204
timestamp 1606256979
transform 1 0 19872 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1606256979
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1606256979
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1606256979
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_210
timestamp 1606256979
transform 1 0 20424 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1606256979
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606256979
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606256979
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606256979
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1606256979
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1606256979
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1606256979
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1606256979
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1606256979
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1606256979
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1606256979
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1606256979
transform 1 0 12972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_141
timestamp 1606256979
transform 1 0 14076 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1606256979
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1606256979
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16560 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1606256979
transform 1 0 17388 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19044 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 20056 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1606256979
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1606256979
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1606256979
transform 1 0 20884 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1606256979
transform 1 0 21252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606256979
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606256979
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1606256979
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1606256979
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1606256979
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1606256979
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_117
timestamp 1606256979
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606256979
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_139
timestamp 1606256979
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1606256979
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606256979
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16836 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1606256979
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1606256979
transform 1 0 18308 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1606256979
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1606256979
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606256979
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606256979
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606256979
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606256979
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606256979
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606256979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1606256979
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1606256979
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1606256979
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1606256979
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13800 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12788 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1606256979
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15456 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1606256979
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_172
timestamp 1606256979
transform 1 0 16928 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1606256979
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18584 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 20240 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1606256979
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1606256979
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1606256979
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606256979
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1606256979
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1606256979
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1606256979
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606256979
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1606256979
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13340 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_129
timestamp 1606256979
transform 1 0 12972 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606256979
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15916 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606256979
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1606256979
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17572 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1606256979
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19412 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_195
timestamp 1606256979
transform 1 0 19044 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_205
timestamp 1606256979
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606256979
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606256979
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606256979
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606256979
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606256979
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606256979
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606256979
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606256979
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606256979
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606256979
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1606256979
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1606256979
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1606256979
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1606256979
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1606256979
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1606256979
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1606256979
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606256979
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606256979
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606256979
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1606256979
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1606256979
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15088 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1606256979
transform 1 0 14628 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_151
timestamp 1606256979
transform 1 0 14996 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_161
timestamp 1606256979
transform 1 0 15916 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606256979
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606256979
transform 1 0 17480 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1606256979
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 1606256979
transform 1 0 17388 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606256979
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606256979
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_194
timestamp 1606256979
transform 1 0 18952 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_190
timestamp 1606256979
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1606256979
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1606256979
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1606256979
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19596 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19596 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606256979
transform 1 0 19044 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 19044 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1606256979
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1606256979
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20332 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1606256979
transform 1 0 20884 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1606256979
transform 1 0 21252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1606256979
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1606256979
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1606256979
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606256979
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606256979
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1606256979
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1606256979
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_98
timestamp 1606256979
transform 1 0 10120 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10856 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_112
timestamp 1606256979
transform 1 0 11408 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1606256979
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606256979
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16100 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1606256979
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1606256979
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1606256979
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 19320 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 19872 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1606256979
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1606256979
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_216
timestamp 1606256979
transform 1 0 20976 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606256979
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1606256979
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_68
timestamp 1606256979
transform 1 0 7360 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_76
timestamp 1606256979
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1606256979
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1606256979
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1606256979
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1606256979
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1606256979
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1606256979
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1606256979
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1606256979
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1606256979
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1606256979
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1606256979
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606256979
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606256979
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606256979
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1606256979
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1606256979
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606256979
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1606256979
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9752 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_86
timestamp 1606256979
transform 1 0 9016 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_100
timestamp 1606256979
transform 1 0 10304 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_112
timestamp 1606256979
transform 1 0 11408 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606256979
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606256979
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1606256979
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1606256979
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1606256979
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp 1606256979
transform 1 0 19872 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1606256979
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606256979
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606256979
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606256979
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606256979
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1606256979
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1606256979
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1606256979
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1606256979
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11868 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606256979
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1606256979
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13800 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_135
timestamp 1606256979
transform 1 0 13524 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1606256979
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606256979
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606256979
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606256979
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606256979
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1606256979
transform 1 0 19688 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606256979
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606256979
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606256979
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606256979
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606256979
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606256979
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1606256979
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1606256979
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1606256979
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606256979
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1606256979
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1606256979
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1606256979
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19504 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1606256979
transform 1 0 19136 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1606256979
transform 1 0 20056 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_210
timestamp 1606256979
transform 1 0 20424 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606256979
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606256979
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606256979
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606256979
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1606256979
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1606256979
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606256979
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1606256979
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606256979
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606256979
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606256979
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1606256979
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1606256979
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1606256979
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606256979
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1606256979
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1606256979
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14168 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1606256979
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1606256979
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_135
timestamp 1606256979
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1606256979
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_166
timestamp 1606256979
transform 1 0 16376 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_148
timestamp 1606256979
transform 1 0 14720 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_160
timestamp 1606256979
transform 1 0 15824 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17020 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_172
timestamp 1606256979
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1606256979
transform 1 0 17572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_172
timestamp 1606256979
transform 1 0 16928 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1606256979
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 19964 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_191
timestamp 1606256979
transform 1 0 18676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1606256979
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1606256979
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1606256979
transform 1 0 19872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1606256979
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1606256979
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606256979
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606256979
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1606256979
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606256979
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606256979
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606256979
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1606256979
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1606256979
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11316 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_105
timestamp 1606256979
transform 1 0 10764 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1606256979
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1606256979
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1606256979
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1606256979
transform 1 0 15640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_170
timestamp 1606256979
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_182
timestamp 1606256979
transform 1 0 17848 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_194
timestamp 1606256979
transform 1 0 18952 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1606256979
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606256979
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606256979
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1606256979
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1606256979
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1606256979
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7728 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_70
timestamp 1606256979
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_78
timestamp 1606256979
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_90
timestamp 1606256979
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_102
timestamp 1606256979
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1606256979
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1606256979
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1606256979
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1606256979
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606256979
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 19964 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_196
timestamp 1606256979
transform 1 0 19136 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1606256979
transform 1 0 19872 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606256979
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1606256979
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606256979
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606256979
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1606256979
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1606256979
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606256979
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1606256979
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1606256979
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1606256979
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9752 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_93
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_100
timestamp 1606256979
transform 1 0 10304 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12144 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_112
timestamp 1606256979
transform 1 0 11408 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_126
timestamp 1606256979
transform 1 0 12696 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_138
timestamp 1606256979
transform 1 0 13800 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15640 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1606256979
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_164
timestamp 1606256979
transform 1 0 16192 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17664 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1606256979
transform 1 0 17296 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_186
timestamp 1606256979
transform 1 0 18216 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19596 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_198
timestamp 1606256979
transform 1 0 19320 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1606256979
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1606256979
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606256979
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1606256979
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1606256979
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1606256979
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606256979
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1606256979
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1606256979
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1606256979
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1606256979
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1606256979
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 16376 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1606256979
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_159
timestamp 1606256979
transform 1 0 15732 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_165
timestamp 1606256979
transform 1 0 16284 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_170
timestamp 1606256979
transform 1 0 16744 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1606256979
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606256979
transform 1 0 18492 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_188
timestamp 1606256979
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1606256979
transform 1 0 18860 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1606256979
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606256979
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606256979
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606256979
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606256979
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606256979
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606256979
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606256979
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606256979
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606256979
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606256979
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606256979
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606256979
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606256979
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606256979
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 5722 22320 5778 22800 6 SC_IN_TOP
port 0 nsew default input
rlabel metal2 s 22466 0 22522 480 6 SC_OUT_BOT
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_1_
port 2 nsew default input
rlabel metal2 s 17130 22320 17186 22800 6 ccff_head
port 3 nsew default input
rlabel metal3 s 0 11432 480 11552 6 ccff_tail
port 4 nsew default tristate
rlabel metal3 s 22320 3680 22800 3800 6 chanx_right_in[0]
port 5 nsew default input
rlabel metal3 s 22320 8304 22800 8424 6 chanx_right_in[10]
port 6 nsew default input
rlabel metal3 s 22320 8712 22800 8832 6 chanx_right_in[11]
port 7 nsew default input
rlabel metal3 s 22320 9256 22800 9376 6 chanx_right_in[12]
port 8 nsew default input
rlabel metal3 s 22320 9664 22800 9784 6 chanx_right_in[13]
port 9 nsew default input
rlabel metal3 s 22320 10072 22800 10192 6 chanx_right_in[14]
port 10 nsew default input
rlabel metal3 s 22320 10616 22800 10736 6 chanx_right_in[15]
port 11 nsew default input
rlabel metal3 s 22320 11024 22800 11144 6 chanx_right_in[16]
port 12 nsew default input
rlabel metal3 s 22320 11568 22800 11688 6 chanx_right_in[17]
port 13 nsew default input
rlabel metal3 s 22320 11976 22800 12096 6 chanx_right_in[18]
port 14 nsew default input
rlabel metal3 s 22320 12384 22800 12504 6 chanx_right_in[19]
port 15 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal3 s 22320 4632 22800 4752 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal3 s 22320 5040 22800 5160 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal3 s 22320 5584 22800 5704 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal3 s 22320 5992 22800 6112 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal3 s 22320 6536 22800 6656 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal3 s 22320 6944 22800 7064 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal3 s 22320 7352 22800 7472 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal3 s 22320 7896 22800 8016 6 chanx_right_in[9]
port 24 nsew default input
rlabel metal3 s 22320 12928 22800 13048 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal3 s 22320 17416 22800 17536 6 chanx_right_out[10]
port 26 nsew default tristate
rlabel metal3 s 22320 17960 22800 18080 6 chanx_right_out[11]
port 27 nsew default tristate
rlabel metal3 s 22320 18368 22800 18488 6 chanx_right_out[12]
port 28 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[13]
port 29 nsew default tristate
rlabel metal3 s 22320 19320 22800 19440 6 chanx_right_out[14]
port 30 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[15]
port 31 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[16]
port 32 nsew default tristate
rlabel metal3 s 22320 20680 22800 20800 6 chanx_right_out[17]
port 33 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[18]
port 34 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[19]
port 35 nsew default tristate
rlabel metal3 s 22320 13336 22800 13456 6 chanx_right_out[1]
port 36 nsew default tristate
rlabel metal3 s 22320 13744 22800 13864 6 chanx_right_out[2]
port 37 nsew default tristate
rlabel metal3 s 22320 14288 22800 14408 6 chanx_right_out[3]
port 38 nsew default tristate
rlabel metal3 s 22320 14696 22800 14816 6 chanx_right_out[4]
port 39 nsew default tristate
rlabel metal3 s 22320 15104 22800 15224 6 chanx_right_out[5]
port 40 nsew default tristate
rlabel metal3 s 22320 15648 22800 15768 6 chanx_right_out[6]
port 41 nsew default tristate
rlabel metal3 s 22320 16056 22800 16176 6 chanx_right_out[7]
port 42 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[8]
port 43 nsew default tristate
rlabel metal3 s 22320 17008 22800 17128 6 chanx_right_out[9]
port 44 nsew default tristate
rlabel metal2 s 662 0 718 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[10]
port 46 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[11]
port 47 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[12]
port 48 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[13]
port 49 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chany_bottom_in[14]
port 50 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[15]
port 51 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[16]
port 52 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[17]
port 53 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[18]
port 54 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[19]
port 55 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 56 nsew default input
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_in[2]
port 57 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[3]
port 58 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[4]
port 59 nsew default input
rlabel metal2 s 3422 0 3478 480 6 chany_bottom_in[5]
port 60 nsew default input
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_in[6]
port 61 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[7]
port 62 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[8]
port 63 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chany_bottom_in[9]
port 64 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_out[0]
port 65 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[10]
port 66 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[11]
port 67 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[12]
port 68 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[13]
port 69 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[14]
port 70 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[15]
port 71 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[16]
port 72 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[17]
port 73 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[18]
port 74 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[19]
port 75 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_out[1]
port 76 nsew default tristate
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_out[2]
port 77 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[3]
port 78 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[4]
port 79 nsew default tristate
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_out[5]
port 80 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_out[6]
port 81 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[7]
port 82 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[8]
port 83 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[9]
port 84 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 prog_clk_0_E_in
port 85 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 86 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 87 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 88 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 89 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 90 nsew default input
rlabel metal3 s 22320 2320 22800 2440 6 right_bottom_grid_pin_39_
port 91 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 92 nsew default input
rlabel metal3 s 22320 3272 22800 3392 6 right_bottom_grid_pin_41_
port 93 nsew default input
rlabel metal3 s 22320 22448 22800 22568 6 right_top_grid_pin_1_
port 94 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 95 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 96 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
