magic
tech sky130A
magscale 1 2
timestamp 1604668539
<< locali >>
rect 21373 24599 21407 24701
rect 12081 21335 12115 21505
rect 15945 19363 15979 19465
rect 21925 16983 21959 17085
rect 16129 10999 16163 11237
rect 15209 10591 15243 10693
rect 21649 9367 21683 9605
rect 12081 8415 12115 8585
rect 22845 5083 22879 5185
rect 19349 3927 19383 4029
<< viali >>
rect 14473 25449 14507 25483
rect 16865 25449 16899 25483
rect 19625 25449 19659 25483
rect 22201 25449 22235 25483
rect 14289 25313 14323 25347
rect 15577 25313 15611 25347
rect 16681 25313 16715 25347
rect 19441 25313 19475 25347
rect 22017 25313 22051 25347
rect 15301 25245 15335 25279
rect 15761 25177 15795 25211
rect 16221 25109 16255 25143
rect 18153 25109 18187 25143
rect 22017 24837 22051 24871
rect 16037 24769 16071 24803
rect 17509 24769 17543 24803
rect 18705 24769 18739 24803
rect 13185 24701 13219 24735
rect 13737 24701 13771 24735
rect 14289 24701 14323 24735
rect 14841 24701 14875 24735
rect 16957 24701 16991 24735
rect 18429 24701 18463 24735
rect 19901 24701 19935 24735
rect 20453 24701 20487 24735
rect 21005 24701 21039 24735
rect 21373 24701 21407 24735
rect 22201 24701 22235 24735
rect 22753 24701 22787 24735
rect 14197 24633 14231 24667
rect 15209 24633 15243 24667
rect 15853 24633 15887 24667
rect 17877 24633 17911 24667
rect 18521 24633 18555 24667
rect 19533 24633 19567 24667
rect 13369 24565 13403 24599
rect 14473 24565 14507 24599
rect 15393 24565 15427 24599
rect 15761 24565 15795 24599
rect 16773 24565 16807 24599
rect 18061 24565 18095 24599
rect 20085 24565 20119 24599
rect 21189 24565 21223 24599
rect 21373 24565 21407 24599
rect 21649 24565 21683 24599
rect 22385 24565 22419 24599
rect 23673 24565 23707 24599
rect 16313 24361 16347 24395
rect 19809 24361 19843 24395
rect 21465 24361 21499 24395
rect 21925 24361 21959 24395
rect 22569 24361 22603 24395
rect 23673 24361 23707 24395
rect 24777 24361 24811 24395
rect 15485 24293 15519 24327
rect 12173 24225 12207 24259
rect 13277 24225 13311 24259
rect 13737 24225 13771 24259
rect 16221 24225 16255 24259
rect 17693 24225 17727 24259
rect 18153 24225 18187 24259
rect 19625 24225 19659 24259
rect 21281 24225 21315 24259
rect 22385 24225 22419 24259
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 12265 24157 12299 24191
rect 12449 24157 12483 24191
rect 13829 24157 13863 24191
rect 14013 24157 14047 24191
rect 16405 24157 16439 24191
rect 18245 24157 18279 24191
rect 18429 24157 18463 24191
rect 12909 24089 12943 24123
rect 15853 24089 15887 24123
rect 11345 24021 11379 24055
rect 11805 24021 11839 24055
rect 13369 24021 13403 24055
rect 15025 24021 15059 24055
rect 17785 24021 17819 24055
rect 18889 24021 18923 24055
rect 11437 23817 11471 23851
rect 11805 23817 11839 23851
rect 14933 23817 14967 23851
rect 16037 23817 16071 23851
rect 16313 23817 16347 23851
rect 17049 23817 17083 23851
rect 24777 23817 24811 23851
rect 15577 23681 15611 23715
rect 18889 23681 18923 23715
rect 21925 23681 21959 23715
rect 25145 23681 25179 23715
rect 11253 23613 11287 23647
rect 12449 23613 12483 23647
rect 12716 23613 12750 23647
rect 14841 23613 14875 23647
rect 15393 23613 15427 23647
rect 16865 23613 16899 23647
rect 17417 23613 17451 23647
rect 21833 23613 21867 23647
rect 24593 23613 24627 23647
rect 11161 23545 11195 23579
rect 17877 23545 17911 23579
rect 18429 23545 18463 23579
rect 19156 23545 19190 23579
rect 21741 23545 21775 23579
rect 12173 23477 12207 23511
rect 13829 23477 13863 23511
rect 14381 23477 14415 23511
rect 15301 23477 15335 23511
rect 16681 23477 16715 23511
rect 18705 23477 18739 23511
rect 20269 23477 20303 23511
rect 20821 23477 20855 23511
rect 21189 23477 21223 23511
rect 21373 23477 21407 23511
rect 22385 23477 22419 23511
rect 23857 23477 23891 23511
rect 24409 23477 24443 23511
rect 13001 23273 13035 23307
rect 13461 23273 13495 23307
rect 15577 23273 15611 23307
rect 17141 23273 17175 23307
rect 17693 23273 17727 23307
rect 18153 23273 18187 23307
rect 19625 23273 19659 23307
rect 21373 23273 21407 23307
rect 23397 23273 23431 23307
rect 24041 23273 24075 23307
rect 24777 23273 24811 23307
rect 12633 23205 12667 23239
rect 16028 23205 16062 23239
rect 10876 23137 10910 23171
rect 15761 23137 15795 23171
rect 18245 23137 18279 23171
rect 18501 23137 18535 23171
rect 21281 23137 21315 23171
rect 24593 23137 24627 23171
rect 10609 23069 10643 23103
rect 13553 23069 13587 23103
rect 13645 23069 13679 23103
rect 14197 23069 14231 23103
rect 21465 23069 21499 23103
rect 23489 23069 23523 23103
rect 23673 23069 23707 23103
rect 24409 23069 24443 23103
rect 20913 23001 20947 23035
rect 11989 22933 12023 22967
rect 13093 22933 13127 22967
rect 14933 22933 14967 22967
rect 21925 22933 21959 22967
rect 23029 22933 23063 22967
rect 10977 22729 11011 22763
rect 13829 22729 13863 22763
rect 14381 22729 14415 22763
rect 15945 22729 15979 22763
rect 16405 22729 16439 22763
rect 17049 22729 17083 22763
rect 17509 22729 17543 22763
rect 18061 22729 18095 22763
rect 19073 22729 19107 22763
rect 19993 22729 20027 22763
rect 21557 22729 21591 22763
rect 23029 22729 23063 22763
rect 25421 22729 25455 22763
rect 17785 22661 17819 22695
rect 19441 22661 19475 22695
rect 22753 22661 22787 22695
rect 10701 22593 10735 22627
rect 12265 22593 12299 22627
rect 12449 22593 12483 22627
rect 15577 22593 15611 22627
rect 18521 22593 18555 22627
rect 18613 22593 18647 22627
rect 20177 22593 20211 22627
rect 22201 22593 22235 22627
rect 24225 22593 24259 22627
rect 16865 22525 16899 22559
rect 18429 22525 18463 22559
rect 24041 22525 24075 22559
rect 12716 22457 12750 22491
rect 14841 22457 14875 22491
rect 20422 22457 20456 22491
rect 24133 22457 24167 22491
rect 14933 22389 14967 22423
rect 15301 22389 15335 22423
rect 15393 22389 15427 22423
rect 23489 22389 23523 22423
rect 23673 22389 23707 22423
rect 24685 22389 24719 22423
rect 12909 22185 12943 22219
rect 15393 22185 15427 22219
rect 18153 22185 18187 22219
rect 18981 22185 19015 22219
rect 20269 22185 20303 22219
rect 20729 22185 20763 22219
rect 21649 22185 21683 22219
rect 22661 22185 22695 22219
rect 23029 22185 23063 22219
rect 13277 22117 13311 22151
rect 15761 22117 15795 22151
rect 13369 22049 13403 22083
rect 13921 22049 13955 22083
rect 17325 22049 17359 22083
rect 21097 22049 21131 22083
rect 22109 22049 22143 22083
rect 23388 22049 23422 22083
rect 12541 21981 12575 22015
rect 13461 21981 13495 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 17417 21981 17451 22015
rect 17601 21981 17635 22015
rect 19073 21981 19107 22015
rect 19165 21981 19199 22015
rect 22017 21981 22051 22015
rect 23121 21981 23155 22015
rect 18521 21913 18555 21947
rect 10885 21845 10919 21879
rect 12173 21845 12207 21879
rect 15025 21845 15059 21879
rect 16957 21845 16991 21879
rect 18613 21845 18647 21879
rect 19625 21845 19659 21879
rect 21281 21845 21315 21879
rect 22293 21845 22327 21879
rect 24501 21845 24535 21879
rect 10609 21641 10643 21675
rect 13461 21641 13495 21675
rect 14749 21641 14783 21675
rect 15945 21641 15979 21675
rect 16313 21641 16347 21675
rect 16865 21641 16899 21675
rect 17417 21641 17451 21675
rect 18889 21641 18923 21675
rect 20453 21641 20487 21675
rect 22017 21641 22051 21675
rect 21925 21573 21959 21607
rect 11253 21505 11287 21539
rect 11437 21505 11471 21539
rect 12081 21505 12115 21539
rect 13093 21505 13127 21539
rect 14473 21505 14507 21539
rect 15485 21505 15519 21539
rect 19073 21505 19107 21539
rect 21557 21505 21591 21539
rect 22477 21505 22511 21539
rect 22569 21505 22603 21539
rect 11897 21369 11931 21403
rect 15301 21437 15335 21471
rect 19340 21437 19374 21471
rect 22385 21437 22419 21471
rect 24133 21437 24167 21471
rect 24389 21437 24423 21471
rect 12909 21369 12943 21403
rect 15393 21369 15427 21403
rect 10793 21301 10827 21335
rect 11161 21301 11195 21335
rect 12081 21301 12115 21335
rect 12173 21301 12207 21335
rect 12449 21301 12483 21335
rect 12817 21301 12851 21335
rect 14013 21301 14047 21335
rect 14933 21301 14967 21335
rect 16957 21301 16991 21335
rect 17785 21301 17819 21335
rect 18061 21301 18095 21335
rect 18521 21301 18555 21335
rect 21189 21301 21223 21335
rect 23121 21301 23155 21335
rect 23949 21301 23983 21335
rect 25513 21301 25547 21335
rect 13369 21097 13403 21131
rect 13829 21097 13863 21131
rect 13921 21097 13955 21131
rect 15025 21097 15059 21131
rect 17141 21097 17175 21131
rect 17325 21097 17359 21131
rect 19349 21097 19383 21131
rect 19901 21097 19935 21131
rect 21741 21097 21775 21131
rect 23213 21097 23247 21131
rect 23765 21097 23799 21131
rect 11704 21029 11738 21063
rect 17785 21029 17819 21063
rect 18705 21029 18739 21063
rect 24685 21029 24719 21063
rect 1409 20961 1443 20995
rect 15761 20961 15795 20995
rect 16865 20961 16899 20995
rect 17693 20961 17727 20995
rect 19257 20961 19291 20995
rect 22100 20961 22134 20995
rect 11437 20893 11471 20927
rect 15853 20893 15887 20927
rect 16037 20893 16071 20927
rect 17877 20893 17911 20927
rect 19533 20893 19567 20927
rect 21833 20893 21867 20927
rect 24777 20893 24811 20927
rect 24961 20893 24995 20927
rect 1593 20825 1627 20859
rect 10885 20757 10919 20791
rect 12817 20757 12851 20791
rect 15393 20757 15427 20791
rect 18889 20757 18923 20791
rect 20545 20757 20579 20791
rect 24133 20757 24167 20791
rect 24317 20757 24351 20791
rect 11253 20553 11287 20587
rect 12449 20553 12483 20587
rect 16129 20553 16163 20587
rect 17049 20553 17083 20587
rect 19441 20553 19475 20587
rect 20085 20553 20119 20587
rect 22201 20553 22235 20587
rect 23489 20553 23523 20587
rect 25513 20553 25547 20587
rect 25881 20553 25915 20587
rect 12909 20417 12943 20451
rect 13093 20417 13127 20451
rect 21097 20417 21131 20451
rect 24777 20417 24811 20451
rect 1409 20349 1443 20383
rect 13829 20349 13863 20383
rect 14749 20349 14783 20383
rect 17877 20349 17911 20383
rect 18061 20349 18095 20383
rect 20453 20349 20487 20383
rect 21005 20349 21039 20383
rect 22569 20349 22603 20383
rect 24501 20349 24535 20383
rect 12265 20281 12299 20315
rect 12817 20281 12851 20315
rect 14994 20281 15028 20315
rect 17509 20281 17543 20315
rect 18328 20281 18362 20315
rect 24593 20281 24627 20315
rect 1593 20213 1627 20247
rect 1961 20213 1995 20247
rect 10333 20213 10367 20247
rect 11345 20213 11379 20247
rect 11897 20213 11931 20247
rect 13461 20213 13495 20247
rect 14197 20213 14231 20247
rect 14565 20213 14599 20247
rect 16681 20213 16715 20247
rect 20545 20213 20579 20247
rect 20913 20213 20947 20247
rect 21833 20213 21867 20247
rect 23949 20213 23983 20247
rect 24133 20213 24167 20247
rect 25145 20213 25179 20247
rect 14105 20009 14139 20043
rect 17509 20009 17543 20043
rect 18061 20009 18095 20043
rect 18705 20009 18739 20043
rect 20085 20009 20119 20043
rect 20637 20009 20671 20043
rect 22293 20009 22327 20043
rect 23857 20009 23891 20043
rect 12992 19941 13026 19975
rect 15752 19941 15786 19975
rect 19165 19941 19199 19975
rect 24216 19941 24250 19975
rect 10241 19873 10275 19907
rect 10497 19873 10531 19907
rect 12725 19873 12759 19907
rect 14841 19873 14875 19907
rect 15485 19873 15519 19907
rect 18613 19873 18647 19907
rect 19073 19873 19107 19907
rect 19809 19873 19843 19907
rect 21169 19873 21203 19907
rect 23949 19873 23983 19907
rect 19349 19805 19383 19839
rect 20913 19805 20947 19839
rect 1593 19669 1627 19703
rect 11621 19669 11655 19703
rect 12541 19669 12575 19703
rect 16865 19669 16899 19703
rect 25329 19669 25363 19703
rect 9505 19465 9539 19499
rect 13553 19465 13587 19499
rect 14105 19465 14139 19499
rect 15945 19465 15979 19499
rect 16497 19465 16531 19499
rect 18061 19465 18095 19499
rect 21281 19465 21315 19499
rect 22293 19465 22327 19499
rect 25053 19465 25087 19499
rect 9873 19397 9907 19431
rect 16129 19397 16163 19431
rect 20913 19397 20947 19431
rect 10977 19329 11011 19363
rect 11345 19329 11379 19363
rect 13093 19329 13127 19363
rect 14197 19329 14231 19363
rect 15945 19329 15979 19363
rect 17509 19329 17543 19363
rect 18705 19329 18739 19363
rect 20269 19329 20303 19363
rect 21925 19329 21959 19363
rect 24593 19329 24627 19363
rect 10149 19261 10183 19295
rect 10701 19261 10735 19295
rect 11897 19261 11931 19295
rect 12817 19261 12851 19295
rect 16681 19261 16715 19295
rect 18429 19261 18463 19295
rect 20085 19261 20119 19295
rect 23121 19261 23155 19295
rect 24317 19261 24351 19295
rect 25513 19261 25547 19295
rect 26065 19261 26099 19295
rect 12265 19193 12299 19227
rect 14464 19193 14498 19227
rect 21741 19193 21775 19227
rect 23489 19193 23523 19227
rect 24409 19193 24443 19227
rect 25329 19193 25363 19227
rect 10333 19125 10367 19159
rect 10793 19125 10827 19159
rect 12449 19125 12483 19159
rect 12909 19125 12943 19159
rect 15577 19125 15611 19159
rect 16865 19125 16899 19159
rect 17877 19125 17911 19159
rect 18521 19125 18555 19159
rect 19165 19125 19199 19159
rect 19533 19125 19567 19159
rect 19717 19125 19751 19159
rect 20177 19125 20211 19159
rect 21649 19125 21683 19159
rect 22753 19125 22787 19159
rect 23949 19125 23983 19159
rect 25697 19125 25731 19159
rect 12817 18921 12851 18955
rect 13185 18921 13219 18955
rect 13645 18921 13679 18955
rect 14013 18921 14047 18955
rect 14657 18921 14691 18955
rect 15393 18921 15427 18955
rect 16773 18921 16807 18955
rect 18521 18921 18555 18955
rect 19533 18921 19567 18955
rect 20637 18921 20671 18955
rect 21189 18921 21223 18955
rect 22569 18921 22603 18955
rect 23673 18921 23707 18955
rect 14105 18853 14139 18887
rect 15761 18853 15795 18887
rect 16405 18853 16439 18887
rect 21557 18853 21591 18887
rect 24124 18853 24158 18887
rect 10957 18785 10991 18819
rect 15853 18785 15887 18819
rect 17408 18785 17442 18819
rect 19165 18785 19199 18819
rect 19809 18785 19843 18819
rect 10701 18717 10735 18751
rect 14197 18717 14231 18751
rect 16037 18717 16071 18751
rect 17141 18717 17175 18751
rect 21649 18717 21683 18751
rect 21741 18717 21775 18751
rect 22845 18717 22879 18751
rect 23857 18717 23891 18751
rect 10425 18581 10459 18615
rect 12081 18581 12115 18615
rect 15025 18581 15059 18615
rect 19993 18581 20027 18615
rect 22201 18581 22235 18615
rect 25237 18581 25271 18615
rect 10333 18377 10367 18411
rect 10609 18377 10643 18411
rect 14197 18377 14231 18411
rect 15761 18377 15795 18411
rect 16405 18377 16439 18411
rect 17693 18377 17727 18411
rect 20361 18377 20395 18411
rect 22845 18377 22879 18411
rect 23397 18377 23431 18411
rect 24685 18377 24719 18411
rect 25145 18377 25179 18411
rect 11805 18309 11839 18343
rect 16681 18309 16715 18343
rect 17325 18309 17359 18343
rect 18797 18309 18831 18343
rect 11253 18241 11287 18275
rect 11437 18241 11471 18275
rect 12265 18241 12299 18275
rect 13369 18241 13403 18275
rect 13921 18241 13955 18275
rect 18981 18241 19015 18275
rect 22109 18241 22143 18275
rect 22477 18241 22511 18275
rect 24133 18241 24167 18275
rect 24317 18241 24351 18275
rect 9965 18173 9999 18207
rect 13185 18173 13219 18207
rect 14381 18173 14415 18207
rect 16865 18173 16899 18207
rect 18245 18173 18279 18207
rect 21189 18173 21223 18207
rect 24041 18173 24075 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 12725 18105 12759 18139
rect 13277 18105 13311 18139
rect 14626 18105 14660 18139
rect 19226 18105 19260 18139
rect 21925 18105 21959 18139
rect 10793 18037 10827 18071
rect 11161 18037 11195 18071
rect 12817 18037 12851 18071
rect 17049 18037 17083 18071
rect 21465 18037 21499 18071
rect 21833 18037 21867 18071
rect 23673 18037 23707 18071
rect 25421 18037 25455 18071
rect 13737 17833 13771 17867
rect 15761 17833 15795 17867
rect 16313 17833 16347 17867
rect 19993 17833 20027 17867
rect 20361 17833 20395 17867
rect 21925 17833 21959 17867
rect 23121 17833 23155 17867
rect 23673 17833 23707 17867
rect 24225 17833 24259 17867
rect 11498 17765 11532 17799
rect 15669 17765 15703 17799
rect 17224 17765 17258 17799
rect 21373 17765 21407 17799
rect 11253 17697 11287 17731
rect 16957 17697 16991 17731
rect 19809 17697 19843 17731
rect 21281 17697 21315 17731
rect 23581 17697 23615 17731
rect 24777 17697 24811 17731
rect 10885 17629 10919 17663
rect 14197 17629 14231 17663
rect 15853 17629 15887 17663
rect 21557 17629 21591 17663
rect 23765 17629 23799 17663
rect 15025 17561 15059 17595
rect 20913 17561 20947 17595
rect 23213 17561 23247 17595
rect 12633 17493 12667 17527
rect 14749 17493 14783 17527
rect 15301 17493 15335 17527
rect 18337 17493 18371 17527
rect 19073 17493 19107 17527
rect 22293 17493 22327 17527
rect 24961 17493 24995 17527
rect 11805 17289 11839 17323
rect 12173 17289 12207 17323
rect 13829 17289 13863 17323
rect 14473 17289 14507 17323
rect 16313 17289 16347 17323
rect 17049 17289 17083 17323
rect 17417 17289 17451 17323
rect 20545 17289 20579 17323
rect 21097 17289 21131 17323
rect 22477 17289 22511 17323
rect 25053 17289 25087 17323
rect 25605 17289 25639 17323
rect 18429 17221 18463 17255
rect 23397 17221 23431 17255
rect 10333 17153 10367 17187
rect 11437 17153 11471 17187
rect 18613 17153 18647 17187
rect 21005 17153 21039 17187
rect 21649 17153 21683 17187
rect 22845 17153 22879 17187
rect 23673 17153 23707 17187
rect 10701 17085 10735 17119
rect 12449 17085 12483 17119
rect 12716 17085 12750 17119
rect 14933 17085 14967 17119
rect 15189 17085 15223 17119
rect 21465 17085 21499 17119
rect 21925 17085 21959 17119
rect 23940 17085 23974 17119
rect 11161 17017 11195 17051
rect 14841 17017 14875 17051
rect 18880 17017 18914 17051
rect 10793 16949 10827 16983
rect 11253 16949 11287 16983
rect 19993 16949 20027 16983
rect 21557 16949 21591 16983
rect 21925 16949 21959 16983
rect 22109 16949 22143 16983
rect 11253 16745 11287 16779
rect 11345 16745 11379 16779
rect 12541 16745 12575 16779
rect 14381 16745 14415 16779
rect 15025 16745 15059 16779
rect 15301 16745 15335 16779
rect 16405 16745 16439 16779
rect 18889 16745 18923 16779
rect 20361 16745 20395 16779
rect 22293 16745 22327 16779
rect 22937 16745 22971 16779
rect 23397 16745 23431 16779
rect 24501 16745 24535 16779
rect 25145 16745 25179 16779
rect 11713 16677 11747 16711
rect 15761 16677 15795 16711
rect 17132 16677 17166 16711
rect 23213 16677 23247 16711
rect 23765 16677 23799 16711
rect 10885 16609 10919 16643
rect 14197 16609 14231 16643
rect 15669 16609 15703 16643
rect 16865 16609 16899 16643
rect 19809 16609 19843 16643
rect 21169 16609 21203 16643
rect 24961 16609 24995 16643
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 15853 16541 15887 16575
rect 20913 16541 20947 16575
rect 23857 16541 23891 16575
rect 24041 16541 24075 16575
rect 18245 16405 18279 16439
rect 20637 16405 20671 16439
rect 11161 16201 11195 16235
rect 11897 16201 11931 16235
rect 13829 16201 13863 16235
rect 14657 16201 14691 16235
rect 15761 16201 15795 16235
rect 16221 16201 16255 16235
rect 17417 16201 17451 16235
rect 20177 16201 20211 16235
rect 21557 16201 21591 16235
rect 23857 16201 23891 16235
rect 24225 16201 24259 16235
rect 25513 16201 25547 16235
rect 12173 16133 12207 16167
rect 21189 16133 21223 16167
rect 11345 16065 11379 16099
rect 14197 16065 14231 16099
rect 15209 16065 15243 16099
rect 16865 16065 16899 16099
rect 17049 16065 17083 16099
rect 18521 16065 18555 16099
rect 19165 16065 19199 16099
rect 19717 16065 19751 16099
rect 20729 16065 20763 16099
rect 22201 16065 22235 16099
rect 22385 16065 22419 16099
rect 22753 16065 22787 16099
rect 12449 15997 12483 16031
rect 12909 15997 12943 16031
rect 15117 15997 15151 16031
rect 16773 15997 16807 16031
rect 20545 15997 20579 16031
rect 22109 15997 22143 16031
rect 24593 15997 24627 16031
rect 25145 15997 25179 16031
rect 14473 15929 14507 15963
rect 17877 15929 17911 15963
rect 18981 15929 19015 15963
rect 12633 15861 12667 15895
rect 15025 15861 15059 15895
rect 16405 15861 16439 15895
rect 18613 15861 18647 15895
rect 19073 15861 19107 15895
rect 19993 15861 20027 15895
rect 20637 15861 20671 15895
rect 21741 15861 21775 15895
rect 23397 15861 23431 15895
rect 24777 15861 24811 15895
rect 14289 15657 14323 15691
rect 14657 15657 14691 15691
rect 15025 15657 15059 15691
rect 16681 15657 16715 15691
rect 17049 15657 17083 15691
rect 19165 15657 19199 15691
rect 20177 15657 20211 15691
rect 21097 15657 21131 15691
rect 22753 15657 22787 15691
rect 21618 15589 21652 15623
rect 15945 15521 15979 15555
rect 17141 15521 17175 15555
rect 17408 15521 17442 15555
rect 24593 15521 24627 15555
rect 16037 15453 16071 15487
rect 16221 15453 16255 15487
rect 19625 15453 19659 15487
rect 21373 15453 21407 15487
rect 24777 15385 24811 15419
rect 15577 15317 15611 15351
rect 18521 15317 18555 15351
rect 14749 15113 14783 15147
rect 16221 15113 16255 15147
rect 17233 15113 17267 15147
rect 18337 15113 18371 15147
rect 21649 15113 21683 15147
rect 22293 15113 22327 15147
rect 22661 15113 22695 15147
rect 24409 15113 24443 15147
rect 21925 15045 21959 15079
rect 15117 14977 15151 15011
rect 16681 14977 16715 15011
rect 16773 14977 16807 15011
rect 18521 14977 18555 15011
rect 13001 14909 13035 14943
rect 13461 14909 13495 14943
rect 16129 14909 16163 14943
rect 17601 14909 17635 14943
rect 21465 14909 21499 14943
rect 22477 14909 22511 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 16589 14841 16623 14875
rect 18766 14841 18800 14875
rect 13185 14773 13219 14807
rect 14381 14773 14415 14807
rect 15209 14773 15243 14807
rect 15669 14773 15703 14807
rect 19901 14773 19935 14807
rect 21373 14773 21407 14807
rect 23121 14773 23155 14807
rect 24777 14773 24811 14807
rect 15669 14569 15703 14603
rect 17417 14569 17451 14603
rect 18061 14569 18095 14603
rect 19441 14569 19475 14603
rect 21465 14569 21499 14603
rect 23213 14569 23247 14603
rect 24961 14569 24995 14603
rect 15117 14501 15151 14535
rect 16282 14501 16316 14535
rect 13093 14433 13127 14467
rect 14105 14433 14139 14467
rect 16037 14433 16071 14467
rect 20913 14433 20947 14467
rect 22017 14433 22051 14467
rect 23581 14433 23615 14467
rect 23673 14433 23707 14467
rect 24777 14433 24811 14467
rect 18981 14365 19015 14399
rect 19533 14365 19567 14399
rect 19625 14365 19659 14399
rect 23857 14365 23891 14399
rect 14289 14297 14323 14331
rect 20085 14297 20119 14331
rect 13277 14229 13311 14263
rect 18521 14229 18555 14263
rect 19073 14229 19107 14263
rect 21097 14229 21131 14263
rect 22201 14229 22235 14263
rect 23029 14229 23063 14263
rect 13093 14025 13127 14059
rect 13461 14025 13495 14059
rect 14197 14025 14231 14059
rect 14473 14025 14507 14059
rect 15669 14025 15703 14059
rect 17049 14025 17083 14059
rect 18061 14025 18095 14059
rect 19165 14025 19199 14059
rect 19533 14025 19567 14059
rect 23121 14025 23155 14059
rect 25053 14025 25087 14059
rect 25605 14025 25639 14059
rect 15209 13957 15243 13991
rect 16773 13957 16807 13991
rect 21557 13957 21591 13991
rect 22017 13957 22051 13991
rect 23397 13957 23431 13991
rect 16129 13889 16163 13923
rect 16313 13889 16347 13923
rect 18613 13889 18647 13923
rect 23673 13889 23707 13923
rect 13645 13821 13679 13855
rect 14657 13821 14691 13855
rect 15485 13821 15519 13855
rect 16037 13821 16071 13855
rect 17785 13821 17819 13855
rect 18521 13821 18555 13855
rect 19625 13821 19659 13855
rect 19881 13821 19915 13855
rect 22477 13821 22511 13855
rect 18429 13753 18463 13787
rect 23918 13753 23952 13787
rect 13829 13685 13863 13719
rect 14841 13685 14875 13719
rect 21005 13685 21039 13719
rect 22569 13685 22603 13719
rect 14381 13481 14415 13515
rect 15577 13481 15611 13515
rect 17601 13481 17635 13515
rect 18245 13481 18279 13515
rect 19165 13481 19199 13515
rect 23213 13481 23247 13515
rect 24777 13481 24811 13515
rect 16037 13413 16071 13447
rect 19625 13413 19659 13447
rect 23121 13413 23155 13447
rect 14197 13345 14231 13379
rect 15945 13345 15979 13379
rect 17509 13345 17543 13379
rect 19717 13345 19751 13379
rect 21281 13345 21315 13379
rect 24593 13345 24627 13379
rect 16221 13277 16255 13311
rect 17693 13277 17727 13311
rect 19901 13277 19935 13311
rect 21373 13277 21407 13311
rect 21557 13277 21591 13311
rect 23397 13277 23431 13311
rect 16681 13209 16715 13243
rect 17141 13209 17175 13243
rect 18797 13209 18831 13243
rect 19257 13209 19291 13243
rect 20913 13209 20947 13243
rect 22753 13209 22787 13243
rect 16957 13141 16991 13175
rect 20637 13141 20671 13175
rect 21925 13141 21959 13175
rect 22293 13141 22327 13175
rect 23765 13141 23799 13175
rect 14013 12937 14047 12971
rect 16405 12937 16439 12971
rect 16773 12937 16807 12971
rect 17601 12937 17635 12971
rect 20453 12937 20487 12971
rect 21925 12937 21959 12971
rect 22293 12937 22327 12971
rect 23121 12937 23155 12971
rect 24501 12937 24535 12971
rect 16129 12869 16163 12903
rect 20085 12869 20119 12903
rect 22845 12869 22879 12903
rect 14105 12801 14139 12835
rect 19533 12801 19567 12835
rect 21189 12801 21223 12835
rect 16589 12733 16623 12767
rect 18797 12733 18831 12767
rect 19349 12733 19383 12767
rect 20913 12733 20947 12767
rect 22109 12733 22143 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 13645 12665 13679 12699
rect 14350 12665 14384 12699
rect 19441 12665 19475 12699
rect 21005 12665 21039 12699
rect 13093 12597 13127 12631
rect 15485 12597 15519 12631
rect 17233 12597 17267 12631
rect 18429 12597 18463 12631
rect 18981 12597 19015 12631
rect 20545 12597 20579 12631
rect 21557 12597 21591 12631
rect 24777 12597 24811 12631
rect 12449 12393 12483 12427
rect 15117 12393 15151 12427
rect 16957 12393 16991 12427
rect 17509 12393 17543 12427
rect 18061 12393 18095 12427
rect 19257 12393 19291 12427
rect 19625 12393 19659 12427
rect 23765 12393 23799 12427
rect 12541 12325 12575 12359
rect 21364 12325 21398 12359
rect 14013 12257 14047 12291
rect 15844 12257 15878 12291
rect 18705 12257 18739 12291
rect 19717 12257 19751 12291
rect 21097 12257 21131 12291
rect 23581 12257 23615 12291
rect 24593 12257 24627 12291
rect 12633 12189 12667 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 15577 12189 15611 12223
rect 19901 12189 19935 12223
rect 17877 12121 17911 12155
rect 23121 12121 23155 12155
rect 12081 12053 12115 12087
rect 13645 12053 13679 12087
rect 14657 12053 14691 12087
rect 19073 12053 19107 12087
rect 20545 12053 20579 12087
rect 22477 12053 22511 12087
rect 24133 12053 24167 12087
rect 24777 12053 24811 12087
rect 11437 11849 11471 11883
rect 12173 11849 12207 11883
rect 13093 11849 13127 11883
rect 15577 11849 15611 11883
rect 16405 11849 16439 11883
rect 17785 11849 17819 11883
rect 20085 11849 20119 11883
rect 20453 11849 20487 11883
rect 21925 11849 21959 11883
rect 22753 11849 22787 11883
rect 24685 11849 24719 11883
rect 11805 11781 11839 11815
rect 16313 11781 16347 11815
rect 16865 11713 16899 11747
rect 16957 11713 16991 11747
rect 18061 11713 18095 11747
rect 23489 11713 23523 11747
rect 24133 11713 24167 11747
rect 24225 11713 24259 11747
rect 13461 11645 13495 11679
rect 13553 11645 13587 11679
rect 16773 11645 16807 11679
rect 20545 11645 20579 11679
rect 12725 11577 12759 11611
rect 13798 11577 13832 11611
rect 18306 11577 18340 11611
rect 20790 11577 20824 11611
rect 24041 11577 24075 11611
rect 14933 11509 14967 11543
rect 17417 11509 17451 11543
rect 19441 11509 19475 11543
rect 23029 11509 23063 11543
rect 23673 11509 23707 11543
rect 12173 11305 12207 11339
rect 13185 11305 13219 11339
rect 13645 11305 13679 11339
rect 14657 11305 14691 11339
rect 15301 11305 15335 11339
rect 18889 11305 18923 11339
rect 19625 11305 19659 11339
rect 19809 11305 19843 11339
rect 21097 11305 21131 11339
rect 21465 11305 21499 11339
rect 15669 11237 15703 11271
rect 16129 11237 16163 11271
rect 22538 11237 22572 11271
rect 25237 11237 25271 11271
rect 11989 11169 12023 11203
rect 14013 11169 14047 11203
rect 14105 11169 14139 11203
rect 15761 11169 15795 11203
rect 13553 11101 13587 11135
rect 14197 11101 14231 11135
rect 15025 11101 15059 11135
rect 15853 11101 15887 11135
rect 16865 11169 16899 11203
rect 17132 11169 17166 11203
rect 21273 11169 21307 11203
rect 22293 11169 22327 11203
rect 25145 11169 25179 11203
rect 21833 11101 21867 11135
rect 25421 11101 25455 11135
rect 16313 11033 16347 11067
rect 18245 11033 18279 11067
rect 19349 11033 19383 11067
rect 24777 11033 24811 11067
rect 1593 10965 1627 10999
rect 11345 10965 11379 10999
rect 12541 10965 12575 10999
rect 16129 10965 16163 10999
rect 16773 10965 16807 10999
rect 20545 10965 20579 10999
rect 22109 10965 22143 10999
rect 23673 10965 23707 10999
rect 24317 10965 24351 10999
rect 11253 10761 11287 10795
rect 11529 10761 11563 10795
rect 14013 10761 14047 10795
rect 15577 10761 15611 10795
rect 16865 10761 16899 10795
rect 17601 10761 17635 10795
rect 18245 10761 18279 10795
rect 21373 10761 21407 10795
rect 22385 10761 22419 10795
rect 22753 10761 22787 10795
rect 25973 10761 26007 10795
rect 12449 10693 12483 10727
rect 15025 10693 15059 10727
rect 15209 10693 15243 10727
rect 18705 10693 18739 10727
rect 23397 10693 23431 10727
rect 12265 10625 12299 10659
rect 13001 10625 13035 10659
rect 13553 10625 13587 10659
rect 14473 10625 14507 10659
rect 14657 10625 14691 10659
rect 16129 10625 16163 10659
rect 17233 10625 17267 10659
rect 18889 10625 18923 10659
rect 21281 10625 21315 10659
rect 21925 10625 21959 10659
rect 23673 10625 23707 10659
rect 1409 10557 1443 10591
rect 1676 10557 1710 10591
rect 11345 10557 11379 10591
rect 15209 10557 15243 10591
rect 16037 10557 16071 10591
rect 19156 10557 19190 10591
rect 23940 10557 23974 10591
rect 11897 10489 11931 10523
rect 12817 10489 12851 10523
rect 20913 10489 20947 10523
rect 21833 10489 21867 10523
rect 2789 10421 2823 10455
rect 12909 10421 12943 10455
rect 13829 10421 13863 10455
rect 14381 10421 14415 10455
rect 15485 10421 15519 10455
rect 15945 10421 15979 10455
rect 20269 10421 20303 10455
rect 21741 10421 21775 10455
rect 25053 10421 25087 10455
rect 25605 10421 25639 10455
rect 1685 10217 1719 10251
rect 11621 10217 11655 10251
rect 13185 10217 13219 10251
rect 15301 10217 15335 10251
rect 16313 10217 16347 10251
rect 16681 10217 16715 10251
rect 18429 10217 18463 10251
rect 21281 10217 21315 10251
rect 22477 10217 22511 10251
rect 13553 10149 13587 10183
rect 23734 10149 23768 10183
rect 11989 10081 12023 10115
rect 14013 10081 14047 10115
rect 15669 10081 15703 10115
rect 17233 10081 17267 10115
rect 18797 10081 18831 10115
rect 18889 10081 18923 10115
rect 12081 10013 12115 10047
rect 12173 10013 12207 10047
rect 14105 10013 14139 10047
rect 14197 10013 14231 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 18981 10013 19015 10047
rect 21373 10013 21407 10047
rect 21465 10013 21499 10047
rect 23489 10013 23523 10047
rect 20913 9945 20947 9979
rect 21925 9945 21959 9979
rect 11161 9877 11195 9911
rect 11437 9877 11471 9911
rect 12633 9877 12667 9911
rect 13645 9877 13679 9911
rect 14841 9877 14875 9911
rect 16865 9877 16899 9911
rect 18153 9877 18187 9911
rect 24869 9877 24903 9911
rect 25421 9877 25455 9911
rect 14013 9673 14047 9707
rect 16129 9673 16163 9707
rect 20729 9673 20763 9707
rect 21741 9673 21775 9707
rect 22109 9673 22143 9707
rect 23397 9673 23431 9707
rect 23949 9673 23983 9707
rect 17417 9605 17451 9639
rect 18061 9605 18095 9639
rect 21649 9605 21683 9639
rect 13001 9537 13035 9571
rect 14749 9537 14783 9571
rect 16773 9537 16807 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 19441 9537 19475 9571
rect 21373 9537 21407 9571
rect 9873 9469 9907 9503
rect 10129 9469 10163 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 21097 9469 21131 9503
rect 15016 9401 15050 9435
rect 17877 9401 17911 9435
rect 20269 9401 20303 9435
rect 21189 9401 21223 9435
rect 22477 9537 22511 9571
rect 24133 9537 24167 9571
rect 24400 9469 24434 9503
rect 9689 9333 9723 9367
rect 11253 9333 11287 9367
rect 11805 9333 11839 9367
rect 12173 9333 12207 9367
rect 12449 9333 12483 9367
rect 13737 9333 13771 9367
rect 14657 9333 14691 9367
rect 17049 9333 17083 9367
rect 18429 9333 18463 9367
rect 19165 9333 19199 9367
rect 21649 9333 21683 9367
rect 23029 9333 23063 9367
rect 25513 9333 25547 9367
rect 9965 9129 9999 9163
rect 12541 9129 12575 9163
rect 13645 9129 13679 9163
rect 14105 9129 14139 9163
rect 17785 9129 17819 9163
rect 18245 9129 18279 9163
rect 19993 9129 20027 9163
rect 20729 9129 20763 9163
rect 21557 9129 21591 9163
rect 22661 9129 22695 9163
rect 23029 9129 23063 9163
rect 23673 9129 23707 9163
rect 24225 9129 24259 9163
rect 11069 9061 11103 9095
rect 13461 9061 13495 9095
rect 14749 9061 14783 9095
rect 15568 9061 15602 9095
rect 17601 9061 17635 9095
rect 24133 9061 24167 9095
rect 11417 8993 11451 9027
rect 14013 8993 14047 9027
rect 15301 8993 15335 9027
rect 18153 8993 18187 9027
rect 19441 8993 19475 9027
rect 21465 8993 21499 9027
rect 24593 8993 24627 9027
rect 11161 8925 11195 8959
rect 14197 8925 14231 8959
rect 18337 8925 18371 8959
rect 21741 8925 21775 8959
rect 22569 8925 22603 8959
rect 23121 8925 23155 8959
rect 23305 8925 23339 8959
rect 24685 8925 24719 8959
rect 24777 8925 24811 8959
rect 17233 8857 17267 8891
rect 19625 8857 19659 8891
rect 21097 8857 21131 8891
rect 25237 8857 25271 8891
rect 16681 8789 16715 8823
rect 18797 8789 18831 8823
rect 22201 8789 22235 8823
rect 10885 8585 10919 8619
rect 11161 8585 11195 8619
rect 12081 8585 12115 8619
rect 12173 8585 12207 8619
rect 14381 8585 14415 8619
rect 14749 8585 14783 8619
rect 17049 8585 17083 8619
rect 17509 8585 17543 8619
rect 21373 8585 21407 8619
rect 22385 8585 22419 8619
rect 23029 8585 23063 8619
rect 23489 8585 23523 8619
rect 25513 8585 25547 8619
rect 11345 8449 11379 8483
rect 11897 8449 11931 8483
rect 21925 8517 21959 8551
rect 22661 8517 22695 8551
rect 14933 8449 14967 8483
rect 18705 8449 18739 8483
rect 24133 8449 24167 8483
rect 12081 8381 12115 8415
rect 12449 8381 12483 8415
rect 12705 8381 12739 8415
rect 17785 8381 17819 8415
rect 18521 8381 18555 8415
rect 19993 8381 20027 8415
rect 20260 8381 20294 8415
rect 22477 8381 22511 8415
rect 24041 8381 24075 8415
rect 15200 8313 15234 8347
rect 18429 8313 18463 8347
rect 19073 8313 19107 8347
rect 19441 8313 19475 8347
rect 19901 8313 19935 8347
rect 24400 8313 24434 8347
rect 13829 8245 13863 8279
rect 16313 8245 16347 8279
rect 18061 8245 18095 8279
rect 12081 8041 12115 8075
rect 13553 8041 13587 8075
rect 14013 8041 14047 8075
rect 14933 8041 14967 8075
rect 15301 8041 15335 8075
rect 17785 8041 17819 8075
rect 18153 8041 18187 8075
rect 21097 8041 21131 8075
rect 24593 8041 24627 8075
rect 24961 8041 24995 8075
rect 11989 7973 12023 8007
rect 12449 7973 12483 8007
rect 14105 7973 14139 8007
rect 15853 7973 15887 8007
rect 13185 7905 13219 7939
rect 16957 7905 16991 7939
rect 18521 7905 18555 7939
rect 21465 7905 21499 7939
rect 22661 7905 22695 7939
rect 22928 7905 22962 7939
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 14289 7837 14323 7871
rect 17049 7837 17083 7871
rect 17233 7837 17267 7871
rect 18613 7837 18647 7871
rect 18705 7837 18739 7871
rect 19717 7837 19751 7871
rect 21557 7837 21591 7871
rect 21741 7837 21775 7871
rect 16129 7769 16163 7803
rect 16589 7769 16623 7803
rect 20729 7769 20763 7803
rect 22477 7769 22511 7803
rect 13645 7701 13679 7735
rect 19441 7701 19475 7735
rect 22201 7701 22235 7735
rect 24041 7701 24075 7735
rect 11529 7497 11563 7531
rect 15025 7497 15059 7531
rect 17417 7497 17451 7531
rect 17785 7497 17819 7531
rect 18521 7497 18555 7531
rect 18889 7497 18923 7531
rect 19349 7497 19383 7531
rect 21833 7497 21867 7531
rect 23121 7497 23155 7531
rect 11897 7429 11931 7463
rect 16037 7429 16071 7463
rect 23673 7429 23707 7463
rect 13001 7361 13035 7395
rect 14565 7361 14599 7395
rect 16589 7361 16623 7395
rect 19441 7361 19475 7395
rect 22477 7361 22511 7395
rect 22661 7361 22695 7395
rect 24317 7361 24351 7395
rect 25053 7361 25087 7395
rect 12909 7293 12943 7327
rect 13921 7293 13955 7327
rect 14381 7293 14415 7327
rect 14473 7293 14507 7327
rect 22385 7293 22419 7327
rect 12265 7225 12299 7259
rect 12817 7225 12851 7259
rect 13553 7225 13587 7259
rect 15577 7225 15611 7259
rect 19686 7225 19720 7259
rect 24041 7225 24075 7259
rect 24777 7225 24811 7259
rect 25237 7225 25271 7259
rect 12449 7157 12483 7191
rect 14013 7157 14047 7191
rect 15853 7157 15887 7191
rect 16405 7157 16439 7191
rect 16497 7157 16531 7191
rect 17141 7157 17175 7191
rect 18061 7157 18095 7191
rect 20821 7157 20855 7191
rect 21465 7157 21499 7191
rect 22017 7157 22051 7191
rect 23489 7157 23523 7191
rect 24133 7157 24167 7191
rect 12449 6953 12483 6987
rect 12909 6953 12943 6987
rect 14657 6953 14691 6987
rect 15669 6953 15703 6987
rect 16497 6953 16531 6987
rect 18889 6953 18923 6987
rect 22661 6953 22695 6987
rect 24133 6953 24167 6987
rect 13645 6885 13679 6919
rect 17325 6885 17359 6919
rect 21557 6885 21591 6919
rect 23020 6885 23054 6919
rect 12173 6817 12207 6851
rect 15117 6817 15151 6851
rect 15761 6817 15795 6851
rect 17417 6817 17451 6851
rect 18981 6817 19015 6851
rect 22293 6817 22327 6851
rect 22753 6817 22787 6851
rect 25237 6817 25271 6851
rect 13737 6749 13771 6783
rect 13829 6749 13863 6783
rect 15945 6749 15979 6783
rect 17601 6749 17635 6783
rect 19165 6749 19199 6783
rect 19993 6749 20027 6783
rect 21649 6749 21683 6783
rect 21833 6749 21867 6783
rect 15301 6681 15335 6715
rect 16865 6681 16899 6715
rect 18521 6681 18555 6715
rect 21189 6681 21223 6715
rect 13277 6613 13311 6647
rect 14381 6613 14415 6647
rect 16957 6613 16991 6647
rect 18153 6613 18187 6647
rect 19717 6613 19751 6647
rect 20729 6613 20763 6647
rect 25421 6613 25455 6647
rect 14565 6409 14599 6443
rect 19073 6409 19107 6443
rect 19441 6409 19475 6443
rect 21925 6409 21959 6443
rect 22753 6409 22787 6443
rect 24041 6409 24075 6443
rect 25237 6409 25271 6443
rect 15025 6341 15059 6375
rect 21649 6341 21683 6375
rect 11897 6273 11931 6307
rect 13737 6273 13771 6307
rect 14197 6273 14231 6307
rect 15485 6273 15519 6307
rect 18705 6273 18739 6307
rect 19625 6273 19659 6307
rect 24777 6273 24811 6307
rect 17877 6205 17911 6239
rect 18429 6205 18463 6239
rect 19881 6205 19915 6239
rect 22109 6205 22143 6239
rect 13001 6137 13035 6171
rect 13553 6137 13587 6171
rect 13645 6137 13679 6171
rect 15752 6137 15786 6171
rect 23489 6137 23523 6171
rect 24593 6137 24627 6171
rect 12265 6069 12299 6103
rect 12633 6069 12667 6103
rect 13185 6069 13219 6103
rect 15393 6069 15427 6103
rect 16865 6069 16899 6103
rect 17509 6069 17543 6103
rect 18061 6069 18095 6103
rect 18521 6069 18555 6103
rect 21005 6069 21039 6103
rect 22293 6069 22327 6103
rect 24225 6069 24259 6103
rect 24685 6069 24719 6103
rect 14197 5865 14231 5899
rect 15301 5865 15335 5899
rect 16405 5865 16439 5899
rect 18429 5865 18463 5899
rect 18981 5865 19015 5899
rect 19441 5865 19475 5899
rect 21373 5865 21407 5899
rect 22017 5865 22051 5899
rect 25145 5865 25179 5899
rect 12081 5797 12115 5831
rect 15669 5797 15703 5831
rect 17316 5797 17350 5831
rect 21281 5797 21315 5831
rect 12440 5729 12474 5763
rect 15761 5729 15795 5763
rect 17049 5729 17083 5763
rect 19717 5729 19751 5763
rect 22477 5729 22511 5763
rect 23949 5729 23983 5763
rect 12173 5661 12207 5695
rect 15945 5661 15979 5695
rect 21465 5661 21499 5695
rect 24041 5661 24075 5695
rect 24225 5661 24259 5695
rect 15117 5593 15151 5627
rect 19901 5593 19935 5627
rect 22385 5593 22419 5627
rect 23581 5593 23615 5627
rect 24961 5593 24995 5627
rect 13553 5525 13587 5559
rect 16957 5525 16991 5559
rect 20361 5525 20395 5559
rect 20913 5525 20947 5559
rect 22661 5525 22695 5559
rect 23121 5525 23155 5559
rect 23489 5525 23523 5559
rect 24685 5525 24719 5559
rect 15945 5321 15979 5355
rect 19533 5321 19567 5355
rect 19901 5321 19935 5355
rect 21005 5321 21039 5355
rect 21373 5321 21407 5355
rect 22017 5321 22051 5355
rect 23029 5321 23063 5355
rect 25697 5321 25731 5355
rect 11897 5253 11931 5287
rect 23397 5253 23431 5287
rect 25145 5253 25179 5287
rect 11345 5185 11379 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 18981 5185 19015 5219
rect 20545 5185 20579 5219
rect 22477 5185 22511 5219
rect 22661 5185 22695 5219
rect 22845 5185 22879 5219
rect 23765 5185 23799 5219
rect 12817 5117 12851 5151
rect 13921 5117 13955 5151
rect 14013 5117 14047 5151
rect 16773 5117 16807 5151
rect 17325 5117 17359 5151
rect 18337 5117 18371 5151
rect 18797 5117 18831 5151
rect 20453 5117 20487 5151
rect 22385 5117 22419 5151
rect 13553 5049 13587 5083
rect 14258 5049 14292 5083
rect 18889 5049 18923 5083
rect 21925 5049 21959 5083
rect 22845 5049 22879 5083
rect 24032 5049 24066 5083
rect 12173 4981 12207 5015
rect 12449 4981 12483 5015
rect 15393 4981 15427 5015
rect 16405 4981 16439 5015
rect 16957 4981 16991 5015
rect 17785 4981 17819 5015
rect 18429 4981 18463 5015
rect 19993 4981 20027 5015
rect 20361 4981 20395 5015
rect 11805 4777 11839 4811
rect 13645 4777 13679 4811
rect 16129 4777 16163 4811
rect 16681 4777 16715 4811
rect 17049 4777 17083 4811
rect 18153 4777 18187 4811
rect 18797 4777 18831 4811
rect 19257 4777 19291 4811
rect 20729 4777 20763 4811
rect 22937 4777 22971 4811
rect 12173 4709 12207 4743
rect 17141 4709 17175 4743
rect 18245 4709 18279 4743
rect 20269 4709 20303 4743
rect 21158 4709 21192 4743
rect 12532 4641 12566 4675
rect 15577 4641 15611 4675
rect 16589 4641 16623 4675
rect 19625 4641 19659 4675
rect 23653 4641 23687 4675
rect 12265 4573 12299 4607
rect 17325 4573 17359 4607
rect 19717 4573 19751 4607
rect 19901 4573 19935 4607
rect 20913 4573 20947 4607
rect 23397 4573 23431 4607
rect 19165 4505 19199 4539
rect 23213 4505 23247 4539
rect 14749 4437 14783 4471
rect 15025 4437 15059 4471
rect 15761 4437 15795 4471
rect 17693 4437 17727 4471
rect 22293 4437 22327 4471
rect 24777 4437 24811 4471
rect 12265 4233 12299 4267
rect 17233 4233 17267 4267
rect 21005 4233 21039 4267
rect 21925 4233 21959 4267
rect 23029 4233 23063 4267
rect 23397 4233 23431 4267
rect 25053 4233 25087 4267
rect 16589 4097 16623 4131
rect 16773 4097 16807 4131
rect 18521 4097 18555 4131
rect 18705 4097 18739 4131
rect 19165 4097 19199 4131
rect 23673 4097 23707 4131
rect 11345 4029 11379 4063
rect 11897 4029 11931 4063
rect 13369 4029 13403 4063
rect 13636 4029 13670 4063
rect 15669 4029 15703 4063
rect 18429 4029 18463 4063
rect 19349 4029 19383 4063
rect 19625 4029 19659 4063
rect 21557 4029 21591 4063
rect 22109 4029 22143 4063
rect 22661 4029 22695 4063
rect 16497 3961 16531 3995
rect 19870 3961 19904 3995
rect 23918 3961 23952 3995
rect 11529 3893 11563 3927
rect 12725 3893 12759 3927
rect 13277 3893 13311 3927
rect 14749 3893 14783 3927
rect 15945 3893 15979 3927
rect 16129 3893 16163 3927
rect 17785 3893 17819 3927
rect 18061 3893 18095 3927
rect 19349 3893 19383 3927
rect 19441 3893 19475 3927
rect 22293 3893 22327 3927
rect 11713 3689 11747 3723
rect 13461 3689 13495 3723
rect 14657 3689 14691 3723
rect 15117 3689 15151 3723
rect 19349 3689 19383 3723
rect 20361 3689 20395 3723
rect 20913 3689 20947 3723
rect 21373 3689 21407 3723
rect 22109 3689 22143 3723
rect 22569 3689 22603 3723
rect 23305 3689 23339 3723
rect 23765 3689 23799 3723
rect 24869 3689 24903 3723
rect 25237 3689 25271 3723
rect 25329 3689 25363 3723
rect 14013 3621 14047 3655
rect 16221 3621 16255 3655
rect 16764 3621 16798 3655
rect 20085 3621 20119 3655
rect 23673 3621 23707 3655
rect 10517 3553 10551 3587
rect 11529 3553 11563 3587
rect 12541 3553 12575 3587
rect 15393 3553 15427 3587
rect 21281 3553 21315 3587
rect 14105 3485 14139 3519
rect 14289 3485 14323 3519
rect 16497 3485 16531 3519
rect 19441 3485 19475 3519
rect 19533 3485 19567 3519
rect 21465 3485 21499 3519
rect 23949 3485 23983 3519
rect 25513 3485 25547 3519
rect 18889 3417 18923 3451
rect 24409 3417 24443 3451
rect 10701 3349 10735 3383
rect 12725 3349 12759 3383
rect 13645 3349 13679 3383
rect 15577 3349 15611 3383
rect 17877 3349 17911 3383
rect 18429 3349 18463 3383
rect 18981 3349 19015 3383
rect 10793 3145 10827 3179
rect 11161 3145 11195 3179
rect 12265 3145 12299 3179
rect 12909 3145 12943 3179
rect 13369 3145 13403 3179
rect 14381 3145 14415 3179
rect 15945 3145 15979 3179
rect 17325 3145 17359 3179
rect 19717 3145 19751 3179
rect 20269 3145 20303 3179
rect 20821 3145 20855 3179
rect 22201 3145 22235 3179
rect 23305 3145 23339 3179
rect 23857 3145 23891 3179
rect 25237 3145 25271 3179
rect 25881 3145 25915 3179
rect 10425 3077 10459 3111
rect 14105 3077 14139 3111
rect 20729 3077 20763 3111
rect 21833 3077 21867 3111
rect 24409 3077 24443 3111
rect 12449 3009 12483 3043
rect 14565 3009 14599 3043
rect 21373 3009 21407 3043
rect 25513 3009 25547 3043
rect 10241 2941 10275 2975
rect 11253 2941 11287 2975
rect 11805 2941 11839 2975
rect 13461 2941 13495 2975
rect 14832 2941 14866 2975
rect 18337 2941 18371 2975
rect 18593 2941 18627 2975
rect 21189 2941 21223 2975
rect 22477 2941 22511 2975
rect 24593 2941 24627 2975
rect 16497 2873 16531 2907
rect 17785 2873 17819 2907
rect 21281 2873 21315 2907
rect 11437 2805 11471 2839
rect 13645 2805 13679 2839
rect 16957 2805 16991 2839
rect 22661 2805 22695 2839
rect 24777 2805 24811 2839
rect 5733 2601 5767 2635
rect 8309 2601 8343 2635
rect 13829 2601 13863 2635
rect 14197 2601 14231 2635
rect 15669 2601 15703 2635
rect 17693 2601 17727 2635
rect 18153 2601 18187 2635
rect 19809 2601 19843 2635
rect 20913 2601 20947 2635
rect 21373 2601 21407 2635
rect 23857 2601 23891 2635
rect 12449 2533 12483 2567
rect 2789 2465 2823 2499
rect 3341 2465 3375 2499
rect 5549 2465 5583 2499
rect 6101 2465 6135 2499
rect 8125 2465 8159 2499
rect 10333 2465 10367 2499
rect 10885 2465 10919 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 13185 2465 13219 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 16313 2465 16347 2499
rect 17049 2465 17083 2499
rect 18705 2465 18739 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 21741 2465 21775 2499
rect 22293 2465 22327 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 13093 2397 13127 2431
rect 16405 2397 16439 2431
rect 16497 2397 16531 2431
rect 18797 2397 18831 2431
rect 18889 2397 18923 2431
rect 2973 2329 3007 2363
rect 15945 2329 15979 2363
rect 18337 2329 18371 2363
rect 23029 2329 23063 2363
rect 24777 2329 24811 2363
rect 8677 2261 8711 2295
rect 10517 2261 10551 2295
rect 11621 2261 11655 2295
rect 13369 2261 13403 2295
rect 14473 2261 14507 2295
rect 15301 2261 15335 2295
rect 17325 2261 17359 2295
rect 19349 2261 19383 2295
rect 20085 2261 20119 2295
rect 21925 2261 21959 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 15930 25480 15936 25492
rect 14507 25452 15936 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 15930 25440 15936 25452
rect 15988 25440 15994 25492
rect 16853 25483 16911 25489
rect 16853 25449 16865 25483
rect 16899 25480 16911 25483
rect 17954 25480 17960 25492
rect 16899 25452 17960 25480
rect 16899 25449 16911 25452
rect 16853 25443 16911 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 19613 25483 19671 25489
rect 19613 25449 19625 25483
rect 19659 25480 19671 25483
rect 20070 25480 20076 25492
rect 19659 25452 20076 25480
rect 19659 25449 19671 25452
rect 19613 25443 19671 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 22189 25483 22247 25489
rect 22189 25449 22201 25483
rect 22235 25480 22247 25483
rect 22738 25480 22744 25492
rect 22235 25452 22744 25480
rect 22235 25449 22247 25452
rect 22189 25443 22247 25449
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 14277 25347 14335 25353
rect 14277 25313 14289 25347
rect 14323 25344 14335 25347
rect 14366 25344 14372 25356
rect 14323 25316 14372 25344
rect 14323 25313 14335 25316
rect 14277 25307 14335 25313
rect 14366 25304 14372 25316
rect 14424 25304 14430 25356
rect 15565 25347 15623 25353
rect 15565 25313 15577 25347
rect 15611 25313 15623 25347
rect 15565 25307 15623 25313
rect 16669 25347 16727 25353
rect 16669 25313 16681 25347
rect 16715 25344 16727 25347
rect 16942 25344 16948 25356
rect 16715 25316 16948 25344
rect 16715 25313 16727 25316
rect 16669 25307 16727 25313
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25276 15347 25279
rect 15580 25276 15608 25307
rect 16942 25304 16948 25316
rect 17000 25304 17006 25356
rect 19426 25344 19432 25356
rect 19387 25316 19432 25344
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 22002 25344 22008 25356
rect 21963 25316 22008 25344
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 17586 25276 17592 25288
rect 15335 25248 17592 25276
rect 15335 25245 15347 25248
rect 15289 25239 15347 25245
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 15749 25211 15807 25217
rect 15749 25177 15761 25211
rect 15795 25208 15807 25211
rect 17310 25208 17316 25220
rect 15795 25180 17316 25208
rect 15795 25177 15807 25180
rect 15749 25171 15807 25177
rect 17310 25168 17316 25180
rect 17368 25168 17374 25220
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16390 25140 16396 25152
rect 16255 25112 16396 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 16390 25100 16396 25112
rect 16448 25100 16454 25152
rect 18138 25140 18144 25152
rect 18099 25112 18144 25140
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 21634 25100 21640 25152
rect 21692 25140 21698 25152
rect 24670 25140 24676 25152
rect 21692 25112 24676 25140
rect 21692 25100 21698 25112
rect 24670 25100 24676 25112
rect 24728 25100 24734 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 18966 24896 18972 24948
rect 19024 24936 19030 24948
rect 23566 24936 23572 24948
rect 19024 24908 23572 24936
rect 19024 24896 19030 24908
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 16390 24868 16396 24880
rect 16040 24840 16396 24868
rect 16040 24809 16068 24840
rect 16390 24828 16396 24840
rect 16448 24868 16454 24880
rect 21726 24868 21732 24880
rect 16448 24840 21732 24868
rect 16448 24828 16454 24840
rect 17512 24809 17540 24840
rect 18708 24809 18736 24840
rect 21726 24828 21732 24840
rect 21784 24828 21790 24880
rect 22002 24868 22008 24880
rect 21963 24840 22008 24868
rect 22002 24828 22008 24840
rect 22060 24828 22066 24880
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24769 16083 24803
rect 16025 24763 16083 24769
rect 17497 24803 17555 24809
rect 17497 24769 17509 24803
rect 17543 24769 17555 24803
rect 17497 24763 17555 24769
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24769 18751 24803
rect 18693 24763 18751 24769
rect 19518 24760 19524 24812
rect 19576 24760 19582 24812
rect 12894 24692 12900 24744
rect 12952 24732 12958 24744
rect 13173 24735 13231 24741
rect 13173 24732 13185 24735
rect 12952 24704 13185 24732
rect 12952 24692 12958 24704
rect 13173 24701 13185 24704
rect 13219 24732 13231 24735
rect 13725 24735 13783 24741
rect 13725 24732 13737 24735
rect 13219 24704 13737 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 13725 24701 13737 24704
rect 13771 24701 13783 24735
rect 14274 24732 14280 24744
rect 14235 24704 14280 24732
rect 13725 24695 13783 24701
rect 14274 24692 14280 24704
rect 14332 24732 14338 24744
rect 14829 24735 14887 24741
rect 14829 24732 14841 24735
rect 14332 24704 14841 24732
rect 14332 24692 14338 24704
rect 14829 24701 14841 24704
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 16945 24735 17003 24741
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 18138 24732 18144 24744
rect 16991 24704 18144 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 18138 24692 18144 24704
rect 18196 24732 18202 24744
rect 18417 24735 18475 24741
rect 18417 24732 18429 24735
rect 18196 24704 18429 24732
rect 18196 24692 18202 24704
rect 18417 24701 18429 24704
rect 18463 24701 18475 24735
rect 19536 24732 19564 24760
rect 19889 24735 19947 24741
rect 19889 24732 19901 24735
rect 19536 24704 19901 24732
rect 18417 24695 18475 24701
rect 19889 24701 19901 24704
rect 19935 24732 19947 24735
rect 20441 24735 20499 24741
rect 20441 24732 20453 24735
rect 19935 24704 20453 24732
rect 19935 24701 19947 24704
rect 19889 24695 19947 24701
rect 20441 24701 20453 24704
rect 20487 24701 20499 24735
rect 20441 24695 20499 24701
rect 20993 24735 21051 24741
rect 20993 24701 21005 24735
rect 21039 24732 21051 24735
rect 21361 24735 21419 24741
rect 21361 24732 21373 24735
rect 21039 24704 21373 24732
rect 21039 24701 21051 24704
rect 20993 24695 21051 24701
rect 21361 24701 21373 24704
rect 21407 24701 21419 24735
rect 21361 24695 21419 24701
rect 21542 24692 21548 24744
rect 21600 24732 21606 24744
rect 22189 24735 22247 24741
rect 22189 24732 22201 24735
rect 21600 24704 22201 24732
rect 21600 24692 21606 24704
rect 22189 24701 22201 24704
rect 22235 24732 22247 24735
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 22235 24704 22753 24732
rect 22235 24701 22247 24704
rect 22189 24695 22247 24701
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 14185 24667 14243 24673
rect 14185 24633 14197 24667
rect 14231 24664 14243 24667
rect 14366 24664 14372 24676
rect 14231 24636 14372 24664
rect 14231 24633 14243 24636
rect 14185 24627 14243 24633
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 15194 24664 15200 24676
rect 15155 24636 15200 24664
rect 15194 24624 15200 24636
rect 15252 24664 15258 24676
rect 15841 24667 15899 24673
rect 15841 24664 15853 24667
rect 15252 24636 15853 24664
rect 15252 24624 15258 24636
rect 15841 24633 15853 24636
rect 15887 24633 15899 24667
rect 15841 24627 15899 24633
rect 17494 24624 17500 24676
rect 17552 24664 17558 24676
rect 17865 24667 17923 24673
rect 17865 24664 17877 24667
rect 17552 24636 17877 24664
rect 17552 24624 17558 24636
rect 17865 24633 17877 24636
rect 17911 24664 17923 24667
rect 18509 24667 18567 24673
rect 18509 24664 18521 24667
rect 17911 24636 18521 24664
rect 17911 24633 17923 24636
rect 17865 24627 17923 24633
rect 18509 24633 18521 24636
rect 18555 24633 18567 24667
rect 18509 24627 18567 24633
rect 19426 24624 19432 24676
rect 19484 24664 19490 24676
rect 19521 24667 19579 24673
rect 19521 24664 19533 24667
rect 19484 24636 19533 24664
rect 19484 24624 19490 24636
rect 19521 24633 19533 24636
rect 19567 24664 19579 24667
rect 20162 24664 20168 24676
rect 19567 24636 20168 24664
rect 19567 24633 19579 24636
rect 19521 24627 19579 24633
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 22094 24664 22100 24676
rect 21192 24636 22100 24664
rect 13354 24596 13360 24608
rect 13315 24568 13360 24596
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 14458 24596 14464 24608
rect 14419 24568 14464 24596
rect 14458 24556 14464 24568
rect 14516 24556 14522 24608
rect 15378 24596 15384 24608
rect 15339 24568 15384 24596
rect 15378 24556 15384 24568
rect 15436 24556 15442 24608
rect 15746 24596 15752 24608
rect 15707 24568 15752 24596
rect 15746 24556 15752 24568
rect 15804 24556 15810 24608
rect 16761 24599 16819 24605
rect 16761 24565 16773 24599
rect 16807 24596 16819 24599
rect 16942 24596 16948 24608
rect 16807 24568 16948 24596
rect 16807 24565 16819 24568
rect 16761 24559 16819 24565
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 18049 24599 18107 24605
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18138 24596 18144 24608
rect 18095 24568 18144 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 20070 24596 20076 24608
rect 20031 24568 20076 24596
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 21192 24605 21220 24636
rect 22094 24624 22100 24636
rect 22152 24624 22158 24676
rect 21177 24599 21235 24605
rect 21177 24565 21189 24599
rect 21223 24565 21235 24599
rect 21177 24559 21235 24565
rect 21361 24599 21419 24605
rect 21361 24565 21373 24599
rect 21407 24596 21419 24599
rect 21637 24599 21695 24605
rect 21637 24596 21649 24599
rect 21407 24568 21649 24596
rect 21407 24565 21419 24568
rect 21361 24559 21419 24565
rect 21637 24565 21649 24568
rect 21683 24596 21695 24599
rect 21818 24596 21824 24608
rect 21683 24568 21824 24596
rect 21683 24565 21695 24568
rect 21637 24559 21695 24565
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22370 24596 22376 24608
rect 22331 24568 22376 24596
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 23658 24596 23664 24608
rect 23619 24568 23664 24596
rect 23658 24556 23664 24568
rect 23716 24556 23722 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 15378 24352 15384 24404
rect 15436 24392 15442 24404
rect 16298 24392 16304 24404
rect 15436 24364 16304 24392
rect 15436 24352 15442 24364
rect 16298 24352 16304 24364
rect 16356 24352 16362 24404
rect 19797 24395 19855 24401
rect 19797 24361 19809 24395
rect 19843 24392 19855 24395
rect 20622 24392 20628 24404
rect 19843 24364 20628 24392
rect 19843 24361 19855 24364
rect 19797 24355 19855 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 21450 24392 21456 24404
rect 21411 24364 21456 24392
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 21910 24392 21916 24404
rect 21871 24364 21916 24392
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 22554 24392 22560 24404
rect 22515 24364 22560 24392
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 23661 24395 23719 24401
rect 23661 24361 23673 24395
rect 23707 24392 23719 24395
rect 23750 24392 23756 24404
rect 23707 24364 23756 24392
rect 23707 24361 23719 24364
rect 23661 24355 23719 24361
rect 23750 24352 23756 24364
rect 23808 24352 23814 24404
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 10134 24284 10140 24336
rect 10192 24324 10198 24336
rect 15473 24327 15531 24333
rect 15473 24324 15485 24327
rect 10192 24296 15485 24324
rect 10192 24284 10198 24296
rect 15473 24293 15485 24296
rect 15519 24324 15531 24327
rect 15562 24324 15568 24336
rect 15519 24296 15568 24324
rect 15519 24293 15531 24296
rect 15473 24287 15531 24293
rect 15562 24284 15568 24296
rect 15620 24324 15626 24336
rect 15746 24324 15752 24336
rect 15620 24296 15752 24324
rect 15620 24284 15626 24296
rect 15746 24284 15752 24296
rect 15804 24284 15810 24336
rect 12066 24216 12072 24268
rect 12124 24256 12130 24268
rect 12161 24259 12219 24265
rect 12161 24256 12173 24259
rect 12124 24228 12173 24256
rect 12124 24216 12130 24228
rect 12161 24225 12173 24228
rect 12207 24225 12219 24259
rect 12161 24219 12219 24225
rect 13265 24259 13323 24265
rect 13265 24225 13277 24259
rect 13311 24256 13323 24259
rect 13722 24256 13728 24268
rect 13311 24228 13728 24256
rect 13311 24225 13323 24228
rect 13265 24219 13323 24225
rect 13722 24216 13728 24228
rect 13780 24216 13786 24268
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 16666 24256 16672 24268
rect 16255 24228 16672 24256
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 17681 24259 17739 24265
rect 17681 24225 17693 24259
rect 17727 24256 17739 24259
rect 18046 24256 18052 24268
rect 17727 24228 18052 24256
rect 17727 24225 17739 24228
rect 17681 24219 17739 24225
rect 18046 24216 18052 24228
rect 18104 24256 18110 24268
rect 18141 24259 18199 24265
rect 18141 24256 18153 24259
rect 18104 24228 18153 24256
rect 18104 24216 18110 24228
rect 18141 24225 18153 24228
rect 18187 24225 18199 24259
rect 18141 24219 18199 24225
rect 18322 24216 18328 24268
rect 18380 24256 18386 24268
rect 19613 24259 19671 24265
rect 19613 24256 19625 24259
rect 18380 24228 19625 24256
rect 18380 24216 18386 24228
rect 19613 24225 19625 24228
rect 19659 24225 19671 24259
rect 19613 24219 19671 24225
rect 21082 24216 21088 24268
rect 21140 24256 21146 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 21140 24228 21281 24256
rect 21140 24216 21146 24228
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 22370 24256 22376 24268
rect 22331 24228 22376 24256
rect 21269 24219 21327 24225
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 23106 24216 23112 24268
rect 23164 24256 23170 24268
rect 23477 24259 23535 24265
rect 23477 24256 23489 24259
rect 23164 24228 23489 24256
rect 23164 24216 23170 24228
rect 23477 24225 23489 24228
rect 23523 24225 23535 24259
rect 23477 24219 23535 24225
rect 24210 24216 24216 24268
rect 24268 24256 24274 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24268 24228 24593 24256
rect 24268 24216 24274 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 11790 24148 11796 24200
rect 11848 24188 11854 24200
rect 12253 24191 12311 24197
rect 12253 24188 12265 24191
rect 11848 24160 12265 24188
rect 11848 24148 11854 24160
rect 12253 24157 12265 24160
rect 12299 24157 12311 24191
rect 12253 24151 12311 24157
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24188 12495 24191
rect 12710 24188 12716 24200
rect 12483 24160 12716 24188
rect 12483 24157 12495 24160
rect 12437 24151 12495 24157
rect 12710 24148 12716 24160
rect 12768 24188 12774 24200
rect 12768 24160 12940 24188
rect 12768 24148 12774 24160
rect 12912 24129 12940 24160
rect 13630 24148 13636 24200
rect 13688 24188 13694 24200
rect 13817 24191 13875 24197
rect 13817 24188 13829 24191
rect 13688 24160 13829 24188
rect 13688 24148 13694 24160
rect 13817 24157 13829 24160
rect 13863 24157 13875 24191
rect 13998 24188 14004 24200
rect 13959 24160 14004 24188
rect 13817 24151 13875 24157
rect 13998 24148 14004 24160
rect 14056 24148 14062 24200
rect 16114 24148 16120 24200
rect 16172 24188 16178 24200
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 16172 24160 16405 24188
rect 16172 24148 16178 24160
rect 16393 24157 16405 24160
rect 16439 24188 16451 24191
rect 16482 24188 16488 24200
rect 16439 24160 16488 24188
rect 16439 24157 16451 24160
rect 16393 24151 16451 24157
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18414 24188 18420 24200
rect 18375 24160 18420 24188
rect 18233 24151 18291 24157
rect 12897 24123 12955 24129
rect 12897 24089 12909 24123
rect 12943 24120 12955 24123
rect 15841 24123 15899 24129
rect 12943 24092 15056 24120
rect 12943 24089 12955 24092
rect 12897 24083 12955 24089
rect 11330 24052 11336 24064
rect 11291 24024 11336 24052
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 11793 24055 11851 24061
rect 11793 24021 11805 24055
rect 11839 24052 11851 24055
rect 12342 24052 12348 24064
rect 11839 24024 12348 24052
rect 11839 24021 11851 24024
rect 11793 24015 11851 24021
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 13354 24052 13360 24064
rect 13315 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 15028 24061 15056 24092
rect 15841 24089 15853 24123
rect 15887 24120 15899 24123
rect 17678 24120 17684 24132
rect 15887 24092 17684 24120
rect 15887 24089 15899 24092
rect 15841 24083 15899 24089
rect 17678 24080 17684 24092
rect 17736 24120 17742 24132
rect 18248 24120 18276 24151
rect 18414 24148 18420 24160
rect 18472 24148 18478 24200
rect 17736 24092 18276 24120
rect 17736 24080 17742 24092
rect 15013 24055 15071 24061
rect 15013 24021 15025 24055
rect 15059 24052 15071 24055
rect 15746 24052 15752 24064
rect 15059 24024 15752 24052
rect 15059 24021 15071 24024
rect 15013 24015 15071 24021
rect 15746 24012 15752 24024
rect 15804 24012 15810 24064
rect 17770 24052 17776 24064
rect 17731 24024 17776 24052
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 18874 24052 18880 24064
rect 18835 24024 18880 24052
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 11422 23848 11428 23860
rect 11383 23820 11428 23848
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 11790 23848 11796 23860
rect 11751 23820 11796 23848
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 13722 23808 13728 23860
rect 13780 23848 13786 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 13780 23820 14933 23848
rect 13780 23808 13786 23820
rect 14921 23817 14933 23820
rect 14967 23817 14979 23851
rect 14921 23811 14979 23817
rect 16025 23851 16083 23857
rect 16025 23817 16037 23851
rect 16071 23848 16083 23851
rect 16114 23848 16120 23860
rect 16071 23820 16120 23848
rect 16071 23817 16083 23820
rect 16025 23811 16083 23817
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 16298 23848 16304 23860
rect 16259 23820 16304 23848
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 17034 23848 17040 23860
rect 16995 23820 17040 23848
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23712 15623 23715
rect 15746 23712 15752 23724
rect 15611 23684 15752 23712
rect 15611 23681 15623 23684
rect 15565 23675 15623 23681
rect 15746 23672 15752 23684
rect 15804 23672 15810 23724
rect 18874 23712 18880 23724
rect 18835 23684 18880 23712
rect 18874 23672 18880 23684
rect 18932 23672 18938 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 21913 23715 21971 23721
rect 21913 23712 21925 23715
rect 21784 23684 21925 23712
rect 21784 23672 21790 23684
rect 21913 23681 21925 23684
rect 21959 23681 21971 23715
rect 21913 23675 21971 23681
rect 24210 23672 24216 23724
rect 24268 23712 24274 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 24268 23684 25145 23712
rect 24268 23672 24274 23684
rect 25133 23681 25145 23684
rect 25179 23681 25191 23715
rect 25133 23675 25191 23681
rect 11241 23647 11299 23653
rect 11241 23613 11253 23647
rect 11287 23644 11299 23647
rect 11330 23644 11336 23656
rect 11287 23616 11336 23644
rect 11287 23613 11299 23616
rect 11241 23607 11299 23613
rect 11330 23604 11336 23616
rect 11388 23644 11394 23656
rect 12250 23644 12256 23656
rect 11388 23616 12256 23644
rect 11388 23604 11394 23616
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 12434 23644 12440 23656
rect 12395 23616 12440 23644
rect 12434 23604 12440 23616
rect 12492 23604 12498 23656
rect 12710 23653 12716 23656
rect 12704 23644 12716 23653
rect 12636 23616 12716 23644
rect 11149 23579 11207 23585
rect 11149 23545 11161 23579
rect 11195 23576 11207 23579
rect 12636 23576 12664 23616
rect 12704 23607 12716 23616
rect 12710 23604 12716 23607
rect 12768 23604 12774 23656
rect 14829 23647 14887 23653
rect 14829 23613 14841 23647
rect 14875 23644 14887 23647
rect 15381 23647 15439 23653
rect 15381 23644 15393 23647
rect 14875 23616 15393 23644
rect 14875 23613 14887 23616
rect 14829 23607 14887 23613
rect 15381 23613 15393 23616
rect 15427 23644 15439 23647
rect 16206 23644 16212 23656
rect 15427 23616 16212 23644
rect 15427 23613 15439 23616
rect 15381 23607 15439 23613
rect 16206 23604 16212 23616
rect 16264 23644 16270 23656
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 16264 23616 16865 23644
rect 16264 23604 16270 23616
rect 16853 23613 16865 23616
rect 16899 23644 16911 23647
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16899 23616 17417 23644
rect 16899 23613 16911 23616
rect 16853 23607 16911 23613
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 21634 23644 21640 23656
rect 17405 23607 17463 23613
rect 20824 23616 21640 23644
rect 11195 23548 12664 23576
rect 17865 23579 17923 23585
rect 11195 23545 11207 23548
rect 11149 23539 11207 23545
rect 17865 23545 17877 23579
rect 17911 23576 17923 23579
rect 18414 23576 18420 23588
rect 17911 23548 18420 23576
rect 17911 23545 17923 23548
rect 17865 23539 17923 23545
rect 18414 23536 18420 23548
rect 18472 23576 18478 23588
rect 19144 23579 19202 23585
rect 19144 23576 19156 23579
rect 18472 23548 19156 23576
rect 18472 23536 18478 23548
rect 19144 23545 19156 23548
rect 19190 23576 19202 23579
rect 19242 23576 19248 23588
rect 19190 23548 19248 23576
rect 19190 23545 19202 23548
rect 19144 23539 19202 23545
rect 19242 23536 19248 23548
rect 19300 23536 19306 23588
rect 20824 23520 20852 23616
rect 21634 23604 21640 23616
rect 21692 23644 21698 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21692 23616 21833 23644
rect 21692 23604 21698 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 21821 23607 21879 23613
rect 24412 23616 24593 23644
rect 21729 23579 21787 23585
rect 21729 23545 21741 23579
rect 21775 23576 21787 23579
rect 21910 23576 21916 23588
rect 21775 23548 21916 23576
rect 21775 23545 21787 23548
rect 21729 23539 21787 23545
rect 21910 23536 21916 23548
rect 21968 23576 21974 23588
rect 22922 23576 22928 23588
rect 21968 23548 22928 23576
rect 21968 23536 21974 23548
rect 22922 23536 22928 23548
rect 22980 23536 22986 23588
rect 8386 23468 8392 23520
rect 8444 23508 8450 23520
rect 9582 23508 9588 23520
rect 8444 23480 9588 23508
rect 8444 23468 8450 23480
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 12066 23468 12072 23520
rect 12124 23508 12130 23520
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 12124 23480 12173 23508
rect 12124 23468 12130 23480
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 12161 23471 12219 23477
rect 13446 23468 13452 23520
rect 13504 23508 13510 23520
rect 13817 23511 13875 23517
rect 13817 23508 13829 23511
rect 13504 23480 13829 23508
rect 13504 23468 13510 23480
rect 13817 23477 13829 23480
rect 13863 23508 13875 23511
rect 13998 23508 14004 23520
rect 13863 23480 14004 23508
rect 13863 23477 13875 23480
rect 13817 23471 13875 23477
rect 13998 23468 14004 23480
rect 14056 23508 14062 23520
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 14056 23480 14381 23508
rect 14056 23468 14062 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 15286 23508 15292 23520
rect 15247 23480 15292 23508
rect 14369 23471 14427 23477
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 16666 23508 16672 23520
rect 16627 23480 16672 23508
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 18322 23468 18328 23520
rect 18380 23508 18386 23520
rect 18693 23511 18751 23517
rect 18693 23508 18705 23511
rect 18380 23480 18705 23508
rect 18380 23468 18386 23480
rect 18693 23477 18705 23480
rect 18739 23477 18751 23511
rect 18693 23471 18751 23477
rect 20257 23511 20315 23517
rect 20257 23477 20269 23511
rect 20303 23508 20315 23511
rect 20622 23508 20628 23520
rect 20303 23480 20628 23508
rect 20303 23477 20315 23480
rect 20257 23471 20315 23477
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 20806 23508 20812 23520
rect 20767 23480 20812 23508
rect 20806 23468 20812 23480
rect 20864 23468 20870 23520
rect 21082 23468 21088 23520
rect 21140 23508 21146 23520
rect 21177 23511 21235 23517
rect 21177 23508 21189 23511
rect 21140 23480 21189 23508
rect 21140 23468 21146 23480
rect 21177 23477 21189 23480
rect 21223 23477 21235 23511
rect 21358 23508 21364 23520
rect 21319 23480 21364 23508
rect 21177 23471 21235 23477
rect 21358 23468 21364 23480
rect 21416 23468 21422 23520
rect 22370 23508 22376 23520
rect 22331 23480 22376 23508
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 23106 23468 23112 23520
rect 23164 23508 23170 23520
rect 23845 23511 23903 23517
rect 23845 23508 23857 23511
rect 23164 23480 23857 23508
rect 23164 23468 23170 23480
rect 23845 23477 23857 23480
rect 23891 23477 23903 23511
rect 23845 23471 23903 23477
rect 24118 23468 24124 23520
rect 24176 23508 24182 23520
rect 24412 23517 24440 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24176 23480 24409 23508
rect 24176 23468 24182 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 12989 23307 13047 23313
rect 12989 23273 13001 23307
rect 13035 23304 13047 23307
rect 13354 23304 13360 23316
rect 13035 23276 13360 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 13354 23264 13360 23276
rect 13412 23304 13418 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 13412 23276 13461 23304
rect 13412 23264 13418 23276
rect 13449 23273 13461 23276
rect 13495 23273 13507 23307
rect 13449 23267 13507 23273
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 15746 23304 15752 23316
rect 15611 23276 15752 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 15746 23264 15752 23276
rect 15804 23264 15810 23316
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 17129 23307 17187 23313
rect 17129 23304 17141 23307
rect 16632 23276 17141 23304
rect 16632 23264 16638 23276
rect 17129 23273 17141 23276
rect 17175 23304 17187 23307
rect 17402 23304 17408 23316
rect 17175 23276 17408 23304
rect 17175 23273 17187 23276
rect 17129 23267 17187 23273
rect 17402 23264 17408 23276
rect 17460 23264 17466 23316
rect 17678 23304 17684 23316
rect 17639 23276 17684 23304
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 18138 23304 18144 23316
rect 18099 23276 18144 23304
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 19613 23307 19671 23313
rect 19613 23304 19625 23307
rect 19392 23276 19625 23304
rect 19392 23264 19398 23276
rect 19613 23273 19625 23276
rect 19659 23273 19671 23307
rect 19613 23267 19671 23273
rect 21361 23307 21419 23313
rect 21361 23273 21373 23307
rect 21407 23304 21419 23307
rect 21634 23304 21640 23316
rect 21407 23276 21640 23304
rect 21407 23273 21419 23276
rect 21361 23267 21419 23273
rect 21634 23264 21640 23276
rect 21692 23304 21698 23316
rect 23382 23304 23388 23316
rect 21692 23276 23388 23304
rect 21692 23264 21698 23276
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 23658 23264 23664 23316
rect 23716 23304 23722 23316
rect 24026 23304 24032 23316
rect 23716 23276 24032 23304
rect 23716 23264 23722 23276
rect 24026 23264 24032 23276
rect 24084 23264 24090 23316
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 12621 23239 12679 23245
rect 12621 23236 12633 23239
rect 12492 23208 12633 23236
rect 12492 23196 12498 23208
rect 12621 23205 12633 23208
rect 12667 23236 12679 23239
rect 16016 23239 16074 23245
rect 12667 23208 15792 23236
rect 12667 23205 12679 23208
rect 12621 23199 12679 23205
rect 10870 23177 10876 23180
rect 10864 23131 10876 23177
rect 10928 23168 10934 23180
rect 15764 23177 15792 23208
rect 16016 23205 16028 23239
rect 16062 23236 16074 23239
rect 16390 23236 16396 23248
rect 16062 23208 16396 23236
rect 16062 23205 16074 23208
rect 16016 23199 16074 23205
rect 16390 23196 16396 23208
rect 16448 23196 16454 23248
rect 18874 23236 18880 23248
rect 18248 23208 18880 23236
rect 15749 23171 15807 23177
rect 10928 23140 13676 23168
rect 10870 23128 10876 23131
rect 10928 23128 10934 23140
rect 10594 23100 10600 23112
rect 10555 23072 10600 23100
rect 10594 23060 10600 23072
rect 10652 23060 10658 23112
rect 13538 23100 13544 23112
rect 13499 23072 13544 23100
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 13648 23109 13676 23140
rect 15749 23137 15761 23171
rect 15795 23168 15807 23171
rect 15838 23168 15844 23180
rect 15795 23140 15844 23168
rect 15795 23137 15807 23140
rect 15749 23131 15807 23137
rect 15838 23128 15844 23140
rect 15896 23168 15902 23180
rect 18248 23177 18276 23208
rect 18874 23196 18880 23208
rect 18932 23196 18938 23248
rect 18233 23171 18291 23177
rect 18233 23168 18245 23171
rect 15896 23140 18245 23168
rect 15896 23128 15902 23140
rect 18233 23137 18245 23140
rect 18279 23137 18291 23171
rect 18489 23171 18547 23177
rect 18489 23168 18501 23171
rect 18233 23131 18291 23137
rect 18340 23140 18501 23168
rect 13633 23103 13691 23109
rect 13633 23069 13645 23103
rect 13679 23100 13691 23103
rect 13814 23100 13820 23112
rect 13679 23072 13820 23100
rect 13679 23069 13691 23072
rect 13633 23063 13691 23069
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 14182 23100 14188 23112
rect 14143 23072 14188 23100
rect 14182 23060 14188 23072
rect 14240 23060 14246 23112
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 18340 23100 18368 23140
rect 18489 23137 18501 23140
rect 18535 23137 18547 23171
rect 18489 23131 18547 23137
rect 20990 23128 20996 23180
rect 21048 23168 21054 23180
rect 21269 23171 21327 23177
rect 21269 23168 21281 23171
rect 21048 23140 21281 23168
rect 21048 23128 21054 23140
rect 21269 23137 21281 23140
rect 21315 23137 21327 23171
rect 21269 23131 21327 23137
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 17460 23072 18368 23100
rect 17460 23060 17466 23072
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 21453 23103 21511 23109
rect 21453 23100 21465 23103
rect 20772 23072 21465 23100
rect 20772 23060 20778 23072
rect 21453 23069 21465 23072
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 23014 23060 23020 23112
rect 23072 23100 23078 23112
rect 23477 23103 23535 23109
rect 23477 23100 23489 23103
rect 23072 23072 23489 23100
rect 23072 23060 23078 23072
rect 23477 23069 23489 23072
rect 23523 23069 23535 23103
rect 23477 23063 23535 23069
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 23934 23100 23940 23112
rect 23707 23072 23940 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 23934 23060 23940 23072
rect 23992 23100 23998 23112
rect 24397 23103 24455 23109
rect 24397 23100 24409 23103
rect 23992 23072 24409 23100
rect 23992 23060 23998 23072
rect 24397 23069 24409 23072
rect 24443 23069 24455 23103
rect 24397 23063 24455 23069
rect 20898 23032 20904 23044
rect 20859 23004 20904 23032
rect 20898 22992 20904 23004
rect 20956 22992 20962 23044
rect 11974 22964 11980 22976
rect 11935 22936 11980 22964
rect 11974 22924 11980 22936
rect 12032 22924 12038 22976
rect 13078 22964 13084 22976
rect 13039 22936 13084 22964
rect 13078 22924 13084 22936
rect 13136 22924 13142 22976
rect 14826 22924 14832 22976
rect 14884 22964 14890 22976
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14884 22936 14933 22964
rect 14884 22924 14890 22936
rect 14921 22933 14933 22936
rect 14967 22964 14979 22967
rect 15286 22964 15292 22976
rect 14967 22936 15292 22964
rect 14967 22933 14979 22936
rect 14921 22927 14979 22933
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 21726 22924 21732 22976
rect 21784 22964 21790 22976
rect 21910 22964 21916 22976
rect 21784 22936 21916 22964
rect 21784 22924 21790 22936
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 22462 22924 22468 22976
rect 22520 22964 22526 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 22520 22936 23029 22964
rect 22520 22924 22526 22936
rect 23017 22933 23029 22936
rect 23063 22933 23075 22967
rect 23017 22927 23075 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 10870 22720 10876 22772
rect 10928 22760 10934 22772
rect 10965 22763 11023 22769
rect 10965 22760 10977 22763
rect 10928 22732 10977 22760
rect 10928 22720 10934 22732
rect 10965 22729 10977 22732
rect 11011 22729 11023 22763
rect 13814 22760 13820 22772
rect 13775 22732 13820 22760
rect 10965 22723 11023 22729
rect 13814 22720 13820 22732
rect 13872 22760 13878 22772
rect 14369 22763 14427 22769
rect 14369 22760 14381 22763
rect 13872 22732 14381 22760
rect 13872 22720 13878 22732
rect 14369 22729 14381 22732
rect 14415 22729 14427 22763
rect 14369 22723 14427 22729
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 15933 22763 15991 22769
rect 15933 22760 15945 22763
rect 15896 22732 15945 22760
rect 15896 22720 15902 22732
rect 15933 22729 15945 22732
rect 15979 22729 15991 22763
rect 16390 22760 16396 22772
rect 16351 22732 16396 22760
rect 15933 22723 15991 22729
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 16482 22720 16488 22772
rect 16540 22720 16546 22772
rect 17034 22760 17040 22772
rect 16995 22732 17040 22760
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 17494 22760 17500 22772
rect 17455 22732 17500 22760
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 18046 22760 18052 22772
rect 18007 22732 18052 22760
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 18874 22720 18880 22772
rect 18932 22760 18938 22772
rect 19061 22763 19119 22769
rect 19061 22760 19073 22763
rect 18932 22732 19073 22760
rect 18932 22720 18938 22732
rect 19061 22729 19073 22732
rect 19107 22760 19119 22763
rect 19981 22763 20039 22769
rect 19981 22760 19993 22763
rect 19107 22732 19993 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19981 22729 19993 22732
rect 20027 22729 20039 22763
rect 19981 22723 20039 22729
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 21910 22760 21916 22772
rect 21591 22732 21916 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 10652 22596 10701 22624
rect 10652 22584 10658 22596
rect 10689 22593 10701 22596
rect 10735 22624 10747 22627
rect 12253 22627 12311 22633
rect 12253 22624 12265 22627
rect 10735 22596 12265 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 12253 22593 12265 22596
rect 12299 22624 12311 22627
rect 12434 22624 12440 22636
rect 12299 22596 12440 22624
rect 12299 22593 12311 22596
rect 12253 22587 12311 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22624 15623 22627
rect 15746 22624 15752 22636
rect 15611 22596 15752 22624
rect 15611 22593 15623 22596
rect 15565 22587 15623 22593
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 16390 22516 16396 22568
rect 16448 22556 16454 22568
rect 16500 22556 16528 22720
rect 17402 22652 17408 22704
rect 17460 22692 17466 22704
rect 17773 22695 17831 22701
rect 17773 22692 17785 22695
rect 17460 22664 17785 22692
rect 17460 22652 17466 22664
rect 17773 22661 17785 22664
rect 17819 22692 17831 22695
rect 19429 22695 19487 22701
rect 19429 22692 19441 22695
rect 17819 22664 19441 22692
rect 17819 22661 17831 22664
rect 17773 22655 17831 22661
rect 18506 22624 18512 22636
rect 18467 22596 18512 22624
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 18616 22633 18644 22664
rect 19429 22661 19441 22664
rect 19475 22661 19487 22695
rect 19429 22655 19487 22661
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 19996 22624 20024 22723
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 23014 22760 23020 22772
rect 22975 22732 23020 22760
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 23382 22720 23388 22772
rect 23440 22720 23446 22772
rect 25406 22760 25412 22772
rect 25367 22732 25412 22760
rect 25406 22720 25412 22732
rect 25464 22720 25470 22772
rect 22741 22695 22799 22701
rect 22741 22661 22753 22695
rect 22787 22692 22799 22695
rect 23400 22692 23428 22720
rect 22787 22664 23428 22692
rect 22787 22661 22799 22664
rect 22741 22655 22799 22661
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 19996 22596 20177 22624
rect 18601 22587 18659 22593
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 22189 22627 22247 22633
rect 22189 22624 22201 22627
rect 20165 22587 20223 22593
rect 21836 22596 22201 22624
rect 16448 22528 16528 22556
rect 16448 22516 16454 22528
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16816 22528 16865 22556
rect 16816 22516 16822 22528
rect 16853 22525 16865 22528
rect 16899 22556 16911 22559
rect 17494 22556 17500 22568
rect 16899 22528 17500 22556
rect 16899 22525 16911 22528
rect 16853 22519 16911 22525
rect 17494 22516 17500 22528
rect 17552 22516 17558 22568
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 18196 22528 18429 22556
rect 18196 22516 18202 22528
rect 18417 22525 18429 22528
rect 18463 22525 18475 22559
rect 18417 22519 18475 22525
rect 20898 22516 20904 22568
rect 20956 22556 20962 22568
rect 21836 22556 21864 22596
rect 22189 22593 22201 22596
rect 22235 22624 22247 22627
rect 23290 22624 23296 22636
rect 22235 22596 23296 22624
rect 22235 22593 22247 22596
rect 22189 22587 22247 22593
rect 23290 22584 23296 22596
rect 23348 22584 23354 22636
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 23934 22624 23940 22636
rect 23440 22596 23940 22624
rect 23440 22584 23446 22596
rect 23934 22584 23940 22596
rect 23992 22624 23998 22636
rect 24213 22627 24271 22633
rect 24213 22624 24225 22627
rect 23992 22596 24225 22624
rect 23992 22584 23998 22596
rect 24213 22593 24225 22596
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 24026 22556 24032 22568
rect 20956 22528 21864 22556
rect 23987 22528 24032 22556
rect 20956 22516 20962 22528
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 12704 22491 12762 22497
rect 12704 22457 12716 22491
rect 12750 22488 12762 22491
rect 13446 22488 13452 22500
rect 12750 22460 13452 22488
rect 12750 22457 12762 22460
rect 12704 22451 12762 22457
rect 13446 22448 13452 22460
rect 13504 22448 13510 22500
rect 14829 22491 14887 22497
rect 14829 22457 14841 22491
rect 14875 22488 14887 22491
rect 14875 22460 15424 22488
rect 14875 22457 14887 22460
rect 14829 22451 14887 22457
rect 15396 22432 15424 22460
rect 20254 22448 20260 22500
rect 20312 22488 20318 22500
rect 20410 22491 20468 22497
rect 20410 22488 20422 22491
rect 20312 22460 20422 22488
rect 20312 22448 20318 22460
rect 20410 22457 20422 22460
rect 20456 22457 20468 22491
rect 20410 22451 20468 22457
rect 21726 22448 21732 22500
rect 21784 22488 21790 22500
rect 23106 22488 23112 22500
rect 21784 22460 23112 22488
rect 21784 22448 21790 22460
rect 23106 22448 23112 22460
rect 23164 22448 23170 22500
rect 24121 22491 24179 22497
rect 24121 22488 24133 22491
rect 23492 22460 24133 22488
rect 14918 22420 14924 22432
rect 14879 22392 14924 22420
rect 14918 22380 14924 22392
rect 14976 22380 14982 22432
rect 15286 22420 15292 22432
rect 15247 22392 15292 22420
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15436 22392 15481 22420
rect 15436 22380 15442 22392
rect 23290 22380 23296 22432
rect 23348 22420 23354 22432
rect 23492 22429 23520 22460
rect 24121 22457 24133 22460
rect 24167 22457 24179 22491
rect 24121 22451 24179 22457
rect 23477 22423 23535 22429
rect 23477 22420 23489 22423
rect 23348 22392 23489 22420
rect 23348 22380 23354 22392
rect 23477 22389 23489 22392
rect 23523 22389 23535 22423
rect 23658 22420 23664 22432
rect 23619 22392 23664 22420
rect 23477 22383 23535 22389
rect 23658 22380 23664 22392
rect 23716 22380 23722 22432
rect 23750 22380 23756 22432
rect 23808 22420 23814 22432
rect 24210 22420 24216 22432
rect 23808 22392 24216 22420
rect 23808 22380 23814 22392
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 24670 22420 24676 22432
rect 24631 22392 24676 22420
rect 24670 22380 24676 22392
rect 24728 22380 24734 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 12897 22219 12955 22225
rect 12897 22185 12909 22219
rect 12943 22216 12955 22219
rect 13538 22216 13544 22228
rect 12943 22188 13544 22216
rect 12943 22185 12955 22188
rect 12897 22179 12955 22185
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 15381 22219 15439 22225
rect 15381 22185 15393 22219
rect 15427 22216 15439 22219
rect 16666 22216 16672 22228
rect 15427 22188 16672 22216
rect 15427 22185 15439 22188
rect 15381 22179 15439 22185
rect 16666 22176 16672 22188
rect 16724 22176 16730 22228
rect 18141 22219 18199 22225
rect 18141 22185 18153 22219
rect 18187 22216 18199 22219
rect 18506 22216 18512 22228
rect 18187 22188 18512 22216
rect 18187 22185 18199 22188
rect 18141 22179 18199 22185
rect 18506 22176 18512 22188
rect 18564 22176 18570 22228
rect 18966 22216 18972 22228
rect 18927 22188 18972 22216
rect 18966 22176 18972 22188
rect 19024 22216 19030 22228
rect 19150 22216 19156 22228
rect 19024 22188 19156 22216
rect 19024 22176 19030 22188
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 20254 22216 20260 22228
rect 20215 22188 20260 22216
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 20714 22216 20720 22228
rect 20675 22188 20720 22216
rect 20714 22176 20720 22188
rect 20772 22176 20778 22228
rect 21634 22216 21640 22228
rect 21595 22188 21640 22216
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 22649 22219 22707 22225
rect 22649 22185 22661 22219
rect 22695 22216 22707 22219
rect 23017 22219 23075 22225
rect 23017 22216 23029 22219
rect 22695 22188 23029 22216
rect 22695 22185 22707 22188
rect 22649 22179 22707 22185
rect 23017 22185 23029 22188
rect 23063 22216 23075 22219
rect 23382 22216 23388 22228
rect 23063 22188 23388 22216
rect 23063 22185 23075 22188
rect 23017 22179 23075 22185
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 13265 22151 13323 22157
rect 13265 22117 13277 22151
rect 13311 22148 13323 22151
rect 13814 22148 13820 22160
rect 13311 22120 13820 22148
rect 13311 22117 13323 22120
rect 13265 22111 13323 22117
rect 13814 22108 13820 22120
rect 13872 22148 13878 22160
rect 14918 22148 14924 22160
rect 13872 22120 14924 22148
rect 13872 22108 13878 22120
rect 14918 22108 14924 22120
rect 14976 22108 14982 22160
rect 15749 22151 15807 22157
rect 15749 22148 15761 22151
rect 15120 22120 15761 22148
rect 12434 22040 12440 22092
rect 12492 22080 12498 22092
rect 13354 22080 13360 22092
rect 12492 22052 13360 22080
rect 12492 22040 12498 22052
rect 13354 22040 13360 22052
rect 13412 22040 13418 22092
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 13909 22083 13967 22089
rect 13909 22080 13921 22083
rect 13596 22052 13921 22080
rect 13596 22040 13602 22052
rect 13909 22049 13921 22052
rect 13955 22049 13967 22083
rect 13909 22043 13967 22049
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 13446 22012 13452 22024
rect 12575 21984 13452 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 13446 21972 13452 21984
rect 13504 21972 13510 22024
rect 14642 21972 14648 22024
rect 14700 22012 14706 22024
rect 15120 22012 15148 22120
rect 15749 22117 15761 22120
rect 15795 22117 15807 22151
rect 23658 22148 23664 22160
rect 15749 22111 15807 22117
rect 23216 22120 23664 22148
rect 17310 22080 17316 22092
rect 17271 22052 17316 22080
rect 17310 22040 17316 22052
rect 17368 22040 17374 22092
rect 19242 22080 19248 22092
rect 19076 22052 19248 22080
rect 15838 22012 15844 22024
rect 14700 21984 15148 22012
rect 15799 21984 15844 22012
rect 14700 21972 14706 21984
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 16298 22012 16304 22024
rect 16071 21984 16304 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 17402 22012 17408 22024
rect 16632 21984 17408 22012
rect 16632 21972 16638 21984
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 21981 17647 22015
rect 17589 21975 17647 21981
rect 16850 21904 16856 21956
rect 16908 21944 16914 21956
rect 17604 21944 17632 21975
rect 18138 21972 18144 22024
rect 18196 22012 18202 22024
rect 19076 22021 19104 22052
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22080 21143 22083
rect 21266 22080 21272 22092
rect 21131 22052 21272 22080
rect 21131 22049 21143 22052
rect 21085 22043 21143 22049
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 22094 22040 22100 22092
rect 22152 22080 22158 22092
rect 23216 22080 23244 22120
rect 23658 22108 23664 22120
rect 23716 22108 23722 22160
rect 23382 22089 23388 22092
rect 23376 22080 23388 22089
rect 22152 22052 22197 22080
rect 22572 22052 23244 22080
rect 23343 22052 23388 22080
rect 22152 22040 22158 22052
rect 19061 22015 19119 22021
rect 19061 22012 19073 22015
rect 18196 21984 19073 22012
rect 18196 21972 18202 21984
rect 19061 21981 19073 21984
rect 19107 21981 19119 22015
rect 19061 21975 19119 21981
rect 19153 22015 19211 22021
rect 19153 21981 19165 22015
rect 19199 21981 19211 22015
rect 19153 21975 19211 21981
rect 18509 21947 18567 21953
rect 18509 21944 18521 21947
rect 16908 21916 18521 21944
rect 16908 21904 16914 21916
rect 18509 21913 18521 21916
rect 18555 21944 18567 21947
rect 18690 21944 18696 21956
rect 18555 21916 18696 21944
rect 18555 21913 18567 21916
rect 18509 21907 18567 21913
rect 18690 21904 18696 21916
rect 18748 21944 18754 21956
rect 19168 21944 19196 21975
rect 21174 21972 21180 22024
rect 21232 22012 21238 22024
rect 21910 22012 21916 22024
rect 21232 21984 21916 22012
rect 21232 21972 21238 21984
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 22012 22063 22015
rect 22370 22012 22376 22024
rect 22051 21984 22376 22012
rect 22051 21981 22063 21984
rect 22005 21975 22063 21981
rect 22370 21972 22376 21984
rect 22428 22012 22434 22024
rect 22572 22012 22600 22052
rect 23376 22043 23388 22052
rect 23382 22040 23388 22043
rect 23440 22040 23446 22092
rect 24118 22040 24124 22092
rect 24176 22080 24182 22092
rect 24578 22080 24584 22092
rect 24176 22052 24584 22080
rect 24176 22040 24182 22052
rect 24578 22040 24584 22052
rect 24636 22040 24642 22092
rect 23106 22012 23112 22024
rect 22428 21984 22600 22012
rect 23067 21984 23112 22012
rect 22428 21972 22434 21984
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 18748 21916 19196 21944
rect 18748 21904 18754 21916
rect 10873 21879 10931 21885
rect 10873 21845 10885 21879
rect 10919 21876 10931 21879
rect 11974 21876 11980 21888
rect 10919 21848 11980 21876
rect 10919 21845 10931 21848
rect 10873 21839 10931 21845
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 12158 21876 12164 21888
rect 12119 21848 12164 21876
rect 12158 21836 12164 21848
rect 12216 21836 12222 21888
rect 15013 21879 15071 21885
rect 15013 21845 15025 21879
rect 15059 21876 15071 21879
rect 15286 21876 15292 21888
rect 15059 21848 15292 21876
rect 15059 21845 15071 21848
rect 15013 21839 15071 21845
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 16945 21879 17003 21885
rect 16945 21845 16957 21879
rect 16991 21876 17003 21879
rect 17126 21876 17132 21888
rect 16991 21848 17132 21876
rect 16991 21845 17003 21848
rect 16945 21839 17003 21845
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 18598 21876 18604 21888
rect 18559 21848 18604 21876
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19610 21876 19616 21888
rect 19571 21848 19616 21876
rect 19610 21836 19616 21848
rect 19668 21836 19674 21888
rect 21269 21879 21327 21885
rect 21269 21845 21281 21879
rect 21315 21876 21327 21879
rect 21910 21876 21916 21888
rect 21315 21848 21916 21876
rect 21315 21845 21327 21848
rect 21269 21839 21327 21845
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 22281 21879 22339 21885
rect 22281 21845 22293 21879
rect 22327 21876 22339 21879
rect 23290 21876 23296 21888
rect 22327 21848 23296 21876
rect 22327 21845 22339 21848
rect 22281 21839 22339 21845
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 24210 21836 24216 21888
rect 24268 21876 24274 21888
rect 24489 21879 24547 21885
rect 24489 21876 24501 21879
rect 24268 21848 24501 21876
rect 24268 21836 24274 21848
rect 24489 21845 24501 21848
rect 24535 21845 24547 21879
rect 24489 21839 24547 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 10594 21672 10600 21684
rect 10555 21644 10600 21672
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 13446 21672 13452 21684
rect 13407 21644 13452 21672
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 14642 21632 14648 21684
rect 14700 21672 14706 21684
rect 14737 21675 14795 21681
rect 14737 21672 14749 21675
rect 14700 21644 14749 21672
rect 14700 21632 14706 21644
rect 14737 21641 14749 21644
rect 14783 21641 14795 21675
rect 15930 21672 15936 21684
rect 15891 21644 15936 21672
rect 14737 21635 14795 21641
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 16298 21672 16304 21684
rect 16259 21644 16304 21672
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 16850 21672 16856 21684
rect 16811 21644 16856 21672
rect 16850 21632 16856 21644
rect 16908 21632 16914 21684
rect 17402 21672 17408 21684
rect 17363 21644 17408 21672
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 18874 21672 18880 21684
rect 18835 21644 18880 21672
rect 18874 21632 18880 21644
rect 18932 21632 18938 21684
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 20441 21675 20499 21681
rect 20441 21672 20453 21675
rect 20312 21644 20453 21672
rect 20312 21632 20318 21644
rect 20441 21641 20453 21644
rect 20487 21641 20499 21675
rect 20441 21635 20499 21641
rect 22005 21675 22063 21681
rect 22005 21641 22017 21675
rect 22051 21672 22063 21675
rect 22094 21672 22100 21684
rect 22051 21644 22100 21672
rect 22051 21641 22063 21644
rect 22005 21635 22063 21641
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 10612 21536 10640 21632
rect 11241 21539 11299 21545
rect 11241 21536 11253 21539
rect 10612 21508 11253 21536
rect 11241 21505 11253 21508
rect 11287 21505 11299 21539
rect 11241 21499 11299 21505
rect 11425 21539 11483 21545
rect 11425 21505 11437 21539
rect 11471 21536 11483 21539
rect 11974 21536 11980 21548
rect 11471 21508 11980 21536
rect 11471 21505 11483 21508
rect 11425 21499 11483 21505
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12115 21508 13093 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 13081 21505 13093 21508
rect 13127 21536 13139 21539
rect 13998 21536 14004 21548
rect 13127 21508 14004 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 15473 21539 15531 21545
rect 15473 21536 15485 21539
rect 14507 21508 15485 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 15473 21505 15485 21508
rect 15519 21536 15531 21539
rect 16022 21536 16028 21548
rect 15519 21508 16028 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 18892 21536 18920 21632
rect 21913 21607 21971 21613
rect 21913 21573 21925 21607
rect 21959 21604 21971 21607
rect 21959 21576 22600 21604
rect 21959 21573 21971 21576
rect 21913 21567 21971 21573
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 18892 21508 19073 21536
rect 19061 21505 19073 21508
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 21545 21539 21603 21545
rect 21545 21505 21557 21539
rect 21591 21536 21603 21539
rect 22462 21536 22468 21548
rect 21591 21508 22468 21536
rect 21591 21505 21603 21508
rect 21545 21499 21603 21505
rect 22462 21496 22468 21508
rect 22520 21496 22526 21548
rect 22572 21545 22600 21576
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21536 22615 21539
rect 23750 21536 23756 21548
rect 22603 21508 23756 21536
rect 22603 21505 22615 21508
rect 22557 21499 22615 21505
rect 23750 21496 23756 21508
rect 23808 21536 23814 21548
rect 23808 21508 24256 21536
rect 23808 21496 23814 21508
rect 24228 21480 24256 21508
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 12710 21468 12716 21480
rect 12216 21440 12716 21468
rect 12216 21428 12222 21440
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 14366 21428 14372 21480
rect 14424 21468 14430 21480
rect 14734 21468 14740 21480
rect 14424 21440 14740 21468
rect 14424 21428 14430 21440
rect 14734 21428 14740 21440
rect 14792 21428 14798 21480
rect 15286 21468 15292 21480
rect 15247 21440 15292 21468
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 19328 21471 19386 21477
rect 19328 21437 19340 21471
rect 19374 21468 19386 21471
rect 19610 21468 19616 21480
rect 19374 21440 19616 21468
rect 19374 21437 19386 21440
rect 19328 21431 19386 21437
rect 19610 21428 19616 21440
rect 19668 21428 19674 21480
rect 22370 21468 22376 21480
rect 22331 21440 22376 21468
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 24121 21471 24179 21477
rect 24121 21468 24133 21471
rect 23952 21440 24133 21468
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 12526 21400 12532 21412
rect 11931 21372 12532 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 12526 21360 12532 21372
rect 12584 21400 12590 21412
rect 12897 21403 12955 21409
rect 12897 21400 12909 21403
rect 12584 21372 12909 21400
rect 12584 21360 12590 21372
rect 12897 21369 12909 21372
rect 12943 21369 12955 21403
rect 15381 21403 15439 21409
rect 15381 21400 15393 21403
rect 12897 21363 12955 21369
rect 14016 21372 15393 21400
rect 10778 21332 10784 21344
rect 10739 21304 10784 21332
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11149 21335 11207 21341
rect 11149 21332 11161 21335
rect 11112 21304 11161 21332
rect 11112 21292 11118 21304
rect 11149 21301 11161 21304
rect 11195 21301 11207 21335
rect 11149 21295 11207 21301
rect 11238 21292 11244 21344
rect 11296 21332 11302 21344
rect 12069 21335 12127 21341
rect 12069 21332 12081 21335
rect 11296 21304 12081 21332
rect 11296 21292 11302 21304
rect 12069 21301 12081 21304
rect 12115 21332 12127 21335
rect 12161 21335 12219 21341
rect 12161 21332 12173 21335
rect 12115 21304 12173 21332
rect 12115 21301 12127 21304
rect 12069 21295 12127 21301
rect 12161 21301 12173 21304
rect 12207 21301 12219 21335
rect 12161 21295 12219 21301
rect 12437 21335 12495 21341
rect 12437 21301 12449 21335
rect 12483 21332 12495 21335
rect 12618 21332 12624 21344
rect 12483 21304 12624 21332
rect 12483 21301 12495 21304
rect 12437 21295 12495 21301
rect 12618 21292 12624 21304
rect 12676 21292 12682 21344
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 12805 21335 12863 21341
rect 12805 21332 12817 21335
rect 12768 21304 12817 21332
rect 12768 21292 12774 21304
rect 12805 21301 12817 21304
rect 12851 21301 12863 21335
rect 12805 21295 12863 21301
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 14016 21341 14044 21372
rect 15381 21369 15393 21372
rect 15427 21369 15439 21403
rect 15381 21363 15439 21369
rect 14001 21335 14059 21341
rect 14001 21332 14013 21335
rect 13780 21304 14013 21332
rect 13780 21292 13786 21304
rect 14001 21301 14013 21304
rect 14047 21301 14059 21335
rect 14918 21332 14924 21344
rect 14879 21304 14924 21332
rect 14001 21295 14059 21301
rect 14918 21292 14924 21304
rect 14976 21292 14982 21344
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17218 21332 17224 21344
rect 16991 21304 17224 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 17773 21335 17831 21341
rect 17773 21332 17785 21335
rect 17368 21304 17785 21332
rect 17368 21292 17374 21304
rect 17773 21301 17785 21304
rect 17819 21301 17831 21335
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 17773 21295 17831 21301
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 18196 21304 18521 21332
rect 18196 21292 18202 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 21177 21335 21235 21341
rect 21177 21301 21189 21335
rect 21223 21332 21235 21335
rect 21266 21332 21272 21344
rect 21223 21304 21272 21332
rect 21223 21301 21235 21304
rect 21177 21295 21235 21301
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 21818 21292 21824 21344
rect 21876 21332 21882 21344
rect 23106 21332 23112 21344
rect 21876 21304 23112 21332
rect 21876 21292 21882 21304
rect 23106 21292 23112 21304
rect 23164 21332 23170 21344
rect 23842 21332 23848 21344
rect 23164 21304 23848 21332
rect 23164 21292 23170 21304
rect 23842 21292 23848 21304
rect 23900 21332 23906 21344
rect 23952 21341 23980 21440
rect 24121 21437 24133 21440
rect 24167 21437 24179 21471
rect 24121 21431 24179 21437
rect 24210 21428 24216 21480
rect 24268 21468 24274 21480
rect 24377 21471 24435 21477
rect 24377 21468 24389 21471
rect 24268 21440 24389 21468
rect 24268 21428 24274 21440
rect 24377 21437 24389 21440
rect 24423 21437 24435 21471
rect 24377 21431 24435 21437
rect 23937 21335 23995 21341
rect 23937 21332 23949 21335
rect 23900 21304 23949 21332
rect 23900 21292 23906 21304
rect 23937 21301 23949 21304
rect 23983 21301 23995 21335
rect 25498 21332 25504 21344
rect 25459 21304 25504 21332
rect 23937 21295 23995 21301
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 13354 21128 13360 21140
rect 13315 21100 13360 21128
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 13814 21128 13820 21140
rect 13775 21100 13820 21128
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 13909 21131 13967 21137
rect 13909 21097 13921 21131
rect 13955 21128 13967 21131
rect 14826 21128 14832 21140
rect 13955 21100 14832 21128
rect 13955 21097 13967 21100
rect 13909 21091 13967 21097
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 15013 21131 15071 21137
rect 15013 21097 15025 21131
rect 15059 21128 15071 21131
rect 15286 21128 15292 21140
rect 15059 21100 15292 21128
rect 15059 21097 15071 21100
rect 15013 21091 15071 21097
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 17126 21128 17132 21140
rect 17087 21100 17132 21128
rect 17126 21088 17132 21100
rect 17184 21088 17190 21140
rect 17313 21131 17371 21137
rect 17313 21097 17325 21131
rect 17359 21128 17371 21131
rect 19337 21131 19395 21137
rect 19337 21128 19349 21131
rect 17359 21100 19349 21128
rect 17359 21097 17371 21100
rect 17313 21091 17371 21097
rect 19337 21097 19349 21100
rect 19383 21128 19395 21131
rect 19889 21131 19947 21137
rect 19889 21128 19901 21131
rect 19383 21100 19901 21128
rect 19383 21097 19395 21100
rect 19337 21091 19395 21097
rect 19889 21097 19901 21100
rect 19935 21097 19947 21131
rect 19889 21091 19947 21097
rect 21729 21131 21787 21137
rect 21729 21097 21741 21131
rect 21775 21128 21787 21131
rect 22094 21128 22100 21140
rect 21775 21100 22100 21128
rect 21775 21097 21787 21100
rect 21729 21091 21787 21097
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 23201 21131 23259 21137
rect 23201 21097 23213 21131
rect 23247 21128 23259 21131
rect 23382 21128 23388 21140
rect 23247 21100 23388 21128
rect 23247 21097 23259 21100
rect 23201 21091 23259 21097
rect 23382 21088 23388 21100
rect 23440 21088 23446 21140
rect 23750 21128 23756 21140
rect 23711 21100 23756 21128
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 11692 21063 11750 21069
rect 11692 21029 11704 21063
rect 11738 21060 11750 21063
rect 11974 21060 11980 21072
rect 11738 21032 11980 21060
rect 11738 21029 11750 21032
rect 11692 21023 11750 21029
rect 11974 21020 11980 21032
rect 12032 21020 12038 21072
rect 17144 21060 17172 21088
rect 17773 21063 17831 21069
rect 17773 21060 17785 21063
rect 17144 21032 17785 21060
rect 17773 21029 17785 21032
rect 17819 21029 17831 21063
rect 17773 21023 17831 21029
rect 18693 21063 18751 21069
rect 18693 21029 18705 21063
rect 18739 21060 18751 21063
rect 19150 21060 19156 21072
rect 18739 21032 19156 21060
rect 18739 21029 18751 21032
rect 18693 21023 18751 21029
rect 19150 21020 19156 21032
rect 19208 21020 19214 21072
rect 22922 21020 22928 21072
rect 22980 21060 22986 21072
rect 23566 21060 23572 21072
rect 22980 21032 23572 21060
rect 22980 21020 22986 21032
rect 23566 21020 23572 21032
rect 23624 21060 23630 21072
rect 24673 21063 24731 21069
rect 24673 21060 24685 21063
rect 23624 21032 24685 21060
rect 23624 21020 23630 21032
rect 24673 21029 24685 21032
rect 24719 21029 24731 21063
rect 24673 21023 24731 21029
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1946 20992 1952 21004
rect 1443 20964 1952 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1946 20952 1952 20964
rect 2004 20952 2010 21004
rect 15654 20952 15660 21004
rect 15712 20992 15718 21004
rect 15749 20995 15807 21001
rect 15749 20992 15761 20995
rect 15712 20964 15761 20992
rect 15712 20952 15718 20964
rect 15749 20961 15761 20964
rect 15795 20961 15807 20995
rect 15749 20955 15807 20961
rect 16853 20995 16911 21001
rect 16853 20961 16865 20995
rect 16899 20992 16911 20995
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 16899 20964 17693 20992
rect 16899 20961 16911 20964
rect 16853 20955 16911 20961
rect 17681 20961 17693 20964
rect 17727 20992 17739 20995
rect 18598 20992 18604 21004
rect 17727 20964 18604 20992
rect 17727 20961 17739 20964
rect 17681 20955 17739 20961
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 19242 20992 19248 21004
rect 19203 20964 19248 20992
rect 19242 20952 19248 20964
rect 19300 20952 19306 21004
rect 22094 21001 22100 21004
rect 22088 20955 22100 21001
rect 22152 20992 22158 21004
rect 22152 20964 22188 20992
rect 22094 20952 22100 20955
rect 22152 20952 22158 20964
rect 11422 20924 11428 20936
rect 11383 20896 11428 20924
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 15286 20884 15292 20936
rect 15344 20924 15350 20936
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 15344 20896 15853 20924
rect 15344 20884 15350 20896
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 16022 20924 16028 20936
rect 15983 20896 16028 20924
rect 15841 20887 15899 20893
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 17862 20924 17868 20936
rect 17823 20896 17868 20924
rect 17862 20884 17868 20896
rect 17920 20884 17926 20936
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 20254 20924 20260 20936
rect 19567 20896 20260 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 21818 20924 21824 20936
rect 21779 20896 21824 20924
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 23750 20884 23756 20936
rect 23808 20924 23814 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 23808 20896 24777 20924
rect 23808 20884 23814 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 25498 20924 25504 20936
rect 24995 20896 25504 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 1578 20856 1584 20868
rect 1539 20828 1584 20856
rect 1578 20816 1584 20828
rect 1636 20816 1642 20868
rect 24780 20856 24808 20887
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 25130 20856 25136 20868
rect 24780 20828 25136 20856
rect 25130 20816 25136 20828
rect 25188 20816 25194 20868
rect 10873 20791 10931 20797
rect 10873 20757 10885 20791
rect 10919 20788 10931 20791
rect 11054 20788 11060 20800
rect 10919 20760 11060 20788
rect 10919 20757 10931 20760
rect 10873 20751 10931 20757
rect 11054 20748 11060 20760
rect 11112 20788 11118 20800
rect 11698 20788 11704 20800
rect 11112 20760 11704 20788
rect 11112 20748 11118 20760
rect 11698 20748 11704 20760
rect 11756 20748 11762 20800
rect 12805 20791 12863 20797
rect 12805 20757 12817 20791
rect 12851 20788 12863 20791
rect 13170 20788 13176 20800
rect 12851 20760 13176 20788
rect 12851 20757 12863 20760
rect 12805 20751 12863 20757
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 15381 20791 15439 20797
rect 15381 20757 15393 20791
rect 15427 20788 15439 20791
rect 15746 20788 15752 20800
rect 15427 20760 15752 20788
rect 15427 20757 15439 20760
rect 15381 20751 15439 20757
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18012 20760 18889 20788
rect 18012 20748 18018 20760
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 18877 20751 18935 20757
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 20533 20791 20591 20797
rect 20533 20788 20545 20791
rect 20496 20760 20545 20788
rect 20496 20748 20502 20760
rect 20533 20757 20545 20760
rect 20579 20757 20591 20791
rect 24118 20788 24124 20800
rect 24079 20760 24124 20788
rect 20533 20751 20591 20757
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 24210 20748 24216 20800
rect 24268 20788 24274 20800
rect 24305 20791 24363 20797
rect 24305 20788 24317 20791
rect 24268 20760 24317 20788
rect 24268 20748 24274 20760
rect 24305 20757 24317 20760
rect 24351 20757 24363 20791
rect 24305 20751 24363 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 11241 20587 11299 20593
rect 11241 20553 11253 20587
rect 11287 20584 11299 20587
rect 11974 20584 11980 20596
rect 11287 20556 11980 20584
rect 11287 20553 11299 20556
rect 11241 20547 11299 20553
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12526 20584 12532 20596
rect 12483 20556 12532 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 16080 20556 16129 20584
rect 16080 20544 16086 20556
rect 16117 20553 16129 20556
rect 16163 20584 16175 20587
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 16163 20556 17049 20584
rect 16163 20553 16175 20556
rect 16117 20547 16175 20553
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 17037 20547 17095 20553
rect 17862 20544 17868 20596
rect 17920 20584 17926 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 17920 20556 19441 20584
rect 17920 20544 17926 20556
rect 19429 20553 19441 20556
rect 19475 20584 19487 20587
rect 19518 20584 19524 20596
rect 19475 20556 19524 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 20073 20587 20131 20593
rect 20073 20553 20085 20587
rect 20119 20584 20131 20587
rect 20254 20584 20260 20596
rect 20119 20556 20260 20584
rect 20119 20553 20131 20556
rect 20073 20547 20131 20553
rect 20254 20544 20260 20556
rect 20312 20544 20318 20596
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 22152 20556 22201 20584
rect 22152 20544 22158 20556
rect 22189 20553 22201 20556
rect 22235 20553 22247 20587
rect 22189 20547 22247 20553
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 23566 20584 23572 20596
rect 23523 20556 23572 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 24026 20544 24032 20596
rect 24084 20584 24090 20596
rect 25314 20584 25320 20596
rect 24084 20556 25320 20584
rect 24084 20544 24090 20556
rect 25314 20544 25320 20556
rect 25372 20544 25378 20596
rect 25498 20584 25504 20596
rect 25459 20556 25504 20584
rect 25498 20544 25504 20556
rect 25556 20584 25562 20596
rect 25869 20587 25927 20593
rect 25869 20584 25881 20587
rect 25556 20556 25881 20584
rect 25556 20544 25562 20556
rect 25869 20553 25881 20556
rect 25915 20553 25927 20587
rect 25869 20547 25927 20553
rect 12894 20448 12900 20460
rect 12855 20420 12900 20448
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 13170 20448 13176 20460
rect 13127 20420 13176 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20772 20420 21097 20448
rect 20772 20408 20778 20420
rect 21085 20417 21097 20420
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20448 24823 20451
rect 25038 20448 25044 20460
rect 24811 20420 25044 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 25038 20408 25044 20420
rect 25096 20448 25102 20460
rect 25516 20448 25544 20544
rect 25096 20420 25544 20448
rect 25096 20408 25102 20420
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 12912 20380 12940 20408
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 12912 20352 13829 20380
rect 13817 20349 13829 20352
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20380 14795 20383
rect 15470 20380 15476 20392
rect 14783 20352 15476 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 15470 20340 15476 20352
rect 15528 20380 15534 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 15528 20352 17877 20380
rect 15528 20340 15534 20352
rect 17865 20349 17877 20352
rect 17911 20380 17923 20383
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 17911 20352 18061 20380
rect 17911 20349 17923 20352
rect 17865 20343 17923 20349
rect 18049 20349 18061 20352
rect 18095 20380 18107 20383
rect 18874 20380 18880 20392
rect 18095 20352 18880 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 20441 20383 20499 20389
rect 20441 20349 20453 20383
rect 20487 20380 20499 20383
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20487 20352 21005 20380
rect 20487 20349 20499 20352
rect 20441 20343 20499 20349
rect 20993 20349 21005 20352
rect 21039 20380 21051 20383
rect 21634 20380 21640 20392
rect 21039 20352 21640 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20380 22615 20383
rect 24118 20380 24124 20392
rect 22603 20352 24124 20380
rect 22603 20349 22615 20352
rect 22557 20343 22615 20349
rect 24118 20340 24124 20352
rect 24176 20380 24182 20392
rect 24489 20383 24547 20389
rect 24489 20380 24501 20383
rect 24176 20352 24501 20380
rect 24176 20340 24182 20352
rect 24489 20349 24501 20352
rect 24535 20349 24547 20383
rect 24489 20343 24547 20349
rect 12253 20315 12311 20321
rect 12253 20281 12265 20315
rect 12299 20312 12311 20315
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 12299 20284 12817 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 12805 20281 12817 20284
rect 12851 20312 12863 20315
rect 13262 20312 13268 20324
rect 12851 20284 13268 20312
rect 12851 20281 12863 20284
rect 12805 20275 12863 20281
rect 13262 20272 13268 20284
rect 13320 20272 13326 20324
rect 14982 20315 15040 20321
rect 14982 20312 14994 20315
rect 14200 20284 14994 20312
rect 14200 20256 14228 20284
rect 14982 20281 14994 20284
rect 15028 20281 15040 20315
rect 14982 20275 15040 20281
rect 17497 20315 17555 20321
rect 17497 20281 17509 20315
rect 17543 20312 17555 20315
rect 18316 20315 18374 20321
rect 18316 20312 18328 20315
rect 17543 20284 18328 20312
rect 17543 20281 17555 20284
rect 17497 20275 17555 20281
rect 18316 20281 18328 20284
rect 18362 20312 18374 20315
rect 18690 20312 18696 20324
rect 18362 20284 18696 20312
rect 18362 20281 18374 20284
rect 18316 20275 18374 20281
rect 18690 20272 18696 20284
rect 18748 20272 18754 20324
rect 24581 20315 24639 20321
rect 24581 20312 24593 20315
rect 23952 20284 24593 20312
rect 23952 20256 23980 20284
rect 24581 20281 24593 20284
rect 24627 20312 24639 20315
rect 24854 20312 24860 20324
rect 24627 20284 24860 20312
rect 24627 20281 24639 20284
rect 24581 20275 24639 20281
rect 24854 20272 24860 20284
rect 24912 20272 24918 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 10321 20247 10379 20253
rect 10321 20213 10333 20247
rect 10367 20244 10379 20247
rect 10962 20244 10968 20256
rect 10367 20216 10968 20244
rect 10367 20213 10379 20216
rect 10321 20207 10379 20213
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 11330 20244 11336 20256
rect 11291 20216 11336 20244
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11882 20244 11888 20256
rect 11480 20216 11888 20244
rect 11480 20204 11486 20216
rect 11882 20204 11888 20216
rect 11940 20204 11946 20256
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 13449 20247 13507 20253
rect 13449 20244 13461 20247
rect 13228 20216 13461 20244
rect 13228 20204 13234 20216
rect 13449 20213 13461 20216
rect 13495 20213 13507 20247
rect 14182 20244 14188 20256
rect 14143 20216 14188 20244
rect 13449 20207 13507 20213
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 14366 20204 14372 20256
rect 14424 20244 14430 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14424 20216 14565 20244
rect 14424 20204 14430 20216
rect 14553 20213 14565 20216
rect 14599 20244 14611 20247
rect 15286 20244 15292 20256
rect 14599 20216 15292 20244
rect 14599 20213 14611 20216
rect 14553 20207 14611 20213
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 20530 20244 20536 20256
rect 20491 20216 20536 20244
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 21818 20244 21824 20256
rect 21779 20216 21824 20244
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 23934 20244 23940 20256
rect 23895 20216 23940 20244
rect 23934 20204 23940 20216
rect 23992 20204 23998 20256
rect 24118 20244 24124 20256
rect 24079 20216 24124 20244
rect 24118 20204 24124 20216
rect 24176 20204 24182 20256
rect 25130 20244 25136 20256
rect 25091 20216 25136 20244
rect 25130 20204 25136 20216
rect 25188 20204 25194 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 12526 20040 12532 20052
rect 11388 20012 12532 20040
rect 11388 20000 11394 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 13998 20000 14004 20052
rect 14056 20040 14062 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 14056 20012 14105 20040
rect 14056 20000 14062 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 14093 20003 14151 20009
rect 17497 20043 17555 20049
rect 17497 20009 17509 20043
rect 17543 20040 17555 20043
rect 17862 20040 17868 20052
rect 17543 20012 17868 20040
rect 17543 20009 17555 20012
rect 17497 20003 17555 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18046 20040 18052 20052
rect 18007 20012 18052 20040
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19242 20040 19248 20052
rect 18739 20012 19248 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19242 20000 19248 20012
rect 19300 20040 19306 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 19300 20012 20085 20040
rect 19300 20000 19306 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 20073 20003 20131 20009
rect 20625 20043 20683 20049
rect 20625 20009 20637 20043
rect 20671 20040 20683 20043
rect 20898 20040 20904 20052
rect 20671 20012 20904 20040
rect 20671 20009 20683 20012
rect 20625 20003 20683 20009
rect 20898 20000 20904 20012
rect 20956 20000 20962 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 22152 20012 22293 20040
rect 22152 20000 22158 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 22281 20003 22339 20009
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20040 23903 20043
rect 24118 20040 24124 20052
rect 23891 20012 24124 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 11422 19972 11428 19984
rect 10244 19944 11428 19972
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10244 19913 10272 19944
rect 11422 19932 11428 19944
rect 11480 19932 11486 19984
rect 12980 19975 13038 19981
rect 12980 19941 12992 19975
rect 13026 19972 13038 19975
rect 13170 19972 13176 19984
rect 13026 19944 13176 19972
rect 13026 19941 13038 19944
rect 12980 19935 13038 19941
rect 13170 19932 13176 19944
rect 13228 19932 13234 19984
rect 15740 19975 15798 19981
rect 15740 19941 15752 19975
rect 15786 19972 15798 19975
rect 16022 19972 16028 19984
rect 15786 19944 16028 19972
rect 15786 19941 15798 19944
rect 15740 19935 15798 19941
rect 16022 19932 16028 19944
rect 16080 19932 16086 19984
rect 19153 19975 19211 19981
rect 19153 19941 19165 19975
rect 19199 19972 19211 19975
rect 19518 19972 19524 19984
rect 19199 19944 19524 19972
rect 19199 19941 19211 19944
rect 19153 19935 19211 19941
rect 19518 19932 19524 19944
rect 19576 19972 19582 19984
rect 20530 19972 20536 19984
rect 19576 19944 20536 19972
rect 19576 19932 19582 19944
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 24204 19975 24262 19981
rect 24204 19941 24216 19975
rect 24250 19972 24262 19975
rect 25038 19972 25044 19984
rect 24250 19944 25044 19972
rect 24250 19941 24262 19944
rect 24204 19935 24262 19941
rect 25038 19932 25044 19944
rect 25096 19932 25102 19984
rect 10229 19907 10287 19913
rect 10229 19904 10241 19907
rect 9916 19876 10241 19904
rect 9916 19864 9922 19876
rect 10229 19873 10241 19876
rect 10275 19873 10287 19907
rect 10229 19867 10287 19873
rect 10318 19864 10324 19916
rect 10376 19904 10382 19916
rect 10485 19907 10543 19913
rect 10485 19904 10497 19907
rect 10376 19876 10497 19904
rect 10376 19864 10382 19876
rect 10485 19873 10497 19876
rect 10531 19904 10543 19907
rect 11238 19904 11244 19916
rect 10531 19876 11244 19904
rect 10531 19873 10543 19876
rect 10485 19867 10543 19873
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 11940 19876 12725 19904
rect 11940 19864 11946 19876
rect 12713 19873 12725 19876
rect 12759 19904 12771 19907
rect 13538 19904 13544 19916
rect 12759 19876 13544 19904
rect 12759 19873 12771 19876
rect 12713 19867 12771 19873
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 18598 19904 18604 19916
rect 18511 19876 18604 19904
rect 18598 19864 18604 19876
rect 18656 19904 18662 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 18656 19876 19073 19904
rect 18656 19864 18662 19876
rect 19061 19873 19073 19876
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 19797 19907 19855 19913
rect 19797 19873 19809 19907
rect 19843 19904 19855 19907
rect 20070 19904 20076 19916
rect 19843 19876 20076 19904
rect 19843 19873 19855 19876
rect 19797 19867 19855 19873
rect 20070 19864 20076 19876
rect 20128 19904 20134 19916
rect 20622 19904 20628 19916
rect 20128 19876 20628 19904
rect 20128 19864 20134 19876
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 20990 19864 20996 19916
rect 21048 19904 21054 19916
rect 21157 19907 21215 19913
rect 21157 19904 21169 19907
rect 21048 19876 21169 19904
rect 21048 19864 21054 19876
rect 21157 19873 21169 19876
rect 21203 19873 21215 19907
rect 21157 19867 21215 19873
rect 23842 19864 23848 19916
rect 23900 19904 23906 19916
rect 23937 19907 23995 19913
rect 23937 19904 23949 19907
rect 23900 19876 23949 19904
rect 23900 19864 23906 19876
rect 23937 19873 23949 19876
rect 23983 19873 23995 19907
rect 23937 19867 23995 19873
rect 19242 19796 19248 19848
rect 19300 19836 19306 19848
rect 19337 19839 19395 19845
rect 19337 19836 19349 19839
rect 19300 19808 19349 19836
rect 19300 19796 19306 19808
rect 19337 19805 19349 19808
rect 19383 19836 19395 19839
rect 19426 19836 19432 19848
rect 19383 19808 19432 19836
rect 19383 19805 19395 19808
rect 19337 19799 19395 19805
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 20898 19836 20904 19848
rect 20859 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 1581 19703 1639 19709
rect 1581 19700 1593 19703
rect 1452 19672 1593 19700
rect 1452 19660 1458 19672
rect 1581 19669 1593 19672
rect 1627 19669 1639 19703
rect 11606 19700 11612 19712
rect 11567 19672 11612 19700
rect 1581 19663 1639 19669
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 16850 19700 16856 19712
rect 16811 19672 16856 19700
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 25314 19700 25320 19712
rect 25275 19672 25320 19700
rect 25314 19660 25320 19672
rect 25372 19660 25378 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 9493 19499 9551 19505
rect 9493 19465 9505 19499
rect 9539 19496 9551 19499
rect 10318 19496 10324 19508
rect 9539 19468 10324 19496
rect 9539 19465 9551 19468
rect 9493 19459 9551 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 13538 19496 13544 19508
rect 13451 19468 13544 19496
rect 13538 19456 13544 19468
rect 13596 19496 13602 19508
rect 14093 19499 14151 19505
rect 14093 19496 14105 19499
rect 13596 19468 14105 19496
rect 13596 19456 13602 19468
rect 14093 19465 14105 19468
rect 14139 19496 14151 19499
rect 14139 19468 15516 19496
rect 14139 19465 14151 19468
rect 14093 19459 14151 19465
rect 9858 19428 9864 19440
rect 9819 19400 9864 19428
rect 9858 19388 9864 19400
rect 9916 19388 9922 19440
rect 10962 19360 10968 19372
rect 10923 19332 10968 19360
rect 10962 19320 10968 19332
rect 11020 19360 11026 19372
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 11020 19332 11345 19360
rect 11020 19320 11026 19332
rect 11333 19329 11345 19332
rect 11379 19360 11391 19363
rect 11606 19360 11612 19372
rect 11379 19332 11612 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12268 19332 13093 19360
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10137 19295 10195 19301
rect 10137 19292 10149 19295
rect 9732 19264 10149 19292
rect 9732 19252 9738 19264
rect 10137 19261 10149 19264
rect 10183 19292 10195 19295
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 10183 19264 10701 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 11885 19295 11943 19301
rect 11885 19261 11897 19295
rect 11931 19292 11943 19295
rect 12268 19292 12296 19332
rect 13081 19329 13093 19332
rect 13127 19360 13139 19363
rect 13170 19360 13176 19372
rect 13127 19332 13176 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 14200 19369 14228 19468
rect 15488 19440 15516 19468
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 15933 19499 15991 19505
rect 15933 19496 15945 19499
rect 15712 19468 15945 19496
rect 15712 19456 15718 19468
rect 15933 19465 15945 19468
rect 15979 19465 15991 19499
rect 15933 19459 15991 19465
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 16485 19499 16543 19505
rect 16485 19496 16497 19499
rect 16080 19468 16497 19496
rect 16080 19456 16086 19468
rect 16485 19465 16497 19468
rect 16531 19465 16543 19499
rect 16485 19459 16543 19465
rect 18049 19499 18107 19505
rect 18049 19465 18061 19499
rect 18095 19496 18107 19499
rect 18598 19496 18604 19508
rect 18095 19468 18604 19496
rect 18095 19465 18107 19468
rect 18049 19459 18107 19465
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 21266 19496 21272 19508
rect 21227 19468 21272 19496
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22281 19499 22339 19505
rect 22281 19496 22293 19499
rect 22152 19468 22293 19496
rect 22152 19456 22158 19468
rect 22281 19465 22293 19468
rect 22327 19465 22339 19499
rect 24854 19496 24860 19508
rect 22281 19459 22339 19465
rect 23032 19468 24860 19496
rect 15470 19388 15476 19440
rect 15528 19428 15534 19440
rect 16114 19428 16120 19440
rect 15528 19400 16120 19428
rect 15528 19388 15534 19400
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 20898 19428 20904 19440
rect 20859 19400 20904 19428
rect 20898 19388 20904 19400
rect 20956 19428 20962 19440
rect 21818 19428 21824 19440
rect 20956 19400 21824 19428
rect 20956 19388 20962 19400
rect 21818 19388 21824 19400
rect 21876 19388 21882 19440
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 16022 19360 16028 19372
rect 15979 19332 16028 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19360 17555 19363
rect 18690 19360 18696 19372
rect 17543 19332 18696 19360
rect 17543 19329 17555 19332
rect 17497 19323 17555 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 19260 19332 20269 19360
rect 11931 19264 12296 19292
rect 11931 19261 11943 19264
rect 11885 19255 11943 19261
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12584 19264 12817 19292
rect 12584 19252 12590 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 16666 19292 16672 19304
rect 16627 19264 16672 19292
rect 12805 19255 12863 19261
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 18046 19252 18052 19304
rect 18104 19292 18110 19304
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 18104 19264 18429 19292
rect 18104 19252 18110 19264
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 12253 19227 12311 19233
rect 12253 19193 12265 19227
rect 12299 19224 12311 19227
rect 14452 19227 14510 19233
rect 12299 19196 12940 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 12912 19168 12940 19196
rect 14452 19193 14464 19227
rect 14498 19224 14510 19227
rect 14642 19224 14648 19236
rect 14498 19196 14648 19224
rect 14498 19193 14510 19196
rect 14452 19187 14510 19193
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 17770 19224 17776 19236
rect 16868 19196 17776 19224
rect 10321 19159 10379 19165
rect 10321 19125 10333 19159
rect 10367 19156 10379 19159
rect 10686 19156 10692 19168
rect 10367 19128 10692 19156
rect 10367 19125 10379 19128
rect 10321 19119 10379 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 10781 19159 10839 19165
rect 10781 19125 10793 19159
rect 10827 19156 10839 19159
rect 10870 19156 10876 19168
rect 10827 19128 10876 19156
rect 10827 19125 10839 19128
rect 10781 19119 10839 19125
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 12437 19159 12495 19165
rect 12437 19125 12449 19159
rect 12483 19156 12495 19159
rect 12710 19156 12716 19168
rect 12483 19128 12716 19156
rect 12483 19125 12495 19128
rect 12437 19119 12495 19125
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 12894 19156 12900 19168
rect 12855 19128 12900 19156
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 16868 19165 16896 19196
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 14240 19128 15577 19156
rect 14240 19116 14246 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 16853 19159 16911 19165
rect 16853 19125 16865 19159
rect 16899 19125 16911 19159
rect 16853 19119 16911 19125
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17865 19159 17923 19165
rect 17865 19156 17877 19159
rect 17000 19128 17877 19156
rect 17000 19116 17006 19128
rect 17865 19125 17877 19128
rect 17911 19156 17923 19159
rect 18509 19159 18567 19165
rect 18509 19156 18521 19159
rect 17911 19128 18521 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 18509 19125 18521 19128
rect 18555 19156 18567 19159
rect 18690 19156 18696 19168
rect 18555 19128 18696 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19150 19156 19156 19168
rect 19111 19128 19156 19156
rect 19150 19116 19156 19128
rect 19208 19156 19214 19168
rect 19260 19156 19288 19332
rect 20257 19329 20269 19332
rect 20303 19360 20315 19363
rect 20990 19360 20996 19372
rect 20303 19332 20996 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21913 19363 21971 19369
rect 21913 19329 21925 19363
rect 21959 19360 21971 19363
rect 22112 19360 22140 19456
rect 22922 19388 22928 19440
rect 22980 19428 22986 19440
rect 23032 19428 23060 19468
rect 24854 19456 24860 19468
rect 24912 19456 24918 19508
rect 25038 19496 25044 19508
rect 24999 19468 25044 19496
rect 25038 19456 25044 19468
rect 25096 19456 25102 19508
rect 22980 19400 23060 19428
rect 22980 19388 22986 19400
rect 23934 19388 23940 19440
rect 23992 19428 23998 19440
rect 24302 19428 24308 19440
rect 23992 19400 24308 19428
rect 23992 19388 23998 19400
rect 24302 19388 24308 19400
rect 24360 19388 24366 19440
rect 24578 19360 24584 19372
rect 21959 19332 22140 19360
rect 23584 19332 24584 19360
rect 21959 19329 21971 19332
rect 21913 19323 21971 19329
rect 20070 19292 20076 19304
rect 20031 19264 20076 19292
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19292 23167 19295
rect 23584 19292 23612 19332
rect 24578 19320 24584 19332
rect 24636 19360 24642 19372
rect 25314 19360 25320 19372
rect 24636 19332 25320 19360
rect 24636 19320 24642 19332
rect 25314 19320 25320 19332
rect 25372 19320 25378 19372
rect 23155 19264 23612 19292
rect 23155 19261 23167 19264
rect 23109 19255 23167 19261
rect 24118 19252 24124 19304
rect 24176 19292 24182 19304
rect 24305 19295 24363 19301
rect 24305 19292 24317 19295
rect 24176 19264 24317 19292
rect 24176 19252 24182 19264
rect 24305 19261 24317 19264
rect 24351 19261 24363 19295
rect 25498 19292 25504 19304
rect 25459 19264 25504 19292
rect 24305 19255 24363 19261
rect 25498 19252 25504 19264
rect 25556 19292 25562 19304
rect 26053 19295 26111 19301
rect 26053 19292 26065 19295
rect 25556 19264 26065 19292
rect 25556 19252 25562 19264
rect 26053 19261 26065 19264
rect 26099 19261 26111 19295
rect 26053 19255 26111 19261
rect 21729 19227 21787 19233
rect 21729 19224 21741 19227
rect 19996 19196 21741 19224
rect 19996 19168 20024 19196
rect 21729 19193 21741 19196
rect 21775 19193 21787 19227
rect 21729 19187 21787 19193
rect 23477 19227 23535 19233
rect 23477 19193 23489 19227
rect 23523 19224 23535 19227
rect 23842 19224 23848 19236
rect 23523 19196 23848 19224
rect 23523 19193 23535 19196
rect 23477 19187 23535 19193
rect 23842 19184 23848 19196
rect 23900 19184 23906 19236
rect 24210 19184 24216 19236
rect 24268 19224 24274 19236
rect 24397 19227 24455 19233
rect 24397 19224 24409 19227
rect 24268 19196 24409 19224
rect 24268 19184 24274 19196
rect 24397 19193 24409 19196
rect 24443 19224 24455 19227
rect 25317 19227 25375 19233
rect 25317 19224 25329 19227
rect 24443 19196 25329 19224
rect 24443 19193 24455 19196
rect 24397 19187 24455 19193
rect 25317 19193 25329 19196
rect 25363 19193 25375 19227
rect 25317 19187 25375 19193
rect 19208 19128 19288 19156
rect 19208 19116 19214 19128
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19521 19159 19579 19165
rect 19521 19156 19533 19159
rect 19484 19128 19533 19156
rect 19484 19116 19490 19128
rect 19521 19125 19533 19128
rect 19567 19125 19579 19159
rect 19521 19119 19579 19125
rect 19705 19159 19763 19165
rect 19705 19125 19717 19159
rect 19751 19156 19763 19159
rect 19978 19156 19984 19168
rect 19751 19128 19984 19156
rect 19751 19125 19763 19128
rect 19705 19119 19763 19125
rect 19978 19116 19984 19128
rect 20036 19116 20042 19168
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 20128 19128 20177 19156
rect 20128 19116 20134 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 21634 19156 21640 19168
rect 21595 19128 21640 19156
rect 20165 19119 20223 19125
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 22738 19156 22744 19168
rect 22699 19128 22744 19156
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 23934 19156 23940 19168
rect 23895 19128 23940 19156
rect 23934 19116 23940 19128
rect 23992 19116 23998 19168
rect 25682 19156 25688 19168
rect 25643 19128 25688 19156
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 12802 18952 12808 18964
rect 12763 18924 12808 18952
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 13170 18952 13176 18964
rect 13131 18924 13176 18952
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 13722 18952 13728 18964
rect 13679 18924 13728 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14001 18955 14059 18961
rect 14001 18952 14013 18955
rect 13964 18924 14013 18952
rect 13964 18912 13970 18924
rect 14001 18921 14013 18924
rect 14047 18921 14059 18955
rect 14642 18952 14648 18964
rect 14603 18924 14648 18952
rect 14001 18915 14059 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 15381 18955 15439 18961
rect 15381 18921 15393 18955
rect 15427 18952 15439 18955
rect 16666 18952 16672 18964
rect 15427 18924 16672 18952
rect 15427 18921 15439 18924
rect 15381 18915 15439 18921
rect 16666 18912 16672 18924
rect 16724 18952 16730 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 16724 18924 16773 18952
rect 16724 18912 16730 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 18509 18955 18567 18961
rect 18509 18921 18521 18955
rect 18555 18952 18567 18955
rect 19150 18952 19156 18964
rect 18555 18924 19156 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 19518 18952 19524 18964
rect 19479 18924 19524 18952
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 20625 18955 20683 18961
rect 20625 18952 20637 18955
rect 20036 18924 20637 18952
rect 20036 18912 20042 18924
rect 20625 18921 20637 18924
rect 20671 18921 20683 18955
rect 20625 18915 20683 18921
rect 21177 18955 21235 18961
rect 21177 18921 21189 18955
rect 21223 18952 21235 18955
rect 21634 18952 21640 18964
rect 21223 18924 21640 18952
rect 21223 18921 21235 18924
rect 21177 18915 21235 18921
rect 21634 18912 21640 18924
rect 21692 18952 21698 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 21692 18924 22569 18952
rect 21692 18912 21698 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 23658 18952 23664 18964
rect 23619 18924 23664 18952
rect 22557 18915 22615 18921
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 24302 18952 24308 18964
rect 23768 18924 24308 18952
rect 13814 18844 13820 18896
rect 13872 18884 13878 18896
rect 14093 18887 14151 18893
rect 14093 18884 14105 18887
rect 13872 18856 14105 18884
rect 13872 18844 13878 18856
rect 14016 18828 14044 18856
rect 14093 18853 14105 18856
rect 14139 18853 14151 18887
rect 15746 18884 15752 18896
rect 15707 18856 15752 18884
rect 14093 18847 14151 18853
rect 15746 18844 15752 18856
rect 15804 18884 15810 18896
rect 16393 18887 16451 18893
rect 16393 18884 16405 18887
rect 15804 18856 16405 18884
rect 15804 18844 15810 18856
rect 16393 18853 16405 18856
rect 16439 18853 16451 18887
rect 16393 18847 16451 18853
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 20070 18884 20076 18896
rect 19484 18856 20076 18884
rect 19484 18844 19490 18856
rect 20070 18844 20076 18856
rect 20128 18844 20134 18896
rect 21542 18884 21548 18896
rect 21503 18856 21548 18884
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 23768 18884 23796 18924
rect 24302 18912 24308 18924
rect 24360 18912 24366 18964
rect 22572 18856 23796 18884
rect 24112 18887 24170 18893
rect 22572 18828 22600 18856
rect 24112 18853 24124 18887
rect 24158 18884 24170 18887
rect 24210 18884 24216 18896
rect 24158 18856 24216 18884
rect 24158 18853 24170 18856
rect 24112 18847 24170 18853
rect 24210 18844 24216 18856
rect 24268 18884 24274 18896
rect 24578 18884 24584 18896
rect 24268 18856 24584 18884
rect 24268 18844 24274 18856
rect 24578 18844 24584 18856
rect 24636 18844 24642 18896
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10962 18825 10968 18828
rect 10945 18819 10968 18825
rect 10945 18816 10957 18819
rect 10376 18788 10957 18816
rect 10376 18776 10382 18788
rect 10945 18785 10957 18788
rect 11020 18816 11026 18828
rect 11020 18788 11093 18816
rect 10945 18779 10968 18785
rect 10962 18776 10968 18779
rect 11020 18776 11026 18788
rect 13998 18776 14004 18828
rect 14056 18776 14062 18828
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 15841 18819 15899 18825
rect 15841 18816 15853 18819
rect 15344 18788 15853 18816
rect 15344 18776 15350 18788
rect 15841 18785 15853 18788
rect 15887 18816 15899 18819
rect 16574 18816 16580 18828
rect 15887 18788 16580 18816
rect 15887 18785 15899 18788
rect 15841 18779 15899 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 17396 18819 17454 18825
rect 17396 18785 17408 18819
rect 17442 18816 17454 18819
rect 17678 18816 17684 18828
rect 17442 18788 17684 18816
rect 17442 18785 17454 18788
rect 17396 18779 17454 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18816 19211 18819
rect 19242 18816 19248 18828
rect 19199 18788 19248 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19794 18816 19800 18828
rect 19755 18788 19800 18816
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 22554 18776 22560 18828
rect 22612 18776 22618 18828
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23474 18816 23480 18828
rect 23072 18788 23480 18816
rect 23072 18776 23078 18788
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 10652 18720 10701 18748
rect 10652 18708 10658 18720
rect 10689 18717 10701 18720
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14182 18748 14188 18760
rect 13872 18720 14188 18748
rect 13872 18708 13878 18720
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 16022 18748 16028 18760
rect 15983 18720 16028 18748
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 17126 18748 17132 18760
rect 16172 18720 17132 18748
rect 16172 18708 16178 18720
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 21450 18748 21456 18760
rect 21232 18720 21456 18748
rect 21232 18708 21238 18720
rect 21450 18708 21456 18720
rect 21508 18748 21514 18760
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 21508 18720 21649 18748
rect 21508 18708 21514 18720
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18748 21787 18751
rect 22738 18748 22744 18760
rect 21775 18720 22744 18748
rect 21775 18717 21787 18720
rect 21729 18711 21787 18717
rect 20990 18640 20996 18692
rect 21048 18680 21054 18692
rect 21744 18680 21772 18711
rect 22738 18708 22744 18720
rect 22796 18708 22802 18760
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 23382 18748 23388 18760
rect 22879 18720 23388 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 23842 18748 23848 18760
rect 23803 18720 23848 18748
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 21048 18652 21772 18680
rect 21048 18640 21054 18652
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18612 10471 18615
rect 10870 18612 10876 18624
rect 10459 18584 10876 18612
rect 10459 18581 10471 18584
rect 10413 18575 10471 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11422 18572 11428 18624
rect 11480 18612 11486 18624
rect 12069 18615 12127 18621
rect 12069 18612 12081 18615
rect 11480 18584 12081 18612
rect 11480 18572 11486 18584
rect 12069 18581 12081 18584
rect 12115 18581 12127 18615
rect 12069 18575 12127 18581
rect 14826 18572 14832 18624
rect 14884 18612 14890 18624
rect 15013 18615 15071 18621
rect 15013 18612 15025 18615
rect 14884 18584 15025 18612
rect 14884 18572 14890 18584
rect 15013 18581 15025 18584
rect 15059 18581 15071 18615
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 15013 18575 15071 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 22186 18612 22192 18624
rect 22147 18584 22192 18612
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 25222 18612 25228 18624
rect 25183 18584 25228 18612
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10594 18408 10600 18420
rect 10555 18380 10600 18408
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 13906 18368 13912 18420
rect 13964 18408 13970 18420
rect 14185 18411 14243 18417
rect 14185 18408 14197 18411
rect 13964 18380 14197 18408
rect 13964 18368 13970 18380
rect 14185 18377 14197 18380
rect 14231 18377 14243 18411
rect 14185 18371 14243 18377
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 14700 18380 15761 18408
rect 14700 18368 14706 18380
rect 15749 18377 15761 18380
rect 15795 18408 15807 18411
rect 15838 18408 15844 18420
rect 15795 18380 15844 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16393 18411 16451 18417
rect 16393 18408 16405 18411
rect 16080 18380 16405 18408
rect 16080 18368 16086 18380
rect 16393 18377 16405 18380
rect 16439 18408 16451 18411
rect 16850 18408 16856 18420
rect 16439 18380 16856 18408
rect 16439 18377 16451 18380
rect 16393 18371 16451 18377
rect 16850 18368 16856 18380
rect 16908 18408 16914 18420
rect 17678 18408 17684 18420
rect 16908 18380 17684 18408
rect 16908 18368 16914 18380
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 20438 18408 20444 18420
rect 20395 18380 20444 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 22833 18411 22891 18417
rect 22833 18408 22845 18411
rect 22796 18380 22845 18408
rect 22796 18368 22802 18380
rect 22833 18377 22845 18380
rect 22879 18377 22891 18411
rect 22833 18371 22891 18377
rect 23198 18368 23204 18420
rect 23256 18408 23262 18420
rect 23385 18411 23443 18417
rect 23385 18408 23397 18411
rect 23256 18380 23397 18408
rect 23256 18368 23262 18380
rect 23385 18377 23397 18380
rect 23431 18377 23443 18411
rect 23385 18371 23443 18377
rect 11793 18343 11851 18349
rect 11793 18340 11805 18343
rect 11256 18312 11805 18340
rect 10686 18232 10692 18284
rect 10744 18272 10750 18284
rect 11256 18281 11284 18312
rect 11793 18309 11805 18312
rect 11839 18309 11851 18343
rect 11793 18303 11851 18309
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 16669 18343 16727 18349
rect 16669 18340 16681 18343
rect 16632 18312 16681 18340
rect 16632 18300 16638 18312
rect 16669 18309 16681 18312
rect 16715 18309 16727 18343
rect 16669 18303 16727 18309
rect 17126 18300 17132 18352
rect 17184 18340 17190 18352
rect 17313 18343 17371 18349
rect 17313 18340 17325 18343
rect 17184 18312 17325 18340
rect 17184 18300 17190 18312
rect 17313 18309 17325 18312
rect 17359 18340 17371 18343
rect 18785 18343 18843 18349
rect 18785 18340 18797 18343
rect 17359 18312 18797 18340
rect 17359 18309 17371 18312
rect 17313 18303 17371 18309
rect 18785 18309 18797 18312
rect 18831 18340 18843 18343
rect 18831 18312 19012 18340
rect 18831 18309 18843 18312
rect 18785 18303 18843 18309
rect 11241 18275 11299 18281
rect 11241 18272 11253 18275
rect 10744 18244 11253 18272
rect 10744 18232 10750 18244
rect 11241 18241 11253 18244
rect 11287 18241 11299 18275
rect 11422 18272 11428 18284
rect 11383 18244 11428 18272
rect 11241 18235 11299 18241
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18272 12311 18275
rect 13357 18275 13415 18281
rect 13357 18272 13369 18275
rect 12299 18244 13369 18272
rect 12299 18241 12311 18244
rect 12253 18235 12311 18241
rect 13357 18241 13369 18244
rect 13403 18272 13415 18275
rect 13630 18272 13636 18284
rect 13403 18244 13636 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 13998 18272 14004 18284
rect 13955 18244 14004 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 18984 18281 19012 18312
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22465 18275 22523 18281
rect 22465 18272 22477 18275
rect 22152 18244 22477 18272
rect 22152 18232 22158 18244
rect 22465 18241 22477 18244
rect 22511 18241 22523 18275
rect 23400 18272 23428 18371
rect 23842 18368 23848 18420
rect 23900 18408 23906 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 23900 18380 24685 18408
rect 23900 18368 23906 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 24673 18371 24731 18377
rect 25133 18411 25191 18417
rect 25133 18377 25145 18411
rect 25179 18408 25191 18411
rect 25222 18408 25228 18420
rect 25179 18380 25228 18408
rect 25179 18377 25191 18380
rect 25133 18371 25191 18377
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 23400 18244 24133 18272
rect 22465 18235 22523 18241
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18272 24363 18275
rect 24670 18272 24676 18284
rect 24351 18244 24676 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 24670 18232 24676 18244
rect 24728 18272 24734 18284
rect 25148 18272 25176 18371
rect 25222 18368 25228 18380
rect 25280 18368 25286 18420
rect 24728 18244 25176 18272
rect 24728 18232 24734 18244
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 11440 18204 11468 18232
rect 9999 18176 11468 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 12860 18176 13185 18204
rect 12860 18164 12866 18176
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 14366 18204 14372 18216
rect 14327 18176 14372 18204
rect 13173 18167 13231 18173
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 16632 18176 16865 18204
rect 16632 18164 16638 18176
rect 16853 18173 16865 18176
rect 16899 18204 16911 18207
rect 18233 18207 18291 18213
rect 18233 18204 18245 18207
rect 16899 18176 18245 18204
rect 16899 18173 16911 18176
rect 16853 18167 16911 18173
rect 18233 18173 18245 18176
rect 18279 18173 18291 18207
rect 21174 18204 21180 18216
rect 21135 18176 21180 18204
rect 18233 18167 18291 18173
rect 21174 18164 21180 18176
rect 21232 18164 21238 18216
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23716 18176 24041 18204
rect 23716 18164 23722 18176
rect 24029 18173 24041 18176
rect 24075 18173 24087 18207
rect 25222 18204 25228 18216
rect 25183 18176 25228 18204
rect 24029 18167 24087 18173
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25280 18176 25789 18204
rect 25280 18164 25286 18176
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 12434 18096 12440 18148
rect 12492 18136 12498 18148
rect 12713 18139 12771 18145
rect 12713 18136 12725 18139
rect 12492 18108 12725 18136
rect 12492 18096 12498 18108
rect 12713 18105 12725 18108
rect 12759 18136 12771 18139
rect 13262 18136 13268 18148
rect 12759 18108 13268 18136
rect 12759 18105 12771 18108
rect 12713 18099 12771 18105
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 14614 18139 14672 18145
rect 14614 18136 14626 18139
rect 14240 18108 14626 18136
rect 14240 18096 14246 18108
rect 14614 18105 14626 18108
rect 14660 18136 14672 18139
rect 14826 18136 14832 18148
rect 14660 18108 14832 18136
rect 14660 18105 14672 18108
rect 14614 18099 14672 18105
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 19058 18096 19064 18148
rect 19116 18136 19122 18148
rect 19214 18139 19272 18145
rect 19214 18136 19226 18139
rect 19116 18108 19226 18136
rect 19116 18096 19122 18108
rect 19214 18105 19226 18108
rect 19260 18105 19272 18139
rect 19214 18099 19272 18105
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 21913 18139 21971 18145
rect 21913 18136 21925 18139
rect 20772 18108 21925 18136
rect 20772 18096 20778 18108
rect 21913 18105 21925 18108
rect 21959 18136 21971 18139
rect 22186 18136 22192 18148
rect 21959 18108 22192 18136
rect 21959 18105 21971 18108
rect 21913 18099 21971 18105
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 23198 18096 23204 18148
rect 23256 18136 23262 18148
rect 23566 18136 23572 18148
rect 23256 18108 23572 18136
rect 23256 18096 23262 18108
rect 23566 18096 23572 18108
rect 23624 18096 23630 18148
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18068 10839 18071
rect 10962 18068 10968 18080
rect 10827 18040 10968 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11146 18068 11152 18080
rect 11107 18040 11152 18068
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 17218 18068 17224 18080
rect 17083 18040 17224 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 21450 18068 21456 18080
rect 21411 18040 21456 18068
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 21818 18068 21824 18080
rect 21779 18040 21824 18068
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 23658 18068 23664 18080
rect 23619 18040 23664 18068
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 25406 18068 25412 18080
rect 25367 18040 25412 18068
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 13722 17864 13728 17876
rect 13683 17836 13728 17864
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 15746 17864 15752 17876
rect 15707 17836 15752 17864
rect 15746 17824 15752 17836
rect 15804 17864 15810 17876
rect 16301 17867 16359 17873
rect 16301 17864 16313 17867
rect 15804 17836 16313 17864
rect 15804 17824 15810 17836
rect 16301 17833 16313 17836
rect 16347 17833 16359 17867
rect 16301 17827 16359 17833
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20070 17864 20076 17876
rect 20027 17836 20076 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 20346 17864 20352 17876
rect 20307 17836 20352 17864
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 21542 17824 21548 17876
rect 21600 17864 21606 17876
rect 21913 17867 21971 17873
rect 21913 17864 21925 17867
rect 21600 17836 21925 17864
rect 21600 17824 21606 17836
rect 21913 17833 21925 17836
rect 21959 17833 21971 17867
rect 21913 17827 21971 17833
rect 23109 17867 23167 17873
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 23658 17864 23664 17876
rect 23155 17836 23664 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 24210 17864 24216 17876
rect 24171 17836 24216 17864
rect 24210 17824 24216 17836
rect 24268 17824 24274 17876
rect 11422 17756 11428 17808
rect 11480 17805 11486 17808
rect 11480 17799 11544 17805
rect 11480 17765 11498 17799
rect 11532 17765 11544 17799
rect 11480 17759 11544 17765
rect 11480 17756 11486 17759
rect 14550 17756 14556 17808
rect 14608 17796 14614 17808
rect 15654 17796 15660 17808
rect 14608 17768 15660 17796
rect 14608 17756 14614 17768
rect 15654 17756 15660 17768
rect 15712 17756 15718 17808
rect 17212 17799 17270 17805
rect 17212 17765 17224 17799
rect 17258 17796 17270 17799
rect 17402 17796 17408 17808
rect 17258 17768 17408 17796
rect 17258 17765 17270 17768
rect 17212 17759 17270 17765
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 21361 17799 21419 17805
rect 21361 17765 21373 17799
rect 21407 17796 21419 17799
rect 22462 17796 22468 17808
rect 21407 17768 22468 17796
rect 21407 17765 21419 17768
rect 21361 17759 21419 17765
rect 22462 17756 22468 17768
rect 22520 17796 22526 17808
rect 23198 17796 23204 17808
rect 22520 17768 23204 17796
rect 22520 17756 22526 17768
rect 23198 17756 23204 17768
rect 23256 17756 23262 17808
rect 23290 17756 23296 17808
rect 23348 17796 23354 17808
rect 23348 17768 24808 17796
rect 23348 17756 23354 17768
rect 10686 17688 10692 17740
rect 10744 17728 10750 17740
rect 11241 17731 11299 17737
rect 11241 17728 11253 17731
rect 10744 17700 11253 17728
rect 10744 17688 10750 17700
rect 11241 17697 11253 17700
rect 11287 17728 11299 17731
rect 11790 17728 11796 17740
rect 11287 17700 11796 17728
rect 11287 17697 11299 17700
rect 11241 17691 11299 17697
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 17034 17728 17040 17740
rect 16991 17700 17040 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 19794 17728 19800 17740
rect 19755 17700 19800 17728
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 20772 17700 21281 17728
rect 20772 17688 20778 17700
rect 21269 17697 21281 17700
rect 21315 17697 21327 17731
rect 23566 17728 23572 17740
rect 23527 17700 23572 17728
rect 21269 17691 21327 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 24780 17737 24808 17768
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17728 24823 17731
rect 25590 17728 25596 17740
rect 24811 17700 25596 17728
rect 24811 17697 24823 17700
rect 24765 17691 24823 17697
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 10870 17660 10876 17672
rect 10831 17632 10876 17660
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17660 14243 17663
rect 14550 17660 14556 17672
rect 14231 17632 14556 17660
rect 14231 17629 14243 17632
rect 14185 17623 14243 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17660 21603 17663
rect 21634 17660 21640 17672
rect 21591 17632 21640 17660
rect 21591 17629 21603 17632
rect 21545 17623 21603 17629
rect 15013 17595 15071 17601
rect 15013 17592 15025 17595
rect 14200 17564 15025 17592
rect 14200 17536 14228 17564
rect 15013 17561 15025 17564
rect 15059 17592 15071 17595
rect 15856 17592 15884 17623
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23753 17663 23811 17669
rect 23753 17660 23765 17663
rect 23348 17632 23765 17660
rect 23348 17620 23354 17632
rect 23753 17629 23765 17632
rect 23799 17629 23811 17663
rect 23753 17623 23811 17629
rect 16022 17592 16028 17604
rect 15059 17564 16028 17592
rect 15059 17561 15071 17564
rect 15013 17555 15071 17561
rect 16022 17552 16028 17564
rect 16080 17552 16086 17604
rect 20901 17595 20959 17601
rect 20901 17561 20913 17595
rect 20947 17592 20959 17595
rect 22186 17592 22192 17604
rect 20947 17564 22192 17592
rect 20947 17561 20959 17564
rect 20901 17555 20959 17561
rect 22186 17552 22192 17564
rect 22244 17552 22250 17604
rect 23198 17592 23204 17604
rect 23159 17564 23204 17592
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 23934 17552 23940 17604
rect 23992 17592 23998 17604
rect 24578 17592 24584 17604
rect 23992 17564 24584 17592
rect 23992 17552 23998 17564
rect 24578 17552 24584 17564
rect 24636 17552 24642 17604
rect 12621 17527 12679 17533
rect 12621 17493 12633 17527
rect 12667 17524 12679 17527
rect 12710 17524 12716 17536
rect 12667 17496 12716 17524
rect 12667 17493 12679 17496
rect 12621 17487 12679 17493
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 14182 17484 14188 17536
rect 14240 17484 14246 17536
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 14737 17527 14795 17533
rect 14737 17524 14749 17527
rect 14424 17496 14749 17524
rect 14424 17484 14430 17496
rect 14737 17493 14749 17496
rect 14783 17524 14795 17527
rect 14826 17524 14832 17536
rect 14783 17496 14832 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 15289 17527 15347 17533
rect 15289 17493 15301 17527
rect 15335 17524 15347 17527
rect 15378 17524 15384 17536
rect 15335 17496 15384 17524
rect 15335 17493 15347 17496
rect 15289 17487 15347 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 18322 17524 18328 17536
rect 18283 17496 18328 17524
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 19058 17524 19064 17536
rect 19019 17496 19064 17524
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 22278 17524 22284 17536
rect 22239 17496 22284 17524
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 24946 17524 24952 17536
rect 24907 17496 24952 17524
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17320 11854 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 11848 17292 12173 17320
rect 11848 17280 11854 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 13814 17320 13820 17332
rect 13775 17292 13820 17320
rect 12161 17283 12219 17289
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 11238 17184 11244 17196
rect 10367 17156 11244 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 11238 17144 11244 17156
rect 11296 17184 11302 17196
rect 11422 17184 11428 17196
rect 11296 17156 11428 17184
rect 11296 17144 11302 17156
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 12176 17116 12204 17283
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14461 17323 14519 17329
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 14642 17320 14648 17332
rect 14507 17292 14648 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 16022 17280 16028 17332
rect 16080 17320 16086 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 16080 17292 16313 17320
rect 16080 17280 16086 17292
rect 16301 17289 16313 17292
rect 16347 17289 16359 17323
rect 17034 17320 17040 17332
rect 16995 17292 17040 17320
rect 16301 17283 16359 17289
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 17402 17320 17408 17332
rect 17363 17292 17408 17320
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 20496 17292 20545 17320
rect 20496 17280 20502 17292
rect 20533 17289 20545 17292
rect 20579 17320 20591 17323
rect 20990 17320 20996 17332
rect 20579 17292 20996 17320
rect 20579 17289 20591 17292
rect 20533 17283 20591 17289
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 21085 17323 21143 17329
rect 21085 17289 21097 17323
rect 21131 17320 21143 17323
rect 21818 17320 21824 17332
rect 21131 17292 21824 17320
rect 21131 17289 21143 17292
rect 21085 17283 21143 17289
rect 21818 17280 21824 17292
rect 21876 17320 21882 17332
rect 22278 17320 22284 17332
rect 21876 17292 22284 17320
rect 21876 17280 21882 17292
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 22462 17320 22468 17332
rect 22423 17292 22468 17320
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 23348 17292 25053 17320
rect 23348 17280 23354 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25590 17320 25596 17332
rect 25551 17292 25596 17320
rect 25041 17283 25099 17289
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 13832 17184 13860 17280
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 16390 17252 16396 17264
rect 16172 17224 16396 17252
rect 16172 17212 16178 17224
rect 16390 17212 16396 17224
rect 16448 17212 16454 17264
rect 17052 17252 17080 17280
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 17052 17224 18429 17252
rect 18417 17221 18429 17224
rect 18463 17252 18475 17255
rect 18463 17224 18644 17252
rect 18463 17221 18475 17224
rect 18417 17215 18475 17221
rect 18616 17193 18644 17224
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 23385 17255 23443 17261
rect 23385 17252 23397 17255
rect 20956 17224 23397 17252
rect 20956 17212 20962 17224
rect 23385 17221 23397 17224
rect 23431 17252 23443 17255
rect 23431 17224 23704 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 18601 17187 18659 17193
rect 13832 17156 15056 17184
rect 15028 17128 15056 17156
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 20993 17187 21051 17193
rect 20993 17184 21005 17187
rect 20772 17156 21005 17184
rect 20772 17144 20778 17156
rect 20993 17153 21005 17156
rect 21039 17153 21051 17187
rect 21634 17184 21640 17196
rect 21595 17156 21640 17184
rect 20993 17147 21051 17153
rect 21634 17144 21640 17156
rect 21692 17184 21698 17196
rect 23676 17193 23704 17224
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 21692 17156 22845 17184
rect 21692 17144 21698 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 12710 17125 12716 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 10735 17088 11468 17116
rect 12176 17088 12449 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 11149 17051 11207 17057
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 11330 17048 11336 17060
rect 11195 17020 11336 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 11440 16992 11468 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12704 17116 12716 17125
rect 12671 17088 12716 17116
rect 12437 17079 12495 17085
rect 12704 17079 12716 17088
rect 12452 17048 12480 17079
rect 12710 17076 12716 17079
rect 12768 17076 12774 17128
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 14826 17048 14832 17060
rect 12452 17020 14832 17048
rect 14826 17008 14832 17020
rect 14884 17048 14890 17060
rect 14936 17048 14964 17079
rect 15010 17076 15016 17128
rect 15068 17116 15074 17128
rect 15177 17119 15235 17125
rect 15177 17116 15189 17119
rect 15068 17088 15189 17116
rect 15068 17076 15074 17088
rect 15177 17085 15189 17088
rect 15223 17085 15235 17119
rect 15177 17079 15235 17085
rect 20806 17076 20812 17128
rect 20864 17116 20870 17128
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20864 17088 21465 17116
rect 20864 17076 20870 17088
rect 21453 17085 21465 17088
rect 21499 17116 21511 17119
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21499 17088 21925 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 22094 17076 22100 17128
rect 22152 17076 22158 17128
rect 23928 17119 23986 17125
rect 23928 17085 23940 17119
rect 23974 17116 23986 17119
rect 24670 17116 24676 17128
rect 23974 17088 24676 17116
rect 23974 17085 23986 17088
rect 23928 17079 23986 17085
rect 24670 17076 24676 17088
rect 24728 17076 24734 17128
rect 16942 17048 16948 17060
rect 14884 17020 16948 17048
rect 14884 17008 14890 17020
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 18874 17057 18880 17060
rect 18868 17048 18880 17057
rect 18787 17020 18880 17048
rect 18868 17011 18880 17020
rect 18932 17048 18938 17060
rect 22112 17048 22140 17076
rect 18932 17020 22140 17048
rect 18874 17008 18880 17011
rect 18932 17008 18938 17020
rect 10781 16983 10839 16989
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 11054 16980 11060 16992
rect 10827 16952 11060 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11422 16980 11428 16992
rect 11287 16952 11428 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 14274 16980 14280 16992
rect 13596 16952 14280 16980
rect 13596 16940 13602 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 19058 16940 19064 16992
rect 19116 16980 19122 16992
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 19116 16952 19993 16980
rect 19116 16940 19122 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 20990 16940 20996 16992
rect 21048 16980 21054 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 21048 16952 21557 16980
rect 21048 16940 21054 16952
rect 21545 16949 21557 16952
rect 21591 16949 21603 16983
rect 21545 16943 21603 16949
rect 21913 16983 21971 16989
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 22097 16983 22155 16989
rect 22097 16980 22109 16983
rect 21959 16952 22109 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22097 16949 22109 16952
rect 22143 16949 22155 16983
rect 22097 16943 22155 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 11238 16776 11244 16788
rect 11199 16748 11244 16776
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 11333 16779 11391 16785
rect 11333 16745 11345 16779
rect 11379 16776 11391 16779
rect 12434 16776 12440 16788
rect 11379 16748 12440 16776
rect 11379 16745 11391 16748
rect 11333 16739 11391 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 12710 16776 12716 16788
rect 12575 16748 12716 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 11054 16668 11060 16720
rect 11112 16708 11118 16720
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 11112 16680 11713 16708
rect 11112 16668 11118 16680
rect 11701 16677 11713 16680
rect 11747 16677 11759 16711
rect 11701 16671 11759 16677
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11330 16640 11336 16652
rect 10919 16612 11336 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 12544 16640 12572 16739
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 14366 16776 14372 16788
rect 14327 16748 14372 16776
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 15010 16776 15016 16788
rect 14971 16748 15016 16776
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16745 15347 16779
rect 15289 16739 15347 16745
rect 12268 16612 12572 16640
rect 14185 16643 14243 16649
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11790 16572 11796 16584
rect 11204 16544 11796 16572
rect 11204 16532 11210 16544
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11940 16544 11989 16572
rect 11940 16532 11946 16544
rect 11977 16541 11989 16544
rect 12023 16572 12035 16575
rect 12268 16572 12296 16612
rect 14185 16609 14197 16643
rect 14231 16640 14243 16643
rect 14274 16640 14280 16652
rect 14231 16612 14280 16640
rect 14231 16609 14243 16612
rect 14185 16603 14243 16609
rect 14274 16600 14280 16612
rect 14332 16640 14338 16652
rect 15304 16640 15332 16739
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 18874 16776 18880 16788
rect 18835 16748 18880 16776
rect 16393 16739 16451 16745
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 22152 16748 22293 16776
rect 22152 16736 22158 16748
rect 22281 16745 22293 16748
rect 22327 16776 22339 16779
rect 22370 16776 22376 16788
rect 22327 16748 22376 16776
rect 22327 16745 22339 16748
rect 22281 16739 22339 16745
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 22925 16779 22983 16785
rect 22925 16745 22937 16779
rect 22971 16776 22983 16779
rect 23385 16779 23443 16785
rect 23385 16776 23397 16779
rect 22971 16748 23397 16776
rect 22971 16745 22983 16748
rect 22925 16739 22983 16745
rect 23385 16745 23397 16748
rect 23431 16776 23443 16779
rect 23566 16776 23572 16788
rect 23431 16748 23572 16776
rect 23431 16745 23443 16748
rect 23385 16739 23443 16745
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 24489 16779 24547 16785
rect 24489 16745 24501 16779
rect 24535 16776 24547 16779
rect 24670 16776 24676 16788
rect 24535 16748 24676 16776
rect 24535 16745 24547 16748
rect 24489 16739 24547 16745
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 17126 16717 17132 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15436 16680 15761 16708
rect 15436 16668 15442 16680
rect 15749 16677 15761 16680
rect 15795 16677 15807 16711
rect 15749 16671 15807 16677
rect 17120 16671 17132 16717
rect 17184 16708 17190 16720
rect 18322 16708 18328 16720
rect 17184 16680 18328 16708
rect 17126 16668 17132 16671
rect 17184 16668 17190 16680
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 23198 16708 23204 16720
rect 23159 16680 23204 16708
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 23474 16668 23480 16720
rect 23532 16708 23538 16720
rect 23753 16711 23811 16717
rect 23753 16708 23765 16711
rect 23532 16680 23765 16708
rect 23532 16668 23538 16680
rect 23753 16677 23765 16680
rect 23799 16677 23811 16711
rect 23753 16671 23811 16677
rect 14332 16612 15332 16640
rect 14332 16600 14338 16612
rect 12023 16544 12296 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 14826 16532 14832 16584
rect 14884 16572 14890 16584
rect 15396 16572 15424 16668
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 14884 16544 15424 16572
rect 15488 16612 15669 16640
rect 14884 16532 14890 16544
rect 14642 16464 14648 16516
rect 14700 16504 14706 16516
rect 15488 16504 15516 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 16942 16640 16948 16652
rect 16899 16612 16948 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16640 19855 16643
rect 20622 16640 20628 16652
rect 19843 16612 20628 16640
rect 19843 16609 19855 16612
rect 19797 16603 19855 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 21157 16643 21215 16649
rect 21157 16640 21169 16643
rect 20824 16612 21169 16640
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 20824 16504 20852 16612
rect 21157 16609 21169 16612
rect 21203 16640 21215 16643
rect 21634 16640 21640 16652
rect 21203 16612 21640 16640
rect 21203 16609 21215 16612
rect 21157 16603 21215 16609
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 20898 16532 20904 16584
rect 20956 16572 20962 16584
rect 23842 16572 23848 16584
rect 20956 16544 21001 16572
rect 23803 16544 23848 16572
rect 20956 16532 20962 16544
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 24029 16575 24087 16581
rect 24029 16541 24041 16575
rect 24075 16572 24087 16575
rect 24210 16572 24216 16584
rect 24075 16544 24216 16572
rect 24075 16541 24087 16544
rect 24029 16535 24087 16541
rect 24210 16532 24216 16544
rect 24268 16572 24274 16584
rect 24504 16572 24532 16739
rect 24670 16736 24676 16748
rect 24728 16736 24734 16788
rect 25130 16776 25136 16788
rect 25091 16748 25136 16776
rect 25130 16736 25136 16748
rect 25188 16736 25194 16788
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 24949 16643 25007 16649
rect 24949 16640 24961 16643
rect 24912 16612 24961 16640
rect 24912 16600 24918 16612
rect 24949 16609 24961 16612
rect 24995 16609 25007 16643
rect 24949 16603 25007 16609
rect 24268 16544 24532 16572
rect 24268 16532 24274 16544
rect 14700 16476 15516 16504
rect 20640 16476 20852 16504
rect 14700 16464 14706 16476
rect 18230 16436 18236 16448
rect 18191 16408 18236 16436
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 20640 16445 20668 16476
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20496 16408 20637 16436
rect 20496 16396 20502 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20625 16399 20683 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 11112 16204 11161 16232
rect 11112 16192 11118 16204
rect 11149 16201 11161 16204
rect 11195 16201 11207 16235
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11149 16195 11207 16201
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 13817 16235 13875 16241
rect 13817 16201 13829 16235
rect 13863 16232 13875 16235
rect 14642 16232 14648 16244
rect 13863 16204 14648 16232
rect 13863 16201 13875 16204
rect 13817 16195 13875 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 15838 16232 15844 16244
rect 15795 16204 15844 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 16080 16204 16221 16232
rect 16080 16192 16086 16204
rect 16209 16201 16221 16204
rect 16255 16201 16267 16235
rect 16209 16195 16267 16201
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 11848 16136 12173 16164
rect 11848 16124 11854 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12161 16127 12219 16133
rect 11330 16096 11336 16108
rect 11291 16068 11336 16096
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 14182 16096 14188 16108
rect 14095 16068 14188 16096
rect 14182 16056 14188 16068
rect 14240 16096 14246 16108
rect 15197 16099 15255 16105
rect 15197 16096 15209 16099
rect 14240 16068 15209 16096
rect 14240 16056 14246 16068
rect 15197 16065 15209 16068
rect 15243 16065 15255 16099
rect 16224 16096 16252 16195
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 17126 16232 17132 16244
rect 17000 16204 17132 16232
rect 17000 16192 17006 16204
rect 17126 16192 17132 16204
rect 17184 16232 17190 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 17184 16204 17417 16232
rect 17184 16192 17190 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16232 20223 16235
rect 20530 16232 20536 16244
rect 20211 16204 20536 16232
rect 20211 16201 20223 16204
rect 20165 16195 20223 16201
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 21545 16235 21603 16241
rect 21545 16232 21557 16235
rect 20772 16204 21557 16232
rect 20772 16192 20778 16204
rect 21545 16201 21557 16204
rect 21591 16232 21603 16235
rect 21591 16204 22140 16232
rect 21591 16201 21603 16204
rect 21545 16195 21603 16201
rect 20898 16124 20904 16176
rect 20956 16164 20962 16176
rect 21177 16167 21235 16173
rect 21177 16164 21189 16167
rect 20956 16136 21189 16164
rect 20956 16124 20962 16136
rect 21177 16133 21189 16136
rect 21223 16133 21235 16167
rect 21177 16127 21235 16133
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16224 16068 16865 16096
rect 15197 16059 15255 16065
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 17034 16096 17040 16108
rect 16995 16068 17040 16096
rect 16853 16059 16911 16065
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12492 16000 12909 16028
rect 12492 15988 12498 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 15102 16028 15108 16040
rect 15063 16000 15108 16028
rect 12897 15991 12955 15997
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16761 16031 16819 16037
rect 16761 16028 16773 16031
rect 16356 16000 16773 16028
rect 16356 15988 16362 16000
rect 16761 15997 16773 16000
rect 16807 15997 16819 16031
rect 16868 16028 16896 16059
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 19058 16096 19064 16108
rect 18555 16068 19064 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 19058 16056 19064 16068
rect 19116 16096 19122 16108
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 19116 16068 19165 16096
rect 19116 16056 19122 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19153 16059 19211 16065
rect 19705 16099 19763 16105
rect 19705 16065 19717 16099
rect 19751 16096 19763 16099
rect 20438 16096 20444 16108
rect 19751 16068 20444 16096
rect 19751 16065 19763 16068
rect 19705 16059 19763 16065
rect 20438 16056 20444 16068
rect 20496 16096 20502 16108
rect 20717 16099 20775 16105
rect 20717 16096 20729 16099
rect 20496 16068 20729 16096
rect 20496 16056 20502 16068
rect 20717 16065 20729 16068
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 16942 16028 16948 16040
rect 16868 16000 16948 16028
rect 16761 15991 16819 15997
rect 13630 15920 13636 15972
rect 13688 15960 13694 15972
rect 14461 15963 14519 15969
rect 14461 15960 14473 15963
rect 13688 15932 14473 15960
rect 13688 15920 13694 15932
rect 14461 15929 14473 15932
rect 14507 15960 14519 15963
rect 15120 15960 15148 15988
rect 14507 15932 15148 15960
rect 16776 15960 16804 15991
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 20070 16028 20076 16040
rect 17052 16000 20076 16028
rect 17052 15960 17080 16000
rect 20070 15988 20076 16000
rect 20128 16028 20134 16040
rect 22112 16037 22140 16204
rect 23474 16192 23480 16244
rect 23532 16232 23538 16244
rect 23845 16235 23903 16241
rect 23845 16232 23857 16235
rect 23532 16204 23857 16232
rect 23532 16192 23538 16204
rect 23845 16201 23857 16204
rect 23891 16201 23903 16235
rect 24210 16232 24216 16244
rect 24171 16204 24216 16232
rect 23845 16195 23903 16201
rect 24210 16192 24216 16204
rect 24268 16192 24274 16244
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25501 16235 25559 16241
rect 25501 16232 25513 16235
rect 24912 16204 25513 16232
rect 24912 16192 24918 16204
rect 25501 16201 25513 16204
rect 25547 16201 25559 16235
rect 25501 16195 25559 16201
rect 22186 16056 22192 16108
rect 22244 16096 22250 16108
rect 22370 16096 22376 16108
rect 22244 16068 22289 16096
rect 22331 16068 22376 16096
rect 22244 16056 22250 16068
rect 22370 16056 22376 16068
rect 22428 16096 22434 16108
rect 22741 16099 22799 16105
rect 22741 16096 22753 16099
rect 22428 16068 22753 16096
rect 22428 16056 22434 16068
rect 22741 16065 22753 16068
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 24210 16056 24216 16108
rect 24268 16096 24274 16108
rect 25038 16096 25044 16108
rect 24268 16068 25044 16096
rect 24268 16056 24274 16068
rect 25038 16056 25044 16068
rect 25096 16056 25102 16108
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20128 16000 20545 16028
rect 20128 15988 20134 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 22097 16031 22155 16037
rect 22097 15997 22109 16031
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 24118 15988 24124 16040
rect 24176 16028 24182 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24176 16000 24593 16028
rect 24176 15988 24182 16000
rect 24581 15997 24593 16000
rect 24627 16028 24639 16031
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24627 16000 25145 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 16776 15932 17080 15960
rect 17865 15963 17923 15969
rect 14507 15929 14519 15932
rect 14461 15923 14519 15929
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18969 15963 19027 15969
rect 17911 15932 18920 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 12621 15895 12679 15901
rect 12621 15861 12633 15895
rect 12667 15892 12679 15895
rect 13722 15892 13728 15904
rect 12667 15864 13728 15892
rect 12667 15861 12679 15864
rect 12621 15855 12679 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 14608 15864 15025 15892
rect 14608 15852 14614 15864
rect 15013 15861 15025 15864
rect 15059 15861 15071 15895
rect 16390 15892 16396 15904
rect 16351 15864 16396 15892
rect 15013 15855 15071 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 18598 15892 18604 15904
rect 18559 15864 18604 15892
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 18892 15892 18920 15932
rect 18969 15929 18981 15963
rect 19015 15960 19027 15963
rect 19150 15960 19156 15972
rect 19015 15932 19156 15960
rect 19015 15929 19027 15932
rect 18969 15923 19027 15929
rect 19150 15920 19156 15932
rect 19208 15960 19214 15972
rect 19208 15932 21772 15960
rect 19208 15920 19214 15932
rect 19058 15892 19064 15904
rect 18892 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 19518 15852 19524 15904
rect 19576 15892 19582 15904
rect 21744 15901 21772 15932
rect 19981 15895 20039 15901
rect 19981 15892 19993 15895
rect 19576 15864 19993 15892
rect 19576 15852 19582 15864
rect 19981 15861 19993 15864
rect 20027 15892 20039 15895
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 20027 15864 20637 15892
rect 20027 15861 20039 15864
rect 19981 15855 20039 15861
rect 20625 15861 20637 15864
rect 20671 15861 20683 15895
rect 20625 15855 20683 15861
rect 21729 15895 21787 15901
rect 21729 15861 21741 15895
rect 21775 15861 21787 15895
rect 21729 15855 21787 15861
rect 23014 15852 23020 15904
rect 23072 15892 23078 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 23072 15864 23397 15892
rect 23072 15852 23078 15864
rect 23385 15861 23397 15864
rect 23431 15892 23443 15895
rect 23842 15892 23848 15904
rect 23431 15864 23848 15892
rect 23431 15861 23443 15864
rect 23385 15855 23443 15861
rect 23842 15852 23848 15864
rect 23900 15852 23906 15904
rect 24762 15892 24768 15904
rect 24723 15864 24768 15892
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 14274 15688 14280 15700
rect 14235 15660 14280 15688
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14608 15660 14657 15688
rect 14608 15648 14614 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 14884 15660 15025 15688
rect 14884 15648 14890 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15013 15651 15071 15657
rect 16669 15691 16727 15697
rect 16669 15657 16681 15691
rect 16715 15688 16727 15691
rect 17034 15688 17040 15700
rect 16715 15660 17040 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 19150 15688 19156 15700
rect 19111 15660 19156 15688
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 20070 15648 20076 15700
rect 20128 15688 20134 15700
rect 20165 15691 20223 15697
rect 20165 15688 20177 15691
rect 20128 15660 20177 15688
rect 20128 15648 20134 15660
rect 20165 15657 20177 15660
rect 20211 15657 20223 15691
rect 20165 15651 20223 15657
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 21085 15691 21143 15697
rect 21085 15688 21097 15691
rect 20496 15660 21097 15688
rect 20496 15648 20502 15660
rect 21085 15657 21097 15660
rect 21131 15688 21143 15691
rect 22741 15691 22799 15697
rect 22741 15688 22753 15691
rect 21131 15660 22753 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 22741 15657 22753 15660
rect 22787 15657 22799 15691
rect 22741 15651 22799 15657
rect 21358 15580 21364 15632
rect 21416 15620 21422 15632
rect 21606 15623 21664 15629
rect 21606 15620 21618 15623
rect 21416 15592 21618 15620
rect 21416 15580 21422 15592
rect 21606 15589 21618 15592
rect 21652 15589 21664 15623
rect 21606 15583 21664 15589
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 15712 15524 15945 15552
rect 15712 15512 15718 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 16390 15552 16396 15564
rect 15933 15515 15991 15521
rect 16040 15524 16396 15552
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 16040 15493 16068 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 17126 15552 17132 15564
rect 17087 15524 17132 15552
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 17402 15561 17408 15564
rect 17396 15552 17408 15561
rect 17363 15524 17408 15552
rect 17396 15515 17408 15524
rect 17402 15512 17408 15515
rect 17460 15512 17466 15564
rect 24026 15512 24032 15564
rect 24084 15552 24090 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 24084 15524 24593 15552
rect 24084 15512 24090 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 14884 15456 16037 15484
rect 14884 15444 14890 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16206 15484 16212 15496
rect 16167 15456 16212 15484
rect 16025 15447 16083 15453
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19484 15456 19625 15484
rect 19484 15444 19490 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 20898 15444 20904 15496
rect 20956 15484 20962 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 20956 15456 21373 15484
rect 20956 15444 20962 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 24762 15416 24768 15428
rect 24723 15388 24768 15416
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 15286 15308 15292 15360
rect 15344 15348 15350 15360
rect 15565 15351 15623 15357
rect 15565 15348 15577 15351
rect 15344 15320 15577 15348
rect 15344 15308 15350 15320
rect 15565 15317 15577 15320
rect 15611 15348 15623 15351
rect 16482 15348 16488 15360
rect 15611 15320 16488 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 18288 15320 18521 15348
rect 18288 15308 18294 15320
rect 18509 15317 18521 15320
rect 18555 15317 18567 15351
rect 18509 15311 18567 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 14737 15147 14795 15153
rect 14737 15113 14749 15147
rect 14783 15144 14795 15147
rect 14826 15144 14832 15156
rect 14783 15116 14832 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15144 16267 15147
rect 16390 15144 16396 15156
rect 16255 15116 16396 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 17184 15116 17233 15144
rect 17184 15104 17190 15116
rect 17221 15113 17233 15116
rect 17267 15144 17279 15147
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 17267 15116 18337 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 21726 15144 21732 15156
rect 21683 15116 21732 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 15008 15163 15011
rect 16206 15008 16212 15020
rect 15151 14980 16212 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 18340 15008 18368 15107
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 22244 15116 22293 15144
rect 22244 15104 22250 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22281 15107 22339 15113
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 24397 15147 24455 15153
rect 24397 15144 24409 15147
rect 24084 15116 24409 15144
rect 24084 15104 24090 15116
rect 24397 15113 24409 15116
rect 24443 15113 24455 15147
rect 24397 15107 24455 15113
rect 20898 15036 20904 15088
rect 20956 15076 20962 15088
rect 21913 15079 21971 15085
rect 21913 15076 21925 15079
rect 20956 15048 21925 15076
rect 20956 15036 20962 15048
rect 21913 15045 21925 15048
rect 21959 15076 21971 15079
rect 23382 15076 23388 15088
rect 21959 15048 23388 15076
rect 21959 15045 21971 15048
rect 21913 15039 21971 15045
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 18340 14980 18521 15008
rect 16761 14971 16819 14977
rect 18509 14977 18521 14980
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 12676 14912 13001 14940
rect 12676 14900 12682 14912
rect 12989 14909 13001 14912
rect 13035 14940 13047 14943
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13035 14912 13461 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16776 14940 16804 14971
rect 17402 14940 17408 14952
rect 16163 14912 17408 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 17402 14900 17408 14912
rect 17460 14940 17466 14952
rect 17589 14943 17647 14949
rect 17589 14940 17601 14943
rect 17460 14912 17601 14940
rect 17460 14900 17466 14912
rect 17589 14909 17601 14912
rect 17635 14909 17647 14943
rect 21450 14940 21456 14952
rect 21411 14912 21456 14940
rect 17589 14903 17647 14909
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 22465 14943 22523 14949
rect 22465 14909 22477 14943
rect 22511 14940 22523 14943
rect 24578 14940 24584 14952
rect 22511 14912 23152 14940
rect 24539 14912 24584 14940
rect 22511 14909 22523 14912
rect 22465 14903 22523 14909
rect 16577 14875 16635 14881
rect 16577 14872 16589 14875
rect 14844 14844 16589 14872
rect 14844 14816 14872 14844
rect 16577 14841 16589 14844
rect 16623 14841 16635 14875
rect 16577 14835 16635 14841
rect 18230 14832 18236 14884
rect 18288 14872 18294 14884
rect 18754 14875 18812 14881
rect 18754 14872 18766 14875
rect 18288 14844 18766 14872
rect 18288 14832 18294 14844
rect 18754 14841 18766 14844
rect 18800 14841 18812 14875
rect 18754 14835 18812 14841
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 14826 14804 14832 14816
rect 14415 14776 14832 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15194 14804 15200 14816
rect 15155 14776 15200 14804
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 19978 14804 19984 14816
rect 19935 14776 19984 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 21358 14804 21364 14816
rect 21319 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 23124 14813 23152 14912
rect 24578 14900 24584 14912
rect 24636 14940 24642 14952
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24636 14912 25145 14940
rect 24636 14900 24642 14912
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 23109 14807 23167 14813
rect 23109 14773 23121 14807
rect 23155 14804 23167 14807
rect 23750 14804 23756 14816
rect 23155 14776 23756 14804
rect 23155 14773 23167 14776
rect 23109 14767 23167 14773
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 24762 14804 24768 14816
rect 24723 14776 24768 14804
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15657 14603 15715 14609
rect 15657 14600 15669 14603
rect 15252 14572 15669 14600
rect 15252 14560 15258 14572
rect 15657 14569 15669 14572
rect 15703 14600 15715 14603
rect 16022 14600 16028 14612
rect 15703 14572 16028 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 18046 14600 18052 14612
rect 18007 14572 18052 14600
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 21450 14600 21456 14612
rect 21411 14572 21456 14600
rect 21450 14560 21456 14572
rect 21508 14600 21514 14612
rect 23201 14603 23259 14609
rect 23201 14600 23213 14603
rect 21508 14572 23213 14600
rect 21508 14560 21514 14572
rect 23201 14569 23213 14572
rect 23247 14569 23259 14603
rect 23201 14563 23259 14569
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 24949 14603 25007 14609
rect 24949 14600 24961 14603
rect 24912 14572 24961 14600
rect 24912 14560 24918 14572
rect 24949 14569 24961 14572
rect 24995 14569 25007 14603
rect 24949 14563 25007 14569
rect 15105 14535 15163 14541
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 15286 14532 15292 14544
rect 15151 14504 15292 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 16206 14492 16212 14544
rect 16264 14541 16270 14544
rect 16264 14535 16328 14541
rect 16264 14501 16282 14535
rect 16316 14501 16328 14535
rect 16264 14495 16328 14501
rect 16264 14492 16270 14495
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13228 14436 14105 14464
rect 13228 14424 13234 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 16025 14467 16083 14473
rect 16025 14464 16037 14467
rect 15528 14436 16037 14464
rect 15528 14424 15534 14436
rect 16025 14433 16037 14436
rect 16071 14464 16083 14467
rect 16758 14464 16764 14476
rect 16071 14436 16764 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16758 14424 16764 14436
rect 16816 14464 16822 14476
rect 17126 14464 17132 14476
rect 16816 14436 17132 14464
rect 16816 14424 16822 14436
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 20898 14464 20904 14476
rect 20859 14436 20904 14464
rect 20898 14424 20904 14436
rect 20956 14424 20962 14476
rect 21910 14424 21916 14476
rect 21968 14464 21974 14476
rect 22005 14467 22063 14473
rect 22005 14464 22017 14467
rect 21968 14436 22017 14464
rect 21968 14424 21974 14436
rect 22005 14433 22017 14436
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14433 23627 14467
rect 23569 14427 23627 14433
rect 23661 14467 23719 14473
rect 23661 14433 23673 14467
rect 23707 14464 23719 14467
rect 24026 14464 24032 14476
rect 23707 14436 24032 14464
rect 23707 14433 23719 14436
rect 23661 14427 23719 14433
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18969 14399 19027 14405
rect 18969 14396 18981 14399
rect 18104 14368 18981 14396
rect 18104 14356 18110 14368
rect 18969 14365 18981 14368
rect 19015 14396 19027 14399
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19015 14368 19533 14396
rect 19015 14365 19027 14368
rect 18969 14359 19027 14365
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 14274 14328 14280 14340
rect 14235 14300 14280 14328
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19628 14328 19656 14359
rect 19978 14328 19984 14340
rect 19392 14300 19984 14328
rect 19392 14288 19398 14300
rect 19978 14288 19984 14300
rect 20036 14328 20042 14340
rect 20073 14331 20131 14337
rect 20073 14328 20085 14331
rect 20036 14300 20085 14328
rect 20036 14288 20042 14300
rect 20073 14297 20085 14300
rect 20119 14297 20131 14331
rect 20073 14291 20131 14297
rect 13262 14260 13268 14272
rect 13223 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 18288 14232 18521 14260
rect 18288 14220 18294 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 18509 14223 18567 14229
rect 18966 14220 18972 14272
rect 19024 14260 19030 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 19024 14232 19073 14260
rect 19024 14220 19030 14232
rect 19061 14229 19073 14232
rect 19107 14229 19119 14263
rect 21082 14260 21088 14272
rect 21043 14232 21088 14260
rect 19061 14223 19119 14229
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 22186 14260 22192 14272
rect 22147 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23017 14263 23075 14269
rect 23017 14260 23029 14263
rect 22796 14232 23029 14260
rect 22796 14220 22802 14232
rect 23017 14229 23029 14232
rect 23063 14260 23075 14263
rect 23584 14260 23612 14427
rect 24026 14424 24032 14436
rect 24084 14424 24090 14476
rect 24394 14424 24400 14476
rect 24452 14464 24458 14476
rect 24765 14467 24823 14473
rect 24765 14464 24777 14467
rect 24452 14436 24777 14464
rect 24452 14424 24458 14436
rect 24765 14433 24777 14436
rect 24811 14464 24823 14467
rect 25590 14464 25596 14476
rect 24811 14436 25596 14464
rect 24811 14433 24823 14436
rect 24765 14427 24823 14433
rect 25590 14424 25596 14436
rect 25648 14424 25654 14476
rect 23842 14396 23848 14408
rect 23803 14368 23848 14396
rect 23842 14356 23848 14368
rect 23900 14356 23906 14408
rect 23063 14232 23612 14260
rect 23063 14229 23075 14232
rect 23017 14223 23075 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 13078 14056 13084 14068
rect 13039 14028 13084 14056
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13449 14059 13507 14065
rect 13449 14056 13461 14059
rect 13228 14028 13461 14056
rect 13228 14016 13234 14028
rect 13449 14025 13461 14028
rect 13495 14025 13507 14059
rect 14182 14056 14188 14068
rect 14143 14028 14188 14056
rect 13449 14019 13507 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14458 14056 14464 14068
rect 14419 14028 14464 14056
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 14884 14028 15669 14056
rect 14884 14016 14890 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 16264 14028 17049 14056
rect 16264 14016 16270 14028
rect 15197 13991 15255 13997
rect 15197 13957 15209 13991
rect 15243 13988 15255 13991
rect 16316 13988 16344 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 18046 14056 18052 14068
rect 18007 14028 18052 14056
rect 17037 14019 17095 14025
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19426 14056 19432 14068
rect 19199 14028 19432 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19521 14059 19579 14065
rect 19521 14025 19533 14059
rect 19567 14056 19579 14059
rect 19610 14056 19616 14068
rect 19567 14028 19616 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 19610 14016 19616 14028
rect 19668 14056 19674 14068
rect 20806 14056 20812 14068
rect 19668 14028 20812 14056
rect 19668 14016 19674 14028
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 23109 14059 23167 14065
rect 23109 14056 23121 14059
rect 21416 14028 23121 14056
rect 21416 14016 21422 14028
rect 23109 14025 23121 14028
rect 23155 14056 23167 14059
rect 23842 14056 23848 14068
rect 23155 14028 23848 14056
rect 23155 14025 23167 14028
rect 23109 14019 23167 14025
rect 23842 14016 23848 14028
rect 23900 14056 23906 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 23900 14028 25053 14056
rect 23900 14016 23906 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25590 14056 25596 14068
rect 25551 14028 25596 14056
rect 25041 14019 25099 14025
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 16758 13988 16764 14000
rect 15243 13960 16344 13988
rect 16719 13960 16764 13988
rect 15243 13957 15255 13960
rect 15197 13951 15255 13957
rect 16316 13929 16344 13960
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 20898 13948 20904 14000
rect 20956 13988 20962 14000
rect 21545 13991 21603 13997
rect 21545 13988 21557 13991
rect 20956 13960 21557 13988
rect 20956 13948 20962 13960
rect 21545 13957 21557 13960
rect 21591 13957 21603 13991
rect 21545 13951 21603 13957
rect 21910 13948 21916 14000
rect 21968 13988 21974 14000
rect 22005 13991 22063 13997
rect 22005 13988 22017 13991
rect 21968 13960 22017 13988
rect 21968 13948 21974 13960
rect 22005 13957 22017 13960
rect 22051 13957 22063 13991
rect 23382 13988 23388 14000
rect 23343 13960 23388 13988
rect 22005 13951 22063 13957
rect 23382 13948 23388 13960
rect 23440 13988 23446 14000
rect 23440 13960 23704 13988
rect 23440 13948 23446 13960
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15488 13892 16129 13920
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 14182 13852 14188 13864
rect 13679 13824 14188 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14516 13824 14657 13852
rect 14516 13812 14522 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14826 13812 14832 13864
rect 14884 13812 14890 13864
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15488 13861 15516 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18288 13892 18613 13920
rect 18288 13880 18294 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 23676 13929 23704 13960
rect 23661 13923 23719 13929
rect 19392 13892 19748 13920
rect 19392 13880 19398 13892
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15436 13824 15485 13852
rect 15436 13812 15442 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 16022 13852 16028 13864
rect 15983 13824 16028 13852
rect 15473 13815 15531 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 17770 13852 17776 13864
rect 17731 13824 17776 13852
rect 17770 13812 17776 13824
rect 17828 13852 17834 13864
rect 17828 13824 17908 13852
rect 17828 13812 17834 13824
rect 13814 13716 13820 13728
rect 13775 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14844 13725 14872 13812
rect 17880 13784 17908 13824
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 18196 13824 18521 13852
rect 18196 13812 18202 13824
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 19610 13852 19616 13864
rect 19571 13824 19616 13852
rect 18509 13815 18567 13821
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 19720 13852 19748 13892
rect 23661 13889 23673 13923
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 19869 13855 19927 13861
rect 19869 13852 19881 13855
rect 19720 13824 19881 13852
rect 19869 13821 19881 13824
rect 19915 13821 19927 13855
rect 19869 13815 19927 13821
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13852 22523 13855
rect 22511 13824 24072 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 24044 13796 24072 13824
rect 18417 13787 18475 13793
rect 18417 13784 18429 13787
rect 17880 13756 18429 13784
rect 18417 13753 18429 13756
rect 18463 13753 18475 13787
rect 18417 13747 18475 13753
rect 23566 13744 23572 13796
rect 23624 13784 23630 13796
rect 23906 13787 23964 13793
rect 23906 13784 23918 13787
rect 23624 13756 23918 13784
rect 23624 13744 23630 13756
rect 23906 13753 23918 13756
rect 23952 13753 23964 13787
rect 23906 13747 23964 13753
rect 24026 13744 24032 13796
rect 24084 13744 24090 13796
rect 14829 13719 14887 13725
rect 14829 13685 14841 13719
rect 14875 13685 14887 13719
rect 14829 13679 14887 13685
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 17586 13716 17592 13728
rect 16908 13688 17592 13716
rect 16908 13676 16914 13688
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 20990 13716 20996 13728
rect 20903 13688 20996 13716
rect 20990 13676 20996 13688
rect 21048 13716 21054 13728
rect 21634 13716 21640 13728
rect 21048 13688 21640 13716
rect 21048 13676 21054 13688
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 22557 13719 22615 13725
rect 22557 13685 22569 13719
rect 22603 13716 22615 13719
rect 23106 13716 23112 13728
rect 22603 13688 23112 13716
rect 22603 13685 22615 13688
rect 22557 13679 22615 13685
rect 23106 13676 23112 13688
rect 23164 13676 23170 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 14369 13515 14427 13521
rect 14369 13481 14381 13515
rect 14415 13512 14427 13515
rect 14734 13512 14740 13524
rect 14415 13484 14740 13512
rect 14415 13481 14427 13484
rect 14369 13475 14427 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 17126 13512 17132 13524
rect 15611 13484 17132 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 17126 13472 17132 13484
rect 17184 13512 17190 13524
rect 17589 13515 17647 13521
rect 17589 13512 17601 13515
rect 17184 13484 17601 13512
rect 17184 13472 17190 13484
rect 17589 13481 17601 13484
rect 17635 13481 17647 13515
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 17589 13475 17647 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19153 13515 19211 13521
rect 19153 13481 19165 13515
rect 19199 13512 19211 13515
rect 19334 13512 19340 13524
rect 19199 13484 19340 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 23198 13512 23204 13524
rect 23159 13484 23204 13512
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23842 13472 23848 13524
rect 23900 13512 23906 13524
rect 24210 13512 24216 13524
rect 23900 13484 24216 13512
rect 23900 13472 23906 13484
rect 24210 13472 24216 13484
rect 24268 13472 24274 13524
rect 24762 13512 24768 13524
rect 24723 13484 24768 13512
rect 24762 13472 24768 13484
rect 24820 13472 24826 13524
rect 16025 13447 16083 13453
rect 16025 13413 16037 13447
rect 16071 13444 16083 13447
rect 16206 13444 16212 13456
rect 16071 13416 16212 13444
rect 16071 13413 16083 13416
rect 16025 13407 16083 13413
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19610 13444 19616 13456
rect 19484 13416 19616 13444
rect 19484 13404 19490 13416
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 23106 13444 23112 13456
rect 23067 13416 23112 13444
rect 23106 13404 23112 13416
rect 23164 13404 23170 13456
rect 14182 13376 14188 13388
rect 14143 13348 14188 13376
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 16298 13376 16304 13388
rect 15979 13348 16304 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 17494 13376 17500 13388
rect 17455 13348 17500 13376
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 18782 13336 18788 13388
rect 18840 13376 18846 13388
rect 19518 13376 19524 13388
rect 18840 13348 19524 13376
rect 18840 13336 18846 13348
rect 19518 13336 19524 13348
rect 19576 13376 19582 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19576 13348 19717 13376
rect 19576 13336 19582 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 21082 13336 21088 13388
rect 21140 13376 21146 13388
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 21140 13348 21281 13376
rect 21140 13336 21146 13348
rect 21269 13345 21281 13348
rect 21315 13345 21327 13379
rect 24578 13376 24584 13388
rect 24539 13348 24584 13376
rect 21269 13339 21327 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 16206 13308 16212 13320
rect 16167 13280 16212 13308
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 17678 13308 17684 13320
rect 17639 13280 17684 13308
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 18472 13280 19901 13308
rect 18472 13268 18478 13280
rect 19889 13277 19901 13280
rect 19935 13308 19947 13311
rect 20990 13308 20996 13320
rect 19935 13280 20996 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 21634 13308 21640 13320
rect 21591 13280 21640 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 23385 13311 23443 13317
rect 23385 13277 23397 13311
rect 23431 13308 23443 13311
rect 23431 13280 23612 13308
rect 23431 13277 23443 13280
rect 23385 13271 23443 13277
rect 16669 13243 16727 13249
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 16758 13240 16764 13252
rect 16715 13212 16764 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 16758 13200 16764 13212
rect 16816 13240 16822 13252
rect 17129 13243 17187 13249
rect 17129 13240 17141 13243
rect 16816 13212 17141 13240
rect 16816 13200 16822 13212
rect 17129 13209 17141 13212
rect 17175 13209 17187 13243
rect 17129 13203 17187 13209
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13240 18843 13243
rect 19242 13240 19248 13252
rect 18831 13212 19248 13240
rect 18831 13209 18843 13212
rect 18785 13203 18843 13209
rect 19242 13200 19248 13212
rect 19300 13200 19306 13252
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 20901 13243 20959 13249
rect 20901 13240 20913 13243
rect 19392 13212 20913 13240
rect 19392 13200 19398 13212
rect 20901 13209 20913 13212
rect 20947 13209 20959 13243
rect 22738 13240 22744 13252
rect 22699 13212 22744 13240
rect 20901 13203 20959 13209
rect 22738 13200 22744 13212
rect 22796 13200 22802 13252
rect 23584 13184 23612 13280
rect 16942 13172 16948 13184
rect 16903 13144 16948 13172
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 20622 13172 20628 13184
rect 20583 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 21910 13172 21916 13184
rect 21871 13144 21916 13172
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22281 13175 22339 13181
rect 22281 13172 22293 13175
rect 22152 13144 22293 13172
rect 22152 13132 22158 13144
rect 22281 13141 22293 13144
rect 22327 13141 22339 13175
rect 22281 13135 22339 13141
rect 23566 13132 23572 13184
rect 23624 13172 23630 13184
rect 23753 13175 23811 13181
rect 23753 13172 23765 13175
rect 23624 13144 23765 13172
rect 23624 13132 23630 13144
rect 23753 13141 23765 13144
rect 23799 13141 23811 13175
rect 23753 13135 23811 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 14001 12971 14059 12977
rect 14001 12937 14013 12971
rect 14047 12968 14059 12971
rect 15470 12968 15476 12980
rect 14047 12940 15476 12968
rect 14047 12937 14059 12940
rect 14001 12931 14059 12937
rect 14108 12841 14136 12940
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16761 12971 16819 12977
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 16850 12968 16856 12980
rect 16807 12940 16856 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17589 12971 17647 12977
rect 17589 12937 17601 12971
rect 17635 12968 17647 12971
rect 17678 12968 17684 12980
rect 17635 12940 17684 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 20441 12971 20499 12977
rect 20441 12937 20453 12971
rect 20487 12968 20499 12971
rect 20806 12968 20812 12980
rect 20487 12940 20812 12968
rect 20487 12937 20499 12940
rect 20441 12931 20499 12937
rect 20806 12928 20812 12940
rect 20864 12968 20870 12980
rect 21358 12968 21364 12980
rect 20864 12940 21364 12968
rect 20864 12928 20870 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 21634 12928 21640 12980
rect 21692 12968 21698 12980
rect 21913 12971 21971 12977
rect 21913 12968 21925 12971
rect 21692 12940 21925 12968
rect 21692 12928 21698 12940
rect 21913 12937 21925 12940
rect 21959 12937 21971 12971
rect 22278 12968 22284 12980
rect 22239 12940 22284 12968
rect 21913 12931 21971 12937
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 23106 12968 23112 12980
rect 23067 12940 23112 12968
rect 23106 12928 23112 12940
rect 23164 12928 23170 12980
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24670 12968 24676 12980
rect 24535 12940 24676 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 16117 12903 16175 12909
rect 16117 12869 16129 12903
rect 16163 12900 16175 12903
rect 16298 12900 16304 12912
rect 16163 12872 16304 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 19610 12860 19616 12912
rect 19668 12900 19674 12912
rect 20073 12903 20131 12909
rect 20073 12900 20085 12903
rect 19668 12872 20085 12900
rect 19668 12860 19674 12872
rect 20073 12869 20085 12872
rect 20119 12900 20131 12903
rect 22554 12900 22560 12912
rect 20119 12872 22560 12900
rect 20119 12869 20131 12872
rect 20073 12863 20131 12869
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 22833 12903 22891 12909
rect 22833 12869 22845 12903
rect 22879 12900 22891 12903
rect 23198 12900 23204 12912
rect 22879 12872 23204 12900
rect 22879 12869 22891 12872
rect 22833 12863 22891 12869
rect 23198 12860 23204 12872
rect 23256 12860 23262 12912
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 19518 12832 19524 12844
rect 19479 12804 19524 12832
rect 14093 12795 14151 12801
rect 19518 12792 19524 12804
rect 19576 12792 19582 12844
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12832 21235 12835
rect 21358 12832 21364 12844
rect 21223 12804 21364 12832
rect 21223 12801 21235 12804
rect 21177 12795 21235 12801
rect 21358 12792 21364 12804
rect 21416 12832 21422 12844
rect 21910 12832 21916 12844
rect 21416 12804 21916 12832
rect 21416 12792 21422 12804
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 16577 12767 16635 12773
rect 16577 12764 16589 12767
rect 16540 12736 16589 12764
rect 16540 12724 16546 12736
rect 16577 12733 16589 12736
rect 16623 12764 16635 12767
rect 16942 12764 16948 12776
rect 16623 12736 16948 12764
rect 16623 12733 16635 12736
rect 16577 12727 16635 12733
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 18782 12764 18788 12776
rect 18743 12736 18788 12764
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19392 12736 19437 12764
rect 19392 12724 19398 12736
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 20680 12736 20913 12764
rect 20680 12724 20686 12736
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 24578 12764 24584 12776
rect 22152 12736 22197 12764
rect 24539 12736 24584 12764
rect 22152 12724 22158 12736
rect 24578 12724 24584 12736
rect 24636 12764 24642 12776
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24636 12736 25145 12764
rect 24636 12724 24642 12736
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 14366 12705 14372 12708
rect 13633 12699 13691 12705
rect 13633 12696 13645 12699
rect 12676 12668 13645 12696
rect 12676 12656 12682 12668
rect 13633 12665 13645 12668
rect 13679 12696 13691 12699
rect 14338 12699 14372 12705
rect 14338 12696 14350 12699
rect 13679 12668 14350 12696
rect 13679 12665 13691 12668
rect 13633 12659 13691 12665
rect 14338 12665 14350 12668
rect 14338 12659 14372 12665
rect 14366 12656 14372 12659
rect 14424 12656 14430 12708
rect 19242 12656 19248 12708
rect 19300 12696 19306 12708
rect 19429 12699 19487 12705
rect 19429 12696 19441 12699
rect 19300 12668 19441 12696
rect 19300 12656 19306 12668
rect 19429 12665 19441 12668
rect 19475 12665 19487 12699
rect 19429 12659 19487 12665
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 20993 12699 21051 12705
rect 20993 12696 21005 12699
rect 20496 12668 21005 12696
rect 20496 12656 20502 12668
rect 20993 12665 21005 12668
rect 21039 12696 21051 12699
rect 23014 12696 23020 12708
rect 21039 12668 23020 12696
rect 21039 12665 21051 12668
rect 20993 12659 21051 12665
rect 23014 12656 23020 12668
rect 23072 12656 23078 12708
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 12492 12600 13093 12628
rect 12492 12588 12498 12600
rect 13081 12597 13093 12600
rect 13127 12597 13139 12631
rect 15470 12628 15476 12640
rect 15431 12600 15476 12628
rect 13081 12591 13139 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 17221 12631 17279 12637
rect 17221 12597 17233 12631
rect 17267 12628 17279 12631
rect 17494 12628 17500 12640
rect 17267 12600 17500 12628
rect 17267 12597 17279 12600
rect 17221 12591 17279 12597
rect 17494 12588 17500 12600
rect 17552 12628 17558 12640
rect 18046 12628 18052 12640
rect 17552 12600 18052 12628
rect 17552 12588 17558 12600
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18414 12628 18420 12640
rect 18375 12600 18420 12628
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18969 12631 19027 12637
rect 18969 12597 18981 12631
rect 19015 12628 19027 12631
rect 19150 12628 19156 12640
rect 19015 12600 19156 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 20530 12628 20536 12640
rect 20491 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 21545 12631 21603 12637
rect 21545 12628 21557 12631
rect 21140 12600 21557 12628
rect 21140 12588 21146 12600
rect 21545 12597 21557 12600
rect 21591 12597 21603 12631
rect 24762 12628 24768 12640
rect 24723 12600 24768 12628
rect 21545 12591 21603 12597
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12492 12396 12537 12424
rect 12492 12384 12498 12396
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 13538 12424 13544 12436
rect 13136 12396 13544 12424
rect 13136 12384 13142 12396
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 16206 12424 16212 12436
rect 15151 12396 16212 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 16206 12384 16212 12396
rect 16264 12424 16270 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 16264 12396 16957 12424
rect 16264 12384 16270 12396
rect 16945 12393 16957 12396
rect 16991 12424 17003 12427
rect 17494 12424 17500 12436
rect 16991 12396 17172 12424
rect 17455 12396 17500 12424
rect 16991 12393 17003 12396
rect 16945 12387 17003 12393
rect 17144 12368 17172 12396
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 19116 12396 19257 12424
rect 19116 12384 19122 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 19245 12387 19303 12393
rect 19536 12396 19625 12424
rect 19536 12368 19564 12396
rect 19613 12393 19625 12396
rect 19659 12424 19671 12427
rect 20530 12424 20536 12436
rect 19659 12396 20536 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 23750 12424 23756 12436
rect 23711 12396 23756 12424
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 12529 12359 12587 12365
rect 12529 12356 12541 12359
rect 11664 12328 12541 12356
rect 11664 12316 11670 12328
rect 12529 12325 12541 12328
rect 12575 12356 12587 12359
rect 13722 12356 13728 12368
rect 12575 12328 13728 12356
rect 12575 12325 12587 12328
rect 12529 12319 12587 12325
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 14550 12356 14556 12368
rect 14332 12328 14556 12356
rect 14332 12316 14338 12328
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 17126 12316 17132 12368
rect 17184 12316 17190 12368
rect 19518 12316 19524 12368
rect 19576 12316 19582 12368
rect 21358 12365 21364 12368
rect 21352 12356 21364 12365
rect 21319 12328 21364 12356
rect 21352 12319 21364 12328
rect 21358 12316 21364 12319
rect 21416 12316 21422 12368
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13228 12260 14013 12288
rect 13228 12248 13234 12260
rect 14001 12257 14013 12260
rect 14047 12257 14059 12291
rect 15470 12288 15476 12300
rect 14001 12251 14059 12257
rect 14292 12260 15476 12288
rect 14292 12232 14320 12260
rect 15470 12248 15476 12260
rect 15528 12288 15534 12300
rect 15832 12291 15890 12297
rect 15832 12288 15844 12291
rect 15528 12260 15844 12288
rect 15528 12248 15534 12260
rect 15832 12257 15844 12260
rect 15878 12288 15890 12291
rect 16298 12288 16304 12300
rect 15878 12260 16304 12288
rect 15878 12257 15890 12260
rect 15832 12251 15890 12257
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 19242 12288 19248 12300
rect 18739 12260 19248 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12288 19763 12291
rect 19978 12288 19984 12300
rect 19751 12260 19984 12288
rect 19751 12257 19763 12260
rect 19705 12251 19763 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 20898 12248 20904 12300
rect 20956 12288 20962 12300
rect 21085 12291 21143 12297
rect 21085 12288 21097 12291
rect 20956 12260 21097 12288
rect 20956 12248 20962 12260
rect 21085 12257 21097 12260
rect 21131 12257 21143 12291
rect 21085 12251 21143 12257
rect 22738 12248 22744 12300
rect 22796 12288 22802 12300
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 22796 12260 23581 12288
rect 22796 12248 22802 12260
rect 23569 12257 23581 12260
rect 23615 12257 23627 12291
rect 24578 12288 24584 12300
rect 24539 12260 24584 12288
rect 23569 12251 23627 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13630 12220 13636 12232
rect 13587 12192 13636 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13630 12180 13636 12192
rect 13688 12220 13694 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13688 12192 14105 12220
rect 13688 12180 13694 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14274 12220 14280 12232
rect 14187 12192 14280 12220
rect 14093 12183 14151 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 15562 12220 15568 12232
rect 15523 12192 15568 12220
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 20070 12220 20076 12232
rect 19935 12192 20076 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 14734 12152 14740 12164
rect 11756 12124 14740 12152
rect 11756 12112 11762 12124
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 17865 12155 17923 12161
rect 17865 12152 17877 12155
rect 16908 12124 17877 12152
rect 16908 12112 16914 12124
rect 17865 12121 17877 12124
rect 17911 12121 17923 12155
rect 17865 12115 17923 12121
rect 23109 12155 23167 12161
rect 23109 12121 23121 12155
rect 23155 12152 23167 12155
rect 23566 12152 23572 12164
rect 23155 12124 23572 12152
rect 23155 12121 23167 12124
rect 23109 12115 23167 12121
rect 23566 12112 23572 12124
rect 23624 12112 23630 12164
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 13170 12084 13176 12096
rect 12115 12056 13176 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 14182 12084 14188 12096
rect 13679 12056 14188 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 14182 12044 14188 12056
rect 14240 12084 14246 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14240 12056 14657 12084
rect 14240 12044 14246 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 19061 12087 19119 12093
rect 19061 12053 19073 12087
rect 19107 12084 19119 12087
rect 19242 12084 19248 12096
rect 19107 12056 19248 12084
rect 19107 12053 19119 12056
rect 19061 12047 19119 12053
rect 19242 12044 19248 12056
rect 19300 12084 19306 12096
rect 19426 12084 19432 12096
rect 19300 12056 19432 12084
rect 19300 12044 19306 12056
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 20533 12087 20591 12093
rect 20533 12084 20545 12087
rect 20496 12056 20545 12084
rect 20496 12044 20502 12056
rect 20533 12053 20545 12056
rect 20579 12053 20591 12087
rect 22462 12084 22468 12096
rect 22423 12056 22468 12084
rect 20533 12047 20591 12053
rect 22462 12044 22468 12056
rect 22520 12044 22526 12096
rect 24121 12087 24179 12093
rect 24121 12053 24133 12087
rect 24167 12084 24179 12087
rect 24210 12084 24216 12096
rect 24167 12056 24216 12084
rect 24167 12053 24179 12056
rect 24121 12047 24179 12053
rect 24210 12044 24216 12056
rect 24268 12044 24274 12096
rect 24762 12084 24768 12096
rect 24723 12056 24768 12084
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 11425 11883 11483 11889
rect 11425 11849 11437 11883
rect 11471 11880 11483 11883
rect 11606 11880 11612 11892
rect 11471 11852 11612 11880
rect 11471 11849 11483 11852
rect 11425 11843 11483 11849
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12434 11880 12440 11892
rect 12207 11852 12440 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 14274 11880 14280 11892
rect 13127 11852 14280 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 15562 11880 15568 11892
rect 15523 11852 15568 11880
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 16393 11883 16451 11889
rect 16393 11849 16405 11883
rect 16439 11880 16451 11883
rect 16482 11880 16488 11892
rect 16439 11852 16488 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 16632 11852 17785 11880
rect 16632 11840 16638 11852
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 20070 11880 20076 11892
rect 20031 11852 20076 11880
rect 17773 11843 17831 11849
rect 11793 11815 11851 11821
rect 11793 11781 11805 11815
rect 11839 11812 11851 11815
rect 12618 11812 12624 11824
rect 11839 11784 12624 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 15580 11744 15608 11840
rect 16301 11815 16359 11821
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 16347 11784 16988 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 16960 11756 16988 11784
rect 16574 11744 16580 11756
rect 15580 11716 16580 11744
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16850 11744 16856 11756
rect 16811 11716 16856 11744
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17788 11744 17816 11843
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20898 11880 20904 11892
rect 20487 11852 20904 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17000 11716 17093 11744
rect 17788 11716 18061 11744
rect 17000 11704 17006 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 13538 11676 13544 11688
rect 13495 11648 13544 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 16758 11676 16764 11688
rect 16719 11648 16764 11676
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 18064 11676 18092 11707
rect 20456 11676 20484 11843
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21910 11880 21916 11892
rect 21871 11852 21916 11880
rect 21910 11840 21916 11852
rect 21968 11840 21974 11892
rect 22738 11880 22744 11892
rect 22699 11852 22744 11880
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 23934 11744 23940 11756
rect 23523 11716 23940 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23934 11704 23940 11716
rect 23992 11744 23998 11756
rect 24121 11747 24179 11753
rect 24121 11744 24133 11747
rect 23992 11716 24133 11744
rect 23992 11704 23998 11716
rect 24121 11713 24133 11716
rect 24167 11713 24179 11747
rect 24121 11707 24179 11713
rect 24210 11704 24216 11756
rect 24268 11744 24274 11756
rect 24268 11716 24313 11744
rect 24268 11704 24274 11716
rect 20530 11676 20536 11688
rect 18064 11648 20536 11676
rect 20530 11636 20536 11648
rect 20588 11636 20594 11688
rect 12713 11611 12771 11617
rect 12713 11577 12725 11611
rect 12759 11608 12771 11611
rect 13786 11611 13844 11617
rect 13786 11608 13798 11611
rect 12759 11580 13798 11608
rect 12759 11577 12771 11580
rect 12713 11571 12771 11577
rect 13786 11577 13798 11580
rect 13832 11608 13844 11611
rect 14642 11608 14648 11620
rect 13832 11580 14648 11608
rect 13832 11577 13844 11580
rect 13786 11571 13844 11577
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 17586 11608 17592 11620
rect 17420 11580 17592 11608
rect 14918 11540 14924 11552
rect 14879 11512 14924 11540
rect 14918 11500 14924 11512
rect 14976 11500 14982 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 17420 11549 17448 11580
rect 17586 11568 17592 11580
rect 17644 11608 17650 11620
rect 18230 11608 18236 11620
rect 17644 11580 18236 11608
rect 17644 11568 17650 11580
rect 18230 11568 18236 11580
rect 18288 11617 18294 11620
rect 18288 11611 18352 11617
rect 18288 11577 18306 11611
rect 18340 11577 18352 11611
rect 18288 11571 18352 11577
rect 18288 11568 18294 11571
rect 20254 11568 20260 11620
rect 20312 11608 20318 11620
rect 20778 11611 20836 11617
rect 20778 11608 20790 11611
rect 20312 11580 20790 11608
rect 20312 11568 20318 11580
rect 20778 11577 20790 11580
rect 20824 11577 20836 11611
rect 24029 11611 24087 11617
rect 24029 11608 24041 11611
rect 20778 11571 20836 11577
rect 23032 11580 24041 11608
rect 23032 11552 23060 11580
rect 24029 11577 24041 11580
rect 24075 11577 24087 11611
rect 24029 11571 24087 11577
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 16816 11512 17417 11540
rect 16816 11500 16822 11512
rect 17405 11509 17417 11512
rect 17451 11509 17463 11543
rect 19426 11540 19432 11552
rect 19387 11512 19432 11540
rect 17405 11503 17463 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 23014 11540 23020 11552
rect 22975 11512 23020 11540
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 23658 11540 23664 11552
rect 23619 11512 23664 11540
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12250 11336 12256 11348
rect 12207 11308 12256 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 13170 11336 13176 11348
rect 13131 11308 13176 11336
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14642 11336 14648 11348
rect 14603 11308 14648 11336
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 16850 11336 16856 11348
rect 15335 11308 16856 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 17000 11308 18889 11336
rect 17000 11296 17006 11308
rect 18877 11305 18889 11308
rect 18923 11336 18935 11339
rect 19150 11336 19156 11348
rect 18923 11308 19156 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19150 11296 19156 11308
rect 19208 11336 19214 11348
rect 19426 11336 19432 11348
rect 19208 11308 19432 11336
rect 19208 11296 19214 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19576 11308 19625 11336
rect 19576 11296 19582 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 19797 11339 19855 11345
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 20622 11336 20628 11348
rect 19843 11308 20628 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 21085 11339 21143 11345
rect 21085 11336 21097 11339
rect 20956 11308 21097 11336
rect 20956 11296 20962 11308
rect 21085 11305 21097 11308
rect 21131 11305 21143 11339
rect 21085 11299 21143 11305
rect 21453 11339 21511 11345
rect 21453 11305 21465 11339
rect 21499 11336 21511 11339
rect 22002 11336 22008 11348
rect 21499 11308 22008 11336
rect 21499 11305 21511 11308
rect 21453 11299 21511 11305
rect 15657 11271 15715 11277
rect 15657 11237 15669 11271
rect 15703 11268 15715 11271
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 15703 11240 16129 11268
rect 15703 11237 15715 11240
rect 15657 11231 15715 11237
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 21100 11268 21128 11299
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 21100 11240 22324 11268
rect 16117 11231 16175 11237
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11296 11172 11989 11200
rect 11296 11160 11302 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 13998 11200 14004 11212
rect 13959 11172 14004 11200
rect 11977 11163 12035 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14093 11203 14151 11209
rect 14093 11169 14105 11203
rect 14139 11200 14151 11203
rect 15102 11200 15108 11212
rect 14139 11172 15108 11200
rect 14139 11169 14151 11172
rect 14093 11163 14151 11169
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 14108 11132 14136 11163
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 16482 11200 16488 11212
rect 15795 11172 16488 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 17126 11209 17132 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 16632 11172 16865 11200
rect 16632 11160 16638 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 17120 11200 17132 11209
rect 17087 11172 17132 11200
rect 16853 11163 16911 11169
rect 17120 11163 17132 11172
rect 17126 11160 17132 11163
rect 17184 11160 17190 11212
rect 22296 11209 22324 11240
rect 22462 11228 22468 11280
rect 22520 11277 22526 11280
rect 22520 11271 22584 11277
rect 22520 11237 22538 11271
rect 22572 11237 22584 11271
rect 22520 11231 22584 11237
rect 25225 11271 25283 11277
rect 25225 11237 25237 11271
rect 25271 11268 25283 11271
rect 25314 11268 25320 11280
rect 25271 11240 25320 11268
rect 25271 11237 25283 11240
rect 25225 11231 25283 11237
rect 22520 11228 22526 11231
rect 25314 11228 25320 11240
rect 25372 11228 25378 11280
rect 21261 11203 21319 11209
rect 21261 11200 21273 11203
rect 21192 11172 21273 11200
rect 13587 11104 14136 11132
rect 14185 11135 14243 11141
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 14185 11101 14197 11135
rect 14231 11132 14243 11135
rect 14366 11132 14372 11144
rect 14231 11104 14372 11132
rect 14231 11101 14243 11104
rect 14185 11095 14243 11101
rect 13722 11024 13728 11076
rect 13780 11064 13786 11076
rect 14200 11064 14228 11095
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 14918 11132 14924 11144
rect 14424 11104 14924 11132
rect 14424 11092 14430 11104
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15059 11104 15853 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15841 11101 15853 11104
rect 15887 11132 15899 11135
rect 16758 11132 16764 11144
rect 15887 11104 16764 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16298 11064 16304 11076
rect 13780 11036 14228 11064
rect 16259 11036 16304 11064
rect 13780 11024 13786 11036
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 18230 11064 18236 11076
rect 18191 11036 18236 11064
rect 18230 11024 18236 11036
rect 18288 11024 18294 11076
rect 19337 11067 19395 11073
rect 19337 11033 19349 11067
rect 19383 11064 19395 11067
rect 19978 11064 19984 11076
rect 19383 11036 19984 11064
rect 19383 11033 19395 11036
rect 19337 11027 19395 11033
rect 19978 11024 19984 11036
rect 20036 11064 20042 11076
rect 20036 11036 20668 11064
rect 20036 11024 20042 11036
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 1581 10999 1639 11005
rect 1581 10996 1593 10999
rect 1544 10968 1593 10996
rect 1544 10956 1550 10968
rect 1581 10965 1593 10968
rect 1627 10965 1639 10999
rect 11330 10996 11336 11008
rect 11291 10968 11336 10996
rect 1581 10959 1639 10965
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12529 10999 12587 11005
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 12894 10996 12900 11008
rect 12575 10968 12900 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 16117 10999 16175 11005
rect 16117 10965 16129 10999
rect 16163 10996 16175 10999
rect 16758 10996 16764 11008
rect 16163 10968 16764 10996
rect 16163 10965 16175 10968
rect 16117 10959 16175 10965
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 20254 10956 20260 11008
rect 20312 10996 20318 11008
rect 20533 10999 20591 11005
rect 20533 10996 20545 10999
rect 20312 10968 20545 10996
rect 20312 10956 20318 10968
rect 20533 10965 20545 10968
rect 20579 10965 20591 10999
rect 20640 10996 20668 11036
rect 20714 10996 20720 11008
rect 20640 10968 20720 10996
rect 20533 10959 20591 10965
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 21192 10996 21220 11172
rect 21261 11169 21273 11172
rect 21307 11169 21319 11203
rect 21261 11163 21319 11169
rect 22281 11203 22339 11209
rect 22281 11169 22293 11203
rect 22327 11200 22339 11203
rect 22370 11200 22376 11212
rect 22327 11172 22376 11200
rect 22327 11169 22339 11172
rect 22281 11163 22339 11169
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 25133 11203 25191 11209
rect 25133 11169 25145 11203
rect 25179 11200 25191 11203
rect 25590 11200 25596 11212
rect 25179 11172 25596 11200
rect 25179 11169 25191 11172
rect 25133 11163 25191 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 21821 11135 21879 11141
rect 21821 11101 21833 11135
rect 21867 11132 21879 11135
rect 21910 11132 21916 11144
rect 21867 11104 21916 11132
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 25406 11132 25412 11144
rect 25367 11104 25412 11132
rect 25406 11092 25412 11104
rect 25464 11092 25470 11144
rect 24762 11064 24768 11076
rect 24723 11036 24768 11064
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 22094 10996 22100 11008
rect 21192 10968 22100 10996
rect 22094 10956 22100 10968
rect 22152 10956 22158 11008
rect 23661 10999 23719 11005
rect 23661 10965 23673 10999
rect 23707 10996 23719 10999
rect 23934 10996 23940 11008
rect 23707 10968 23940 10996
rect 23707 10965 23719 10968
rect 23661 10959 23719 10965
rect 23934 10956 23940 10968
rect 23992 10996 23998 11008
rect 24305 10999 24363 11005
rect 24305 10996 24317 10999
rect 23992 10968 24317 10996
rect 23992 10956 23998 10968
rect 24305 10965 24317 10968
rect 24351 10996 24363 10999
rect 25406 10996 25412 11008
rect 24351 10968 25412 10996
rect 24351 10965 24363 10968
rect 24305 10959 24363 10965
rect 25406 10956 25412 10968
rect 25464 10956 25470 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 11238 10792 11244 10804
rect 11199 10764 11244 10792
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11514 10792 11520 10804
rect 11475 10764 11520 10792
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13872 10764 14013 10792
rect 13872 10752 13878 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15344 10764 15577 10792
rect 15344 10752 15350 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 16632 10764 16865 10792
rect 16632 10752 16638 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 16853 10755 16911 10761
rect 11256 10724 11284 10752
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 11256 10696 12449 10724
rect 12437 10693 12449 10696
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 13504 10696 15025 10724
rect 13504 10684 13510 10696
rect 15013 10693 15025 10696
rect 15059 10724 15071 10727
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 15059 10696 15209 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 16868 10724 16896 10755
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17589 10795 17647 10801
rect 17589 10792 17601 10795
rect 17184 10764 17601 10792
rect 17184 10752 17190 10764
rect 17589 10761 17601 10764
rect 17635 10792 17647 10795
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 17635 10764 18245 10792
rect 17635 10761 17647 10764
rect 17589 10755 17647 10761
rect 18233 10761 18245 10764
rect 18279 10792 18291 10795
rect 18874 10792 18880 10804
rect 18279 10764 18880 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21361 10795 21419 10801
rect 21361 10792 21373 10795
rect 20772 10764 21373 10792
rect 20772 10752 20778 10764
rect 21361 10761 21373 10764
rect 21407 10761 21419 10795
rect 22370 10792 22376 10804
rect 22331 10764 22376 10792
rect 21361 10755 21419 10761
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22520 10764 22753 10792
rect 22520 10752 22526 10764
rect 22741 10761 22753 10764
rect 22787 10761 22799 10795
rect 22741 10755 22799 10761
rect 25406 10752 25412 10804
rect 25464 10792 25470 10804
rect 25961 10795 26019 10801
rect 25961 10792 25973 10795
rect 25464 10764 25973 10792
rect 25464 10752 25470 10764
rect 25961 10761 25973 10764
rect 26007 10761 26019 10795
rect 25961 10755 26019 10761
rect 18693 10727 18751 10733
rect 18693 10724 18705 10727
rect 16868 10696 18705 10724
rect 15197 10687 15255 10693
rect 18693 10693 18705 10696
rect 18739 10724 18751 10727
rect 22388 10724 22416 10752
rect 23382 10724 23388 10736
rect 18739 10696 18920 10724
rect 22388 10696 23388 10724
rect 18739 10693 18751 10696
rect 18693 10687 18751 10693
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 12526 10656 12532 10668
rect 12299 10628 12532 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 12526 10616 12532 10628
rect 12584 10656 12590 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12584 10628 13001 10656
rect 12584 10616 12590 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 13538 10656 13544 10668
rect 13451 10628 13544 10656
rect 12989 10619 13047 10625
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 14458 10656 14464 10668
rect 13596 10628 14464 10656
rect 13596 10616 13602 10628
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 14642 10656 14648 10668
rect 14603 10628 14648 10656
rect 14642 10616 14648 10628
rect 14700 10656 14706 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 14700 10628 16129 10656
rect 14700 10616 14706 10628
rect 16117 10625 16129 10628
rect 16163 10656 16175 10659
rect 16298 10656 16304 10668
rect 16163 10628 16304 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16298 10616 16304 10628
rect 16356 10656 16362 10668
rect 18892 10665 18920 10696
rect 23382 10684 23388 10696
rect 23440 10724 23446 10736
rect 23440 10696 23704 10724
rect 23440 10684 23446 10696
rect 17221 10659 17279 10665
rect 17221 10656 17233 10659
rect 16356 10628 17233 10656
rect 16356 10616 16362 10628
rect 17221 10625 17233 10628
rect 17267 10625 17279 10659
rect 17221 10619 17279 10625
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21910 10656 21916 10668
rect 21315 10628 21916 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 23676 10665 23704 10696
rect 23661 10659 23719 10665
rect 23661 10625 23673 10659
rect 23707 10625 23719 10659
rect 23661 10619 23719 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1486 10588 1492 10600
rect 1443 10560 1492 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 1670 10597 1676 10600
rect 1664 10588 1676 10597
rect 1631 10560 1676 10588
rect 1664 10551 1676 10560
rect 1670 10548 1676 10551
rect 1728 10548 1734 10600
rect 11330 10588 11336 10600
rect 11291 10560 11336 10588
rect 11330 10548 11336 10560
rect 11388 10588 11394 10600
rect 12618 10588 12624 10600
rect 11388 10560 12624 10588
rect 11388 10548 11394 10560
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10588 15255 10591
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15243 10560 16037 10588
rect 15243 10557 15255 10560
rect 15197 10551 15255 10557
rect 16025 10557 16037 10560
rect 16071 10588 16083 10591
rect 16666 10588 16672 10600
rect 16071 10560 16672 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 19150 10597 19156 10600
rect 19144 10588 19156 10597
rect 19111 10560 19156 10588
rect 19144 10551 19156 10560
rect 19150 10548 19156 10551
rect 19208 10548 19214 10600
rect 23934 10597 23940 10600
rect 23928 10588 23940 10597
rect 23895 10560 23940 10588
rect 23928 10551 23940 10560
rect 23934 10548 23940 10551
rect 23992 10548 23998 10600
rect 11606 10480 11612 10532
rect 11664 10520 11670 10532
rect 11885 10523 11943 10529
rect 11885 10520 11897 10523
rect 11664 10492 11897 10520
rect 11664 10480 11670 10492
rect 11885 10489 11897 10492
rect 11931 10520 11943 10523
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 11931 10492 12817 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 20901 10523 20959 10529
rect 20901 10520 20913 10523
rect 20772 10492 20913 10520
rect 20772 10480 20778 10492
rect 20901 10489 20913 10492
rect 20947 10520 20959 10523
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 20947 10492 21833 10520
rect 20947 10489 20959 10492
rect 20901 10483 20959 10489
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 12894 10452 12900 10464
rect 2832 10424 2877 10452
rect 12855 10424 12900 10452
rect 2832 10412 2838 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13596 10424 13829 10452
rect 13596 10412 13602 10424
rect 13817 10421 13829 10424
rect 13863 10452 13875 10455
rect 14366 10452 14372 10464
rect 13863 10424 14372 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15473 10455 15531 10461
rect 15473 10421 15485 10455
rect 15519 10452 15531 10455
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15519 10424 15945 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 15933 10421 15945 10424
rect 15979 10452 15991 10455
rect 16022 10452 16028 10464
rect 15979 10424 16028 10452
rect 15979 10421 15991 10424
rect 15933 10415 15991 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 20254 10452 20260 10464
rect 20215 10424 20260 10452
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 21726 10452 21732 10464
rect 21687 10424 21732 10452
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 24210 10452 24216 10464
rect 23532 10424 24216 10452
rect 23532 10412 23538 10424
rect 24210 10412 24216 10424
rect 24268 10452 24274 10464
rect 25041 10455 25099 10461
rect 25041 10452 25053 10455
rect 24268 10424 25053 10452
rect 24268 10412 24274 10424
rect 25041 10421 25053 10424
rect 25087 10421 25099 10455
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 25041 10415 25099 10421
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 13173 10251 13231 10257
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 13998 10248 14004 10260
rect 13219 10220 14004 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 13998 10208 14004 10220
rect 14056 10248 14062 10260
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14056 10220 15301 10248
rect 14056 10208 14062 10220
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 16298 10248 16304 10260
rect 16259 10220 16304 10248
rect 15289 10211 15347 10217
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16632 10220 16681 10248
rect 16632 10208 16638 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 16816 10220 18429 10248
rect 16816 10208 16822 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 18417 10211 18475 10217
rect 21266 10208 21272 10220
rect 21324 10248 21330 10260
rect 21818 10248 21824 10260
rect 21324 10220 21824 10248
rect 21324 10208 21330 10220
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 23014 10248 23020 10260
rect 22511 10220 23020 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 13541 10183 13599 10189
rect 11204 10152 12204 10180
rect 11204 10140 11210 10152
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11440 10084 11989 10112
rect 11146 9908 11152 9920
rect 11107 9880 11152 9908
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11330 9868 11336 9920
rect 11388 9908 11394 9920
rect 11440 9917 11468 10084
rect 11977 10081 11989 10084
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 12066 10044 12072 10056
rect 12027 10016 12072 10044
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12176 10053 12204 10152
rect 13541 10149 13553 10183
rect 13587 10180 13599 10183
rect 13722 10180 13728 10192
rect 13587 10152 13728 10180
rect 13587 10149 13599 10152
rect 13541 10143 13599 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 17402 10180 17408 10192
rect 17328 10152 17408 10180
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14001 10115 14059 10121
rect 14001 10112 14013 10115
rect 13872 10084 14013 10112
rect 13872 10072 13878 10084
rect 14001 10081 14013 10084
rect 14047 10081 14059 10115
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 14001 10075 14059 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10013 12219 10047
rect 14090 10044 14096 10056
rect 14051 10016 14096 10044
rect 12161 10007 12219 10013
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14240 10016 14333 10044
rect 14240 10004 14246 10016
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15620 10016 15761 10044
rect 15620 10004 15626 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16298 10044 16304 10056
rect 15979 10016 16304 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 17126 10004 17132 10056
rect 17184 10044 17190 10056
rect 17328 10053 17356 10152
rect 17402 10140 17408 10152
rect 17460 10140 17466 10192
rect 23474 10140 23480 10192
rect 23532 10180 23538 10192
rect 23722 10183 23780 10189
rect 23722 10180 23734 10183
rect 23532 10152 23734 10180
rect 23532 10140 23538 10152
rect 23722 10149 23734 10152
rect 23768 10149 23780 10183
rect 23722 10143 23780 10149
rect 18782 10112 18788 10124
rect 18743 10084 18788 10112
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 18877 10115 18935 10121
rect 18877 10081 18889 10115
rect 18923 10112 18935 10115
rect 19150 10112 19156 10124
rect 18923 10084 19156 10112
rect 18923 10081 18935 10084
rect 18877 10075 18935 10081
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 17184 10016 17325 10044
rect 17184 10004 17190 10016
rect 17313 10013 17325 10016
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 18966 10044 18972 10056
rect 17460 10016 17505 10044
rect 18927 10016 18972 10044
rect 17460 10004 17466 10016
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 21358 10044 21364 10056
rect 21319 10016 21364 10044
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21508 10016 21553 10044
rect 21508 10004 21514 10016
rect 23382 10004 23388 10056
rect 23440 10044 23446 10056
rect 23477 10047 23535 10053
rect 23477 10044 23489 10047
rect 23440 10016 23489 10044
rect 23440 10004 23446 10016
rect 23477 10013 23489 10016
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 13446 9936 13452 9988
rect 13504 9976 13510 9988
rect 14200 9976 14228 10004
rect 13504 9948 14228 9976
rect 20901 9979 20959 9985
rect 13504 9936 13510 9948
rect 20901 9945 20913 9979
rect 20947 9976 20959 9979
rect 21726 9976 21732 9988
rect 20947 9948 21732 9976
rect 20947 9945 20959 9948
rect 20901 9939 20959 9945
rect 21726 9936 21732 9948
rect 21784 9976 21790 9988
rect 21913 9979 21971 9985
rect 21913 9976 21925 9979
rect 21784 9948 21925 9976
rect 21784 9936 21790 9948
rect 21913 9945 21925 9948
rect 21959 9945 21971 9979
rect 21913 9939 21971 9945
rect 11425 9911 11483 9917
rect 11425 9908 11437 9911
rect 11388 9880 11437 9908
rect 11388 9868 11394 9880
rect 11425 9877 11437 9880
rect 11471 9877 11483 9911
rect 11425 9871 11483 9877
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12032 9880 12633 9908
rect 12032 9868 12038 9880
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 13630 9908 13636 9920
rect 13591 9880 13636 9908
rect 12621 9871 12679 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 14826 9908 14832 9920
rect 14787 9880 14832 9908
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 16850 9908 16856 9920
rect 16811 9880 16856 9908
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 18322 9908 18328 9920
rect 18187 9880 18328 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 24854 9908 24860 9920
rect 24815 9880 24860 9908
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 25314 9868 25320 9920
rect 25372 9908 25378 9920
rect 25409 9911 25467 9917
rect 25409 9908 25421 9911
rect 25372 9880 25421 9908
rect 25372 9868 25378 9880
rect 25409 9877 25421 9880
rect 25455 9877 25467 9911
rect 25409 9871 25467 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 13998 9704 14004 9716
rect 13959 9676 14004 9704
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 16117 9707 16175 9713
rect 16117 9673 16129 9707
rect 16163 9704 16175 9707
rect 16298 9704 16304 9716
rect 16163 9676 16304 9704
rect 16163 9673 16175 9676
rect 16117 9667 16175 9673
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 20714 9704 20720 9716
rect 16632 9676 17908 9704
rect 20675 9676 20720 9704
rect 16632 9664 16638 9676
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 12032 9608 13032 9636
rect 12032 9596 12038 9608
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 13004 9577 13032 9608
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 17405 9639 17463 9645
rect 17405 9636 17417 9639
rect 16724 9608 17417 9636
rect 16724 9596 16730 9608
rect 17405 9605 17417 9608
rect 17451 9605 17463 9639
rect 17880 9636 17908 9676
rect 20714 9664 20720 9676
rect 20772 9664 20778 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 21729 9707 21787 9713
rect 21729 9704 21741 9707
rect 21416 9676 21741 9704
rect 21416 9664 21422 9676
rect 21729 9673 21741 9676
rect 21775 9673 21787 9707
rect 21729 9667 21787 9673
rect 21818 9664 21824 9716
rect 21876 9704 21882 9716
rect 22097 9707 22155 9713
rect 22097 9704 22109 9707
rect 21876 9676 22109 9704
rect 21876 9664 21882 9676
rect 22097 9673 22109 9676
rect 22143 9673 22155 9707
rect 23382 9704 23388 9716
rect 23343 9676 23388 9704
rect 22097 9667 22155 9673
rect 23382 9664 23388 9676
rect 23440 9704 23446 9716
rect 23937 9707 23995 9713
rect 23937 9704 23949 9707
rect 23440 9676 23949 9704
rect 23440 9664 23446 9676
rect 23937 9673 23949 9676
rect 23983 9673 23995 9707
rect 23937 9667 23995 9673
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 17880 9608 18061 9636
rect 17405 9599 17463 9605
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 18049 9599 18107 9605
rect 12989 9571 13047 9577
rect 11848 9540 12940 9568
rect 11848 9528 11854 9540
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9692 9472 9873 9500
rect 9692 9376 9720 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10117 9503 10175 9509
rect 10117 9500 10129 9503
rect 10008 9472 10129 9500
rect 10008 9460 10014 9472
rect 10117 9469 10129 9472
rect 10163 9500 10175 9503
rect 11974 9500 11980 9512
rect 10163 9472 11980 9500
rect 10163 9469 10175 9472
rect 10117 9463 10175 9469
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12802 9500 12808 9512
rect 12176 9472 12808 9500
rect 12176 9376 12204 9472
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 12912 9509 12940 9540
rect 12989 9537 13001 9571
rect 13035 9568 13047 9571
rect 13035 9540 13676 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13078 9500 13084 9512
rect 12943 9472 13084 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13648 9500 13676 9540
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14642 9568 14648 9580
rect 13780 9540 14648 9568
rect 13780 9528 13786 9540
rect 14642 9528 14648 9540
rect 14700 9568 14706 9580
rect 14737 9571 14795 9577
rect 14737 9568 14749 9571
rect 14700 9540 14749 9568
rect 14700 9528 14706 9540
rect 14737 9537 14749 9540
rect 14783 9537 14795 9571
rect 16758 9568 16764 9580
rect 16719 9540 16764 9568
rect 14737 9531 14795 9537
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 17420 9568 17448 9599
rect 21450 9596 21456 9648
rect 21508 9596 21514 9648
rect 21634 9636 21640 9648
rect 21595 9608 21640 9636
rect 21634 9596 21640 9608
rect 21692 9596 21698 9648
rect 17678 9568 17684 9580
rect 17420 9540 17684 9568
rect 17678 9528 17684 9540
rect 17736 9568 17742 9580
rect 18230 9568 18236 9580
rect 17736 9540 18236 9568
rect 17736 9528 17742 9540
rect 18230 9528 18236 9540
rect 18288 9568 18294 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18288 9540 18521 9568
rect 18288 9528 18294 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 18874 9568 18880 9580
rect 18739 9540 18880 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 18874 9528 18880 9540
rect 18932 9568 18938 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 18932 9540 19441 9568
rect 18932 9528 18938 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 19429 9531 19487 9537
rect 20364 9540 21373 9568
rect 17034 9500 17040 9512
rect 13648 9472 17040 9500
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20162 9500 20168 9512
rect 19935 9472 20168 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20162 9460 20168 9472
rect 20220 9500 20226 9512
rect 20364 9500 20392 9540
rect 21361 9537 21373 9540
rect 21407 9568 21419 9571
rect 21468 9568 21496 9596
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 21407 9540 22477 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 23952 9568 23980 9667
rect 24121 9571 24179 9577
rect 24121 9568 24133 9571
rect 23952 9540 24133 9568
rect 22465 9531 22523 9537
rect 24121 9537 24133 9540
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 20220 9472 20392 9500
rect 20625 9503 20683 9509
rect 20220 9460 20226 9472
rect 20625 9469 20637 9503
rect 20671 9500 20683 9503
rect 21082 9500 21088 9512
rect 20671 9472 21088 9500
rect 20671 9469 20683 9472
rect 20625 9463 20683 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 24388 9503 24446 9509
rect 24388 9469 24400 9503
rect 24434 9500 24446 9503
rect 24762 9500 24768 9512
rect 24434 9472 24768 9500
rect 24434 9469 24446 9472
rect 24388 9463 24446 9469
rect 24762 9460 24768 9472
rect 24820 9460 24826 9512
rect 14826 9392 14832 9444
rect 14884 9432 14890 9444
rect 15010 9441 15016 9444
rect 15004 9432 15016 9441
rect 14884 9404 15016 9432
rect 14884 9392 14890 9404
rect 15004 9395 15016 9404
rect 15010 9392 15016 9395
rect 15068 9392 15074 9444
rect 17862 9432 17868 9444
rect 17823 9404 17868 9432
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 20257 9435 20315 9441
rect 20257 9401 20269 9435
rect 20303 9432 20315 9435
rect 20806 9432 20812 9444
rect 20303 9404 20812 9432
rect 20303 9401 20315 9404
rect 20257 9395 20315 9401
rect 20806 9392 20812 9404
rect 20864 9432 20870 9444
rect 21177 9435 21235 9441
rect 21177 9432 21189 9435
rect 20864 9404 21189 9432
rect 20864 9392 20870 9404
rect 21177 9401 21189 9404
rect 21223 9401 21235 9435
rect 23474 9432 23480 9444
rect 21177 9395 21235 9401
rect 23032 9404 23480 9432
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11146 9364 11152 9376
rect 10928 9336 11152 9364
rect 10928 9324 10934 9336
rect 11146 9324 11152 9336
rect 11204 9364 11210 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 11204 9336 11253 9364
rect 11204 9324 11210 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11790 9364 11796 9376
rect 11751 9336 11796 9364
rect 11241 9327 11299 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12802 9364 12808 9376
rect 12483 9336 12808 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13722 9364 13728 9376
rect 13683 9336 13728 9364
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14645 9367 14703 9373
rect 14645 9333 14657 9367
rect 14691 9364 14703 9367
rect 15562 9364 15568 9376
rect 14691 9336 15568 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17037 9367 17095 9373
rect 17037 9364 17049 9367
rect 16816 9336 17049 9364
rect 16816 9324 16822 9336
rect 17037 9333 17049 9336
rect 17083 9364 17095 9367
rect 17126 9364 17132 9376
rect 17083 9336 17132 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 18322 9324 18328 9376
rect 18380 9364 18386 9376
rect 18417 9367 18475 9373
rect 18417 9364 18429 9367
rect 18380 9336 18429 9364
rect 18380 9324 18386 9336
rect 18417 9333 18429 9336
rect 18463 9333 18475 9367
rect 19150 9364 19156 9376
rect 19111 9336 19156 9364
rect 18417 9327 18475 9333
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 21450 9324 21456 9376
rect 21508 9364 21514 9376
rect 21637 9367 21695 9373
rect 21637 9364 21649 9367
rect 21508 9336 21649 9364
rect 21508 9324 21514 9336
rect 21637 9333 21649 9336
rect 21683 9333 21695 9367
rect 21637 9327 21695 9333
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 23032 9373 23060 9404
rect 23474 9392 23480 9404
rect 23532 9392 23538 9444
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22336 9336 23029 9364
rect 22336 9324 22342 9336
rect 23017 9333 23029 9336
rect 23063 9333 23075 9367
rect 25498 9364 25504 9376
rect 25459 9336 25504 9364
rect 23017 9327 23075 9333
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 12584 9132 12629 9160
rect 12584 9120 12590 9132
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 12952 9132 13645 9160
rect 12952 9120 12958 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13780 9132 14105 9160
rect 13780 9120 13786 9132
rect 14093 9129 14105 9132
rect 14139 9160 14151 9163
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 14139 9132 17785 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 17773 9123 17831 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 19484 9132 19993 9160
rect 19484 9120 19490 9132
rect 19981 9129 19993 9132
rect 20027 9160 20039 9163
rect 20254 9160 20260 9172
rect 20027 9132 20260 9160
rect 20027 9129 20039 9132
rect 19981 9123 20039 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20717 9163 20775 9169
rect 20717 9129 20729 9163
rect 20763 9160 20775 9163
rect 21542 9160 21548 9172
rect 20763 9132 21548 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22152 9132 22661 9160
rect 22152 9120 22158 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 23017 9163 23075 9169
rect 23017 9129 23029 9163
rect 23063 9160 23075 9163
rect 23658 9160 23664 9172
rect 23063 9132 23664 9160
rect 23063 9129 23075 9132
rect 23017 9123 23075 9129
rect 23658 9120 23664 9132
rect 23716 9120 23722 9172
rect 24026 9120 24032 9172
rect 24084 9160 24090 9172
rect 24213 9163 24271 9169
rect 24213 9160 24225 9163
rect 24084 9132 24225 9160
rect 24084 9120 24090 9132
rect 24213 9129 24225 9132
rect 24259 9129 24271 9163
rect 24213 9123 24271 9129
rect 11057 9095 11115 9101
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 12066 9092 12072 9104
rect 11103 9064 12072 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 12066 9052 12072 9064
rect 12124 9092 12130 9104
rect 12802 9092 12808 9104
rect 12124 9064 12808 9092
rect 12124 9052 12130 9064
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 13446 9092 13452 9104
rect 13407 9064 13452 9092
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 14642 9052 14648 9104
rect 14700 9092 14706 9104
rect 14737 9095 14795 9101
rect 14737 9092 14749 9095
rect 14700 9064 14749 9092
rect 14700 9052 14706 9064
rect 14737 9061 14749 9064
rect 14783 9092 14795 9095
rect 15556 9095 15614 9101
rect 14783 9064 15332 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11405 9027 11463 9033
rect 11405 9024 11417 9027
rect 10928 8996 11417 9024
rect 10928 8984 10934 8996
rect 11405 8993 11417 8996
rect 11451 9024 11463 9027
rect 11451 8996 12204 9024
rect 11451 8993 11463 8996
rect 11405 8987 11463 8993
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 11146 8956 11152 8968
rect 9732 8928 11152 8956
rect 9732 8916 9738 8928
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 12176 8956 12204 8996
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 13170 9024 13176 9036
rect 12952 8996 13176 9024
rect 12952 8984 12958 8996
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13998 9024 14004 9036
rect 13959 8996 14004 9024
rect 13998 8984 14004 8996
rect 14056 8984 14062 9036
rect 15304 9033 15332 9064
rect 15556 9061 15568 9095
rect 15602 9092 15614 9095
rect 16206 9092 16212 9104
rect 15602 9064 16212 9092
rect 15602 9061 15614 9064
rect 15556 9055 15614 9061
rect 16206 9052 16212 9064
rect 16264 9092 16270 9104
rect 17402 9092 17408 9104
rect 16264 9064 17408 9092
rect 16264 9052 16270 9064
rect 17402 9052 17408 9064
rect 17460 9092 17466 9104
rect 17589 9095 17647 9101
rect 17589 9092 17601 9095
rect 17460 9064 17601 9092
rect 17460 9052 17466 9064
rect 17589 9061 17601 9064
rect 17635 9061 17647 9095
rect 17589 9055 17647 9061
rect 24121 9095 24179 9101
rect 24121 9061 24133 9095
rect 24167 9092 24179 9095
rect 24762 9092 24768 9104
rect 24167 9064 24768 9092
rect 24167 9061 24179 9064
rect 24121 9055 24179 9061
rect 15289 9027 15347 9033
rect 15289 8993 15301 9027
rect 15335 8993 15347 9027
rect 18138 9024 18144 9036
rect 18099 8996 18144 9024
rect 15289 8987 15347 8993
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 19392 8996 19441 9024
rect 19392 8984 19398 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 21453 9027 21511 9033
rect 21453 8993 21465 9027
rect 21499 9024 21511 9027
rect 21910 9024 21916 9036
rect 21499 8996 21916 9024
rect 21499 8993 21511 8996
rect 21453 8987 21511 8993
rect 21910 8984 21916 8996
rect 21968 8984 21974 9036
rect 14185 8959 14243 8965
rect 14185 8956 14197 8959
rect 12176 8928 14197 8956
rect 14185 8925 14197 8928
rect 14231 8956 14243 8959
rect 14366 8956 14372 8968
rect 14231 8928 14372 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17770 8956 17776 8968
rect 17092 8928 17776 8956
rect 17092 8916 17098 8928
rect 17770 8916 17776 8928
rect 17828 8956 17834 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 17828 8928 18337 8956
rect 17828 8916 17834 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 21729 8959 21787 8965
rect 21729 8925 21741 8959
rect 21775 8956 21787 8959
rect 22186 8956 22192 8968
rect 21775 8928 22192 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8956 22615 8959
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 22603 8928 23121 8956
rect 22603 8925 22615 8928
rect 22557 8919 22615 8925
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23290 8956 23296 8968
rect 23203 8928 23296 8956
rect 23109 8919 23167 8925
rect 16574 8848 16580 8900
rect 16632 8888 16638 8900
rect 17218 8888 17224 8900
rect 16632 8860 17224 8888
rect 16632 8848 16638 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 19613 8891 19671 8897
rect 19613 8857 19625 8891
rect 19659 8888 19671 8891
rect 20162 8888 20168 8900
rect 19659 8860 20168 8888
rect 19659 8857 19671 8860
rect 19613 8851 19671 8857
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 21085 8891 21143 8897
rect 21085 8857 21097 8891
rect 21131 8888 21143 8891
rect 22572 8888 22600 8919
rect 23290 8916 23296 8928
rect 23348 8956 23354 8968
rect 24136 8956 24164 9055
rect 24762 9052 24768 9064
rect 24820 9052 24826 9104
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 24854 9024 24860 9036
rect 24627 8996 24860 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 24670 8956 24676 8968
rect 23348 8928 24164 8956
rect 24631 8928 24676 8956
rect 23348 8916 23354 8928
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 24762 8916 24768 8968
rect 24820 8956 24826 8968
rect 24820 8928 24865 8956
rect 24820 8916 24826 8928
rect 21131 8860 22600 8888
rect 24688 8888 24716 8916
rect 25225 8891 25283 8897
rect 25225 8888 25237 8891
rect 24688 8860 25237 8888
rect 21131 8857 21143 8860
rect 21085 8851 21143 8857
rect 25225 8857 25237 8860
rect 25271 8857 25283 8891
rect 25225 8851 25283 8857
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 15470 8820 15476 8832
rect 13412 8792 15476 8820
rect 13412 8780 13418 8792
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 16666 8820 16672 8832
rect 16627 8792 16672 8820
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 18782 8820 18788 8832
rect 18743 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 22189 8823 22247 8829
rect 22189 8789 22201 8823
rect 22235 8820 22247 8823
rect 22370 8820 22376 8832
rect 22235 8792 22376 8820
rect 22235 8789 22247 8792
rect 22189 8783 22247 8789
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 23566 8780 23572 8832
rect 23624 8820 23630 8832
rect 24762 8820 24768 8832
rect 23624 8792 24768 8820
rect 23624 8780 23630 8792
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8616 11210 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11204 8588 12081 8616
rect 11204 8576 11210 8588
rect 12069 8585 12081 8588
rect 12115 8616 12127 8619
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12115 8588 12173 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 14366 8616 14372 8628
rect 14327 8588 14372 8616
rect 12161 8579 12219 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 14700 8588 14749 8616
rect 14700 8576 14706 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 14737 8579 14795 8585
rect 11330 8480 11336 8492
rect 11291 8452 11336 8480
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 14752 8480 14780 8579
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17497 8619 17555 8625
rect 17497 8585 17509 8619
rect 17543 8616 17555 8619
rect 18138 8616 18144 8628
rect 17543 8588 18144 8616
rect 17543 8585 17555 8588
rect 17497 8579 17555 8585
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 20772 8588 21373 8616
rect 20772 8576 20778 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 22244 8588 22385 8616
rect 22244 8576 22250 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22373 8579 22431 8585
rect 23017 8619 23075 8625
rect 23017 8585 23029 8619
rect 23063 8616 23075 8619
rect 23290 8616 23296 8628
rect 23063 8588 23296 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23290 8576 23296 8588
rect 23348 8576 23354 8628
rect 23474 8616 23480 8628
rect 23435 8588 23480 8616
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 24820 8588 25513 8616
rect 24820 8576 24826 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 25501 8579 25559 8585
rect 21910 8548 21916 8560
rect 21871 8520 21916 8548
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 22278 8508 22284 8560
rect 22336 8548 22342 8560
rect 22649 8551 22707 8557
rect 22649 8548 22661 8551
rect 22336 8520 22661 8548
rect 22336 8508 22342 8520
rect 22649 8517 22661 8520
rect 22695 8517 22707 8551
rect 22649 8511 22707 8517
rect 14918 8480 14924 8492
rect 11931 8452 12572 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12544 8424 12572 8452
rect 14752 8452 14924 8480
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8412 12127 8415
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12115 8384 12449 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12452 8344 12480 8375
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12693 8415 12751 8421
rect 12693 8412 12705 8415
rect 12584 8384 12705 8412
rect 12584 8372 12590 8384
rect 12693 8381 12705 8384
rect 12739 8381 12751 8415
rect 14090 8412 14096 8424
rect 12693 8375 12751 8381
rect 12820 8384 14096 8412
rect 12820 8344 12848 8384
rect 14090 8372 14096 8384
rect 14148 8412 14154 8424
rect 14752 8412 14780 8452
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 17920 8452 18705 8480
rect 17920 8440 17926 8452
rect 18693 8449 18705 8452
rect 18739 8480 18751 8483
rect 18782 8480 18788 8492
rect 18739 8452 18788 8480
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 23492 8480 23520 8576
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 23492 8452 24133 8480
rect 24121 8449 24133 8452
rect 24167 8449 24179 8483
rect 24121 8443 24179 8449
rect 14148 8384 14780 8412
rect 17773 8415 17831 8421
rect 14148 8372 14154 8384
rect 17773 8381 17785 8415
rect 17819 8412 17831 8415
rect 18322 8412 18328 8424
rect 17819 8384 18328 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 18322 8372 18328 8384
rect 18380 8412 18386 8424
rect 18506 8412 18512 8424
rect 18380 8384 18512 8412
rect 18380 8372 18386 8384
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 20254 8421 20260 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20248 8412 20260 8421
rect 20027 8384 20061 8412
rect 20215 8384 20260 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20248 8375 20260 8384
rect 15188 8347 15246 8353
rect 15188 8344 15200 8347
rect 12452 8316 12848 8344
rect 13832 8316 15200 8344
rect 13832 8285 13860 8316
rect 15188 8313 15200 8316
rect 15234 8344 15246 8347
rect 15838 8344 15844 8356
rect 15234 8316 15844 8344
rect 15234 8313 15246 8316
rect 15188 8307 15246 8313
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 17954 8304 17960 8356
rect 18012 8344 18018 8356
rect 18417 8347 18475 8353
rect 18417 8344 18429 8347
rect 18012 8316 18429 8344
rect 18012 8304 18018 8316
rect 18417 8313 18429 8316
rect 18463 8344 18475 8347
rect 18690 8344 18696 8356
rect 18463 8316 18696 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18690 8304 18696 8316
rect 18748 8344 18754 8356
rect 19061 8347 19119 8353
rect 19061 8344 19073 8347
rect 18748 8316 19073 8344
rect 18748 8304 18754 8316
rect 19061 8313 19073 8316
rect 19107 8313 19119 8347
rect 19061 8307 19119 8313
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 19392 8316 19441 8344
rect 19392 8304 19398 8316
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 19429 8307 19487 8313
rect 19889 8347 19947 8353
rect 19889 8313 19901 8347
rect 19935 8344 19947 8347
rect 19996 8344 20024 8375
rect 20254 8372 20260 8375
rect 20312 8372 20318 8424
rect 22462 8412 22468 8424
rect 22423 8384 22468 8412
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 24026 8412 24032 8424
rect 23939 8384 24032 8412
rect 24026 8372 24032 8384
rect 24084 8412 24090 8424
rect 24854 8412 24860 8424
rect 24084 8384 24860 8412
rect 24084 8372 24090 8384
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 20070 8344 20076 8356
rect 19935 8316 20076 8344
rect 19935 8313 19947 8316
rect 19889 8307 19947 8313
rect 20070 8304 20076 8316
rect 20128 8344 20134 8356
rect 20530 8344 20536 8356
rect 20128 8316 20536 8344
rect 20128 8304 20134 8316
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 21726 8304 21732 8356
rect 21784 8344 21790 8356
rect 24388 8347 24446 8353
rect 24388 8344 24400 8347
rect 21784 8316 24400 8344
rect 21784 8304 21790 8316
rect 24388 8313 24400 8316
rect 24434 8344 24446 8347
rect 24578 8344 24584 8356
rect 24434 8316 24584 8344
rect 24434 8313 24446 8316
rect 24388 8307 24446 8313
rect 24578 8304 24584 8316
rect 24636 8344 24642 8356
rect 25498 8344 25504 8356
rect 24636 8316 25504 8344
rect 24636 8304 24642 8316
rect 25498 8304 25504 8316
rect 25556 8304 25562 8356
rect 13817 8279 13875 8285
rect 13817 8245 13829 8279
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 16301 8279 16359 8285
rect 16301 8276 16313 8279
rect 16264 8248 16313 8276
rect 16264 8236 16270 8248
rect 16301 8245 16313 8248
rect 16347 8245 16359 8279
rect 18046 8276 18052 8288
rect 18007 8248 18052 8276
rect 16301 8239 16359 8245
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 13541 8075 13599 8081
rect 12115 8044 12940 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 11974 8004 11980 8016
rect 11935 7976 11980 8004
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 12912 8004 12940 8044
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13722 8072 13728 8084
rect 13587 8044 13728 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14001 8075 14059 8081
rect 14001 8041 14013 8075
rect 14047 8072 14059 8075
rect 14182 8072 14188 8084
rect 14047 8044 14188 8072
rect 14047 8041 14059 8044
rect 14001 8035 14059 8041
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 14918 8072 14924 8084
rect 14879 8044 14924 8072
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 16482 8072 16488 8084
rect 15335 8044 16488 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17736 8044 17785 8072
rect 17736 8032 17742 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 18138 8072 18144 8084
rect 18099 8044 18144 8072
rect 17773 8035 17831 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 21082 8072 21088 8084
rect 21043 8044 21088 8072
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 24578 8032 24584 8084
rect 24636 8072 24642 8084
rect 24636 8044 24681 8072
rect 24636 8032 24642 8044
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 24949 8075 25007 8081
rect 24949 8072 24961 8075
rect 24912 8044 24961 8072
rect 24912 8032 24918 8044
rect 24949 8041 24961 8044
rect 24995 8041 25007 8075
rect 24949 8035 25007 8041
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 12492 7976 12537 8004
rect 12912 7976 14105 8004
rect 12492 7964 12498 7976
rect 14093 7973 14105 7976
rect 14139 8004 14151 8007
rect 14642 8004 14648 8016
rect 14139 7976 14648 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15838 8004 15844 8016
rect 15751 7976 15844 8004
rect 15838 7964 15844 7976
rect 15896 8004 15902 8016
rect 16298 8004 16304 8016
rect 15896 7976 16304 8004
rect 15896 7964 15902 7976
rect 16298 7964 16304 7976
rect 16356 8004 16362 8016
rect 23382 8004 23388 8016
rect 16356 7976 17264 8004
rect 16356 7964 16362 7976
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13998 7936 14004 7948
rect 13219 7908 14004 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 16942 7936 16948 7948
rect 16903 7908 16948 7936
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 12526 7868 12532 7880
rect 12487 7840 12532 7868
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 12802 7868 12808 7880
rect 12759 7840 12808 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14826 7868 14832 7880
rect 14323 7840 14832 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7868 17095 7871
rect 17126 7868 17132 7880
rect 17083 7840 17132 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17236 7877 17264 7976
rect 22664 7976 23388 8004
rect 18506 7936 18512 7948
rect 18467 7908 18512 7936
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 20898 7896 20904 7948
rect 20956 7936 20962 7948
rect 22664 7945 22692 7976
rect 23382 7964 23388 7976
rect 23440 7964 23446 8016
rect 22922 7945 22928 7948
rect 21453 7939 21511 7945
rect 21453 7936 21465 7939
rect 20956 7908 21465 7936
rect 20956 7896 20962 7908
rect 21453 7905 21465 7908
rect 21499 7905 21511 7939
rect 21453 7899 21511 7905
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7905 22707 7939
rect 22916 7936 22928 7945
rect 22883 7908 22928 7936
rect 22649 7899 22707 7905
rect 22916 7899 22928 7908
rect 22922 7896 22928 7899
rect 22980 7896 22986 7948
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17862 7868 17868 7880
rect 17267 7840 17868 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18598 7868 18604 7880
rect 18559 7840 18604 7868
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 19702 7868 19708 7880
rect 19663 7840 19708 7868
rect 18693 7831 18751 7837
rect 12820 7800 12848 7828
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 12820 7772 16129 7800
rect 16117 7769 16129 7772
rect 16163 7800 16175 7803
rect 16206 7800 16212 7812
rect 16163 7772 16212 7800
rect 16163 7769 16175 7772
rect 16117 7763 16175 7769
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 16574 7800 16580 7812
rect 16535 7772 16580 7800
rect 16574 7760 16580 7772
rect 16632 7760 16638 7812
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 18708 7800 18736 7831
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 21542 7868 21548 7880
rect 21503 7840 21548 7868
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 21726 7828 21732 7880
rect 21784 7868 21790 7880
rect 21784 7840 21829 7868
rect 21784 7828 21790 7840
rect 17828 7772 18736 7800
rect 20717 7803 20775 7809
rect 17828 7760 17834 7772
rect 20717 7769 20729 7803
rect 20763 7800 20775 7803
rect 21744 7800 21772 7828
rect 20763 7772 21772 7800
rect 20763 7769 20775 7772
rect 20717 7763 20775 7769
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22462 7800 22468 7812
rect 22152 7772 22468 7800
rect 22152 7760 22158 7772
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 13633 7735 13691 7741
rect 13633 7732 13645 7735
rect 12676 7704 13645 7732
rect 12676 7692 12682 7704
rect 13633 7701 13645 7704
rect 13679 7701 13691 7735
rect 13633 7695 13691 7701
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19392 7704 19441 7732
rect 19392 7692 19398 7704
rect 19429 7701 19441 7704
rect 19475 7732 19487 7735
rect 20622 7732 20628 7744
rect 19475 7704 20628 7732
rect 19475 7701 19487 7704
rect 19429 7695 19487 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 22186 7732 22192 7744
rect 22147 7704 22192 7732
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22646 7692 22652 7744
rect 22704 7732 22710 7744
rect 24029 7735 24087 7741
rect 24029 7732 24041 7735
rect 22704 7704 24041 7732
rect 22704 7692 22710 7704
rect 24029 7701 24041 7704
rect 24075 7701 24087 7735
rect 24029 7695 24087 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 12434 7528 12440 7540
rect 11563 7500 12440 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13538 7528 13544 7540
rect 13412 7500 13544 7528
rect 13412 7488 13418 7500
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14884 7500 15025 7528
rect 14884 7488 14890 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 17000 7500 17417 7528
rect 17000 7488 17006 7500
rect 17405 7497 17417 7500
rect 17451 7528 17463 7531
rect 17494 7528 17500 7540
rect 17451 7500 17500 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17770 7528 17776 7540
rect 17731 7500 17776 7528
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18506 7528 18512 7540
rect 18467 7500 18512 7528
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 18782 7528 18788 7540
rect 18656 7500 18788 7528
rect 18656 7488 18662 7500
rect 18782 7488 18788 7500
rect 18840 7528 18846 7540
rect 18877 7531 18935 7537
rect 18877 7528 18889 7531
rect 18840 7500 18889 7528
rect 18840 7488 18846 7500
rect 18877 7497 18889 7500
rect 18923 7497 18935 7531
rect 18877 7491 18935 7497
rect 19337 7531 19395 7537
rect 19337 7497 19349 7531
rect 19383 7528 19395 7531
rect 20070 7528 20076 7540
rect 19383 7500 20076 7528
rect 19383 7497 19395 7500
rect 19337 7491 19395 7497
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 12802 7460 12808 7472
rect 11931 7432 12808 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 12802 7420 12808 7432
rect 12860 7420 12866 7472
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 14458 7460 14464 7472
rect 13964 7432 14464 7460
rect 13964 7420 13970 7432
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 16025 7463 16083 7469
rect 16025 7460 16037 7463
rect 15252 7432 16037 7460
rect 15252 7420 15258 7432
rect 16025 7429 16037 7432
rect 16071 7429 16083 7463
rect 16025 7423 16083 7429
rect 19444 7404 19472 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 21450 7488 21456 7540
rect 21508 7528 21514 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21508 7500 21833 7528
rect 21508 7488 21514 7500
rect 21821 7497 21833 7500
rect 21867 7528 21879 7531
rect 22646 7528 22652 7540
rect 21867 7500 22652 7528
rect 21867 7497 21879 7500
rect 21821 7491 21879 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23109 7531 23167 7537
rect 23109 7528 23121 7531
rect 22796 7500 23121 7528
rect 22796 7488 22802 7500
rect 23109 7497 23121 7500
rect 23155 7528 23167 7531
rect 23382 7528 23388 7540
rect 23155 7500 23388 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 22370 7420 22376 7472
rect 22428 7460 22434 7472
rect 23661 7463 23719 7469
rect 23661 7460 23673 7463
rect 22428 7432 23673 7460
rect 22428 7420 22434 7432
rect 23661 7429 23673 7432
rect 23707 7429 23719 7463
rect 23661 7423 23719 7429
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12676 7364 13001 7392
rect 12676 7352 12682 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 12989 7355 13047 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 16577 7395 16635 7401
rect 16577 7392 16589 7395
rect 15896 7364 16589 7392
rect 15896 7352 15902 7364
rect 16577 7361 16589 7364
rect 16623 7361 16635 7395
rect 19426 7392 19432 7404
rect 19339 7364 19432 7392
rect 16577 7355 16635 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 22244 7364 22477 7392
rect 22244 7352 22250 7364
rect 22465 7361 22477 7364
rect 22511 7361 22523 7395
rect 22646 7392 22652 7404
rect 22607 7364 22652 7392
rect 22465 7355 22523 7361
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 24118 7352 24124 7404
rect 24176 7392 24182 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 24176 7364 24317 7392
rect 24176 7352 24182 7364
rect 24305 7361 24317 7364
rect 24351 7392 24363 7395
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24351 7364 25053 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 12894 7324 12900 7336
rect 12807 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7324 12958 7336
rect 13630 7324 13636 7336
rect 12952 7296 13636 7324
rect 12952 7284 12958 7296
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13872 7296 13921 7324
rect 13872 7284 13878 7296
rect 13909 7293 13921 7296
rect 13955 7324 13967 7327
rect 14274 7324 14280 7336
rect 13955 7296 14280 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 14274 7284 14280 7296
rect 14332 7324 14338 7336
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 14332 7296 14381 7324
rect 14332 7284 14338 7296
rect 14369 7293 14381 7296
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 15654 7324 15660 7336
rect 14507 7296 15660 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 12253 7259 12311 7265
rect 12253 7225 12265 7259
rect 12299 7256 12311 7259
rect 12802 7256 12808 7268
rect 12299 7228 12808 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 12802 7216 12808 7228
rect 12860 7216 12866 7268
rect 13541 7259 13599 7265
rect 13541 7225 13553 7259
rect 13587 7256 13599 7259
rect 14476 7256 14504 7287
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 22370 7324 22376 7336
rect 22331 7296 22376 7324
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 13587 7228 14504 7256
rect 15565 7259 15623 7265
rect 13587 7225 13599 7228
rect 13541 7219 13599 7225
rect 15565 7225 15577 7259
rect 15611 7256 15623 7259
rect 15611 7228 16528 7256
rect 15611 7225 15623 7228
rect 15565 7219 15623 7225
rect 16500 7200 16528 7228
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 19674 7259 19732 7265
rect 19674 7256 19686 7259
rect 19392 7228 19686 7256
rect 19392 7216 19398 7228
rect 19674 7225 19686 7228
rect 19720 7225 19732 7259
rect 19674 7219 19732 7225
rect 24029 7259 24087 7265
rect 24029 7225 24041 7259
rect 24075 7256 24087 7259
rect 24765 7259 24823 7265
rect 24765 7256 24777 7259
rect 24075 7228 24777 7256
rect 24075 7225 24087 7228
rect 24029 7219 24087 7225
rect 24765 7225 24777 7228
rect 24811 7256 24823 7259
rect 25225 7259 25283 7265
rect 25225 7256 25237 7259
rect 24811 7228 25237 7256
rect 24811 7225 24823 7228
rect 24765 7219 24823 7225
rect 25225 7225 25237 7228
rect 25271 7225 25283 7259
rect 25225 7219 25283 7225
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 13354 7188 13360 7200
rect 12483 7160 13360 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13906 7148 13912 7200
rect 13964 7188 13970 7200
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13964 7160 14013 7188
rect 13964 7148 13970 7160
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 15838 7188 15844 7200
rect 15799 7160 15844 7188
rect 14001 7151 14059 7157
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16390 7188 16396 7200
rect 16351 7160 16396 7188
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 17129 7191 17187 7197
rect 16540 7160 16585 7188
rect 16540 7148 16546 7160
rect 17129 7157 17141 7191
rect 17175 7188 17187 7191
rect 17218 7188 17224 7200
rect 17175 7160 17224 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 21453 7191 21511 7197
rect 21453 7157 21465 7191
rect 21499 7188 21511 7191
rect 21542 7188 21548 7200
rect 21499 7160 21548 7188
rect 21499 7157 21511 7160
rect 21453 7151 21511 7157
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 22002 7188 22008 7200
rect 21963 7160 22008 7188
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 23477 7191 23535 7197
rect 23477 7157 23489 7191
rect 23523 7188 23535 7191
rect 24121 7191 24179 7197
rect 24121 7188 24133 7191
rect 23523 7160 24133 7188
rect 23523 7157 23535 7160
rect 23477 7151 23535 7157
rect 24121 7157 24133 7160
rect 24167 7188 24179 7191
rect 24670 7188 24676 7200
rect 24167 7160 24676 7188
rect 24167 7157 24179 7160
rect 24121 7151 24179 7157
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12618 6984 12624 6996
rect 12483 6956 12624 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 12894 6984 12900 6996
rect 12855 6956 12900 6984
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 14642 6984 14648 6996
rect 14603 6956 14648 6984
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15620 6956 15669 6984
rect 15620 6944 15626 6956
rect 15657 6953 15669 6956
rect 15703 6984 15715 6987
rect 16206 6984 16212 6996
rect 15703 6956 16212 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 16298 6944 16304 6996
rect 16356 6984 16362 6996
rect 16485 6987 16543 6993
rect 16485 6984 16497 6987
rect 16356 6956 16497 6984
rect 16356 6944 16362 6956
rect 16485 6953 16497 6956
rect 16531 6953 16543 6987
rect 16485 6947 16543 6953
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18104 6956 18889 6984
rect 18104 6944 18110 6956
rect 18877 6953 18889 6956
rect 18923 6984 18935 6987
rect 18966 6984 18972 6996
rect 18923 6956 18972 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 18966 6944 18972 6956
rect 19024 6944 19030 6996
rect 22649 6987 22707 6993
rect 22649 6953 22661 6987
rect 22695 6984 22707 6987
rect 22922 6984 22928 6996
rect 22695 6956 22928 6984
rect 22695 6953 22707 6956
rect 22649 6947 22707 6953
rect 12526 6916 12532 6928
rect 12360 6888 12532 6916
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12360 6848 12388 6888
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 13630 6916 13636 6928
rect 13591 6888 13636 6916
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 16390 6916 16396 6928
rect 15120 6888 16396 6916
rect 15120 6857 15148 6888
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 17313 6919 17371 6925
rect 17313 6885 17325 6919
rect 17359 6916 17371 6919
rect 17678 6916 17684 6928
rect 17359 6888 17684 6916
rect 17359 6885 17371 6888
rect 17313 6879 17371 6885
rect 17678 6876 17684 6888
rect 17736 6876 17742 6928
rect 20346 6876 20352 6928
rect 20404 6876 20410 6928
rect 21545 6919 21603 6925
rect 21545 6885 21557 6919
rect 21591 6916 21603 6919
rect 21634 6916 21640 6928
rect 21591 6888 21640 6916
rect 21591 6885 21603 6888
rect 21545 6879 21603 6885
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 22002 6876 22008 6928
rect 22060 6916 22066 6928
rect 22094 6916 22100 6928
rect 22060 6888 22100 6916
rect 22060 6876 22066 6888
rect 22094 6876 22100 6888
rect 22152 6876 22158 6928
rect 12207 6820 12388 6848
rect 15105 6851 15163 6857
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 15105 6817 15117 6851
rect 15151 6817 15163 6851
rect 15746 6848 15752 6860
rect 15707 6820 15752 6848
rect 15105 6811 15163 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17460 6820 17505 6848
rect 17460 6808 17466 6820
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 18969 6851 19027 6857
rect 18969 6848 18981 6851
rect 18932 6820 18981 6848
rect 18932 6808 18938 6820
rect 18969 6817 18981 6820
rect 19015 6817 19027 6851
rect 18969 6811 19027 6817
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13740 6712 13768 6743
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 15930 6780 15936 6792
rect 13872 6752 13917 6780
rect 15891 6752 15936 6780
rect 13872 6740 13878 6752
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 17586 6780 17592 6792
rect 17547 6752 17592 6780
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 19153 6783 19211 6789
rect 19153 6749 19165 6783
rect 19199 6780 19211 6783
rect 19981 6783 20039 6789
rect 19981 6780 19993 6783
rect 19199 6752 19993 6780
rect 19199 6749 19211 6752
rect 19153 6743 19211 6749
rect 19981 6749 19993 6752
rect 20027 6749 20039 6783
rect 20364 6780 20392 6876
rect 22278 6848 22284 6860
rect 22239 6820 22284 6848
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 21637 6783 21695 6789
rect 21637 6780 21649 6783
rect 20364 6752 21649 6780
rect 19981 6743 20039 6749
rect 21637 6749 21649 6752
rect 21683 6780 21695 6783
rect 21726 6780 21732 6792
rect 21683 6752 21732 6780
rect 21683 6749 21695 6752
rect 21637 6743 21695 6749
rect 14182 6712 14188 6724
rect 13740 6684 14188 6712
rect 14182 6672 14188 6684
rect 14240 6712 14246 6724
rect 15289 6715 15347 6721
rect 15289 6712 15301 6715
rect 14240 6684 15301 6712
rect 14240 6672 14246 6684
rect 15289 6681 15301 6684
rect 15335 6681 15347 6715
rect 15289 6675 15347 6681
rect 16853 6715 16911 6721
rect 16853 6681 16865 6715
rect 16899 6712 16911 6715
rect 17604 6712 17632 6740
rect 18506 6712 18512 6724
rect 16899 6684 17632 6712
rect 18467 6684 18512 6712
rect 16899 6681 16911 6684
rect 16853 6675 16911 6681
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 18598 6672 18604 6724
rect 18656 6712 18662 6724
rect 19168 6712 19196 6743
rect 21726 6740 21732 6752
rect 21784 6740 21790 6792
rect 21821 6783 21879 6789
rect 21821 6749 21833 6783
rect 21867 6780 21879 6783
rect 22094 6780 22100 6792
rect 21867 6752 22100 6780
rect 21867 6749 21879 6752
rect 21821 6743 21879 6749
rect 22094 6740 22100 6752
rect 22152 6780 22158 6792
rect 22664 6780 22692 6947
rect 22922 6944 22928 6956
rect 22980 6984 22986 6996
rect 24118 6984 24124 6996
rect 22980 6956 24124 6984
rect 22980 6944 22986 6956
rect 24118 6944 24124 6956
rect 24176 6944 24182 6996
rect 23008 6919 23066 6925
rect 23008 6885 23020 6919
rect 23054 6916 23066 6919
rect 23106 6916 23112 6928
rect 23054 6888 23112 6916
rect 23054 6885 23066 6888
rect 23008 6879 23066 6885
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 22738 6808 22744 6860
rect 22796 6848 22802 6860
rect 25222 6848 25228 6860
rect 22796 6820 22841 6848
rect 25183 6820 25228 6848
rect 22796 6808 22802 6820
rect 25222 6808 25228 6820
rect 25280 6808 25286 6860
rect 22152 6752 22692 6780
rect 22152 6740 22158 6752
rect 20806 6712 20812 6724
rect 18656 6684 19196 6712
rect 19720 6684 20812 6712
rect 18656 6672 18662 6684
rect 19720 6656 19748 6684
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 21177 6715 21235 6721
rect 21177 6681 21189 6715
rect 21223 6712 21235 6715
rect 21910 6712 21916 6724
rect 21223 6684 21916 6712
rect 21223 6681 21235 6684
rect 21177 6675 21235 6681
rect 21910 6672 21916 6684
rect 21968 6672 21974 6724
rect 12894 6604 12900 6656
rect 12952 6644 12958 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 12952 6616 13277 6644
rect 12952 6604 12958 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 14550 6644 14556 6656
rect 14415 6616 14556 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 14550 6604 14556 6616
rect 14608 6644 14614 6656
rect 15930 6644 15936 6656
rect 14608 6616 15936 6644
rect 14608 6604 14614 6616
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16945 6647 17003 6653
rect 16945 6613 16957 6647
rect 16991 6644 17003 6647
rect 17126 6644 17132 6656
rect 16991 6616 17132 6644
rect 16991 6613 17003 6616
rect 16945 6607 17003 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 18138 6644 18144 6656
rect 18099 6616 18144 6644
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 19702 6644 19708 6656
rect 19663 6616 19708 6644
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 20898 6644 20904 6656
rect 20763 6616 20904 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 25406 6644 25412 6656
rect 25367 6616 25412 6644
rect 25406 6604 25412 6616
rect 25464 6604 25470 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 14148 6412 14565 6440
rect 14148 6400 14154 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 15746 6440 15752 6452
rect 14553 6403 14611 6409
rect 15488 6412 15752 6440
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 13596 6344 13768 6372
rect 13596 6332 13602 6344
rect 13740 6313 13768 6344
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 13725 6307 13783 6313
rect 11931 6276 13676 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 13648 6177 13676 6276
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 13814 6304 13820 6316
rect 13771 6276 13820 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 13814 6264 13820 6276
rect 13872 6304 13878 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13872 6276 14197 6304
rect 13872 6264 13878 6276
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14568 6304 14596 6403
rect 15013 6375 15071 6381
rect 15013 6341 15025 6375
rect 15059 6372 15071 6375
rect 15488 6372 15516 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 18874 6400 18880 6452
rect 18932 6440 18938 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18932 6412 19073 6440
rect 18932 6400 18938 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19426 6440 19432 6452
rect 19387 6412 19432 6440
rect 19061 6403 19119 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 21726 6400 21732 6452
rect 21784 6440 21790 6452
rect 21913 6443 21971 6449
rect 21913 6440 21925 6443
rect 21784 6412 21925 6440
rect 21784 6400 21790 6412
rect 21913 6409 21925 6412
rect 21959 6409 21971 6443
rect 22738 6440 22744 6452
rect 22699 6412 22744 6440
rect 21913 6403 21971 6409
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 24026 6440 24032 6452
rect 23987 6412 24032 6440
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 25222 6440 25228 6452
rect 25183 6412 25228 6440
rect 25222 6400 25228 6412
rect 25280 6400 25286 6452
rect 15059 6344 15516 6372
rect 15059 6341 15071 6344
rect 15013 6335 15071 6341
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 14568 6276 15485 6304
rect 14185 6267 14243 6273
rect 15473 6273 15485 6276
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 15488 6236 15516 6267
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17644 6276 18705 6304
rect 17644 6264 17650 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 19058 6304 19064 6316
rect 18739 6276 19064 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 19058 6264 19064 6276
rect 19116 6264 19122 6316
rect 19444 6304 19472 6400
rect 21634 6372 21640 6384
rect 21595 6344 21640 6372
rect 21634 6332 21640 6344
rect 21692 6332 21698 6384
rect 24044 6372 24072 6400
rect 24486 6372 24492 6384
rect 24044 6344 24492 6372
rect 24486 6332 24492 6344
rect 24544 6332 24550 6384
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19444 6276 19625 6304
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 24765 6307 24823 6313
rect 24765 6304 24777 6307
rect 24728 6276 24777 6304
rect 24728 6264 24734 6276
rect 24765 6273 24777 6276
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 16942 6236 16948 6248
rect 15488 6208 16948 6236
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18414 6236 18420 6248
rect 17911 6208 18420 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 19702 6196 19708 6248
rect 19760 6236 19766 6248
rect 19869 6239 19927 6245
rect 19869 6236 19881 6239
rect 19760 6208 19881 6236
rect 19760 6196 19766 6208
rect 19869 6205 19881 6208
rect 19915 6205 19927 6239
rect 19869 6199 19927 6205
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 22278 6236 22284 6248
rect 22143 6208 22284 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 12989 6171 13047 6177
rect 12989 6168 13001 6171
rect 11388 6140 13001 6168
rect 11388 6128 11394 6140
rect 12989 6137 13001 6140
rect 13035 6168 13047 6171
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 13035 6140 13553 6168
rect 13035 6137 13047 6140
rect 12989 6131 13047 6137
rect 13541 6137 13553 6140
rect 13587 6137 13599 6171
rect 13541 6131 13599 6137
rect 13633 6171 13691 6177
rect 13633 6137 13645 6171
rect 13679 6168 13691 6171
rect 13722 6168 13728 6180
rect 13679 6140 13728 6168
rect 13679 6137 13691 6140
rect 13633 6131 13691 6137
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 15740 6171 15798 6177
rect 15740 6137 15752 6171
rect 15786 6168 15798 6171
rect 16390 6168 16396 6180
rect 15786 6140 16396 6168
rect 15786 6137 15798 6140
rect 15740 6131 15798 6137
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 23477 6171 23535 6177
rect 23477 6137 23489 6171
rect 23523 6168 23535 6171
rect 24581 6171 24639 6177
rect 24581 6168 24593 6171
rect 23523 6140 24593 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 24581 6137 24593 6140
rect 24627 6168 24639 6171
rect 25130 6168 25136 6180
rect 24627 6140 25136 6168
rect 24627 6137 24639 6140
rect 24581 6131 24639 6137
rect 25130 6128 25136 6140
rect 25188 6128 25194 6180
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12621 6103 12679 6109
rect 12621 6100 12633 6103
rect 12584 6072 12633 6100
rect 12584 6060 12590 6072
rect 12621 6069 12633 6072
rect 12667 6069 12679 6103
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 12621 6063 12679 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 15381 6103 15439 6109
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15562 6100 15568 6112
rect 15427 6072 15568 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15562 6060 15568 6072
rect 15620 6100 15626 6112
rect 16206 6100 16212 6112
rect 15620 6072 16212 6100
rect 15620 6060 15626 6072
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16850 6100 16856 6112
rect 16811 6072 16856 6100
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 17497 6103 17555 6109
rect 17497 6069 17509 6103
rect 17543 6100 17555 6103
rect 17678 6100 17684 6112
rect 17543 6072 17684 6100
rect 17543 6069 17555 6072
rect 17497 6063 17555 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 18012 6072 18061 6100
rect 18012 6060 18018 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18506 6100 18512 6112
rect 18196 6072 18512 6100
rect 18196 6060 18202 6072
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 20990 6100 20996 6112
rect 20951 6072 20996 6100
rect 20990 6060 20996 6072
rect 21048 6060 21054 6112
rect 22281 6103 22339 6109
rect 22281 6069 22293 6103
rect 22327 6100 22339 6103
rect 22646 6100 22652 6112
rect 22327 6072 22652 6100
rect 22327 6069 22339 6072
rect 22281 6063 22339 6069
rect 22646 6060 22652 6072
rect 22704 6060 22710 6112
rect 23566 6060 23572 6112
rect 23624 6100 23630 6112
rect 24213 6103 24271 6109
rect 24213 6100 24225 6103
rect 23624 6072 24225 6100
rect 23624 6060 23630 6072
rect 24213 6069 24225 6072
rect 24259 6069 24271 6103
rect 24213 6063 24271 6069
rect 24486 6060 24492 6112
rect 24544 6100 24550 6112
rect 24673 6103 24731 6109
rect 24673 6100 24685 6103
rect 24544 6072 24685 6100
rect 24544 6060 24550 6072
rect 24673 6069 24685 6072
rect 24719 6069 24731 6103
rect 24673 6063 24731 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 15286 5896 15292 5908
rect 15247 5868 15292 5896
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 16390 5896 16396 5908
rect 16303 5868 16396 5896
rect 16390 5856 16396 5868
rect 16448 5896 16454 5908
rect 17402 5896 17408 5908
rect 16448 5868 17408 5896
rect 16448 5856 16454 5868
rect 17402 5856 17408 5868
rect 17460 5896 17466 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 17460 5868 18429 5896
rect 17460 5856 17466 5868
rect 18417 5865 18429 5868
rect 18463 5896 18475 5899
rect 18598 5896 18604 5908
rect 18463 5868 18604 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 18966 5896 18972 5908
rect 18927 5868 18972 5896
rect 18966 5856 18972 5868
rect 19024 5856 19030 5908
rect 19058 5856 19064 5908
rect 19116 5896 19122 5908
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 19116 5868 19441 5896
rect 19116 5856 19122 5868
rect 19429 5865 19441 5868
rect 19475 5896 19487 5899
rect 20990 5896 20996 5908
rect 19475 5868 20996 5896
rect 19475 5865 19487 5868
rect 19429 5859 19487 5865
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 21358 5896 21364 5908
rect 21319 5868 21364 5896
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 22005 5899 22063 5905
rect 22005 5865 22017 5899
rect 22051 5896 22063 5899
rect 22094 5896 22100 5908
rect 22051 5868 22100 5896
rect 22051 5865 22063 5868
rect 22005 5859 22063 5865
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 25130 5896 25136 5908
rect 25091 5868 25136 5896
rect 25130 5856 25136 5868
rect 25188 5856 25194 5908
rect 12069 5831 12127 5837
rect 12069 5797 12081 5831
rect 12115 5828 12127 5831
rect 12894 5828 12900 5840
rect 12115 5800 12900 5828
rect 12115 5797 12127 5800
rect 12069 5791 12127 5797
rect 12894 5788 12900 5800
rect 12952 5788 12958 5840
rect 15654 5828 15660 5840
rect 15615 5800 15660 5828
rect 15654 5788 15660 5800
rect 15712 5788 15718 5840
rect 17304 5831 17362 5837
rect 17304 5797 17316 5831
rect 17350 5828 17362 5831
rect 17586 5828 17592 5840
rect 17350 5800 17592 5828
rect 17350 5797 17362 5800
rect 17304 5791 17362 5797
rect 17586 5788 17592 5800
rect 17644 5788 17650 5840
rect 21266 5828 21272 5840
rect 21227 5800 21272 5828
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 12250 5720 12256 5772
rect 12308 5760 12314 5772
rect 12428 5763 12486 5769
rect 12428 5760 12440 5763
rect 12308 5732 12440 5760
rect 12308 5720 12314 5732
rect 12428 5729 12440 5732
rect 12474 5760 12486 5763
rect 15749 5763 15807 5769
rect 12474 5732 15148 5760
rect 12474 5729 12486 5732
rect 12428 5723 12486 5729
rect 12158 5692 12164 5704
rect 12119 5664 12164 5692
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 15120 5633 15148 5732
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 16022 5760 16028 5772
rect 15795 5732 16028 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 16022 5720 16028 5732
rect 16080 5760 16086 5772
rect 16390 5760 16396 5772
rect 16080 5732 16396 5760
rect 16080 5720 16086 5732
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 17000 5732 17049 5760
rect 17000 5720 17006 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19576 5732 19717 5760
rect 19576 5720 19582 5732
rect 19705 5729 19717 5732
rect 19751 5760 19763 5763
rect 20254 5760 20260 5772
rect 19751 5732 20260 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 22002 5760 22008 5772
rect 21376 5732 22008 5760
rect 15930 5692 15936 5704
rect 15891 5664 15936 5692
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 21376 5692 21404 5732
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5760 22523 5763
rect 22554 5760 22560 5772
rect 22511 5732 22560 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 22554 5720 22560 5732
rect 22612 5760 22618 5772
rect 23014 5760 23020 5772
rect 22612 5732 23020 5760
rect 22612 5720 22618 5732
rect 23014 5720 23020 5732
rect 23072 5720 23078 5772
rect 23937 5763 23995 5769
rect 23937 5729 23949 5763
rect 23983 5760 23995 5763
rect 24854 5760 24860 5772
rect 23983 5732 24860 5760
rect 23983 5729 23995 5732
rect 23937 5723 23995 5729
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 19904 5664 21404 5692
rect 21453 5695 21511 5701
rect 15105 5627 15163 5633
rect 15105 5593 15117 5627
rect 15151 5624 15163 5627
rect 15948 5624 15976 5652
rect 19904 5633 19932 5664
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 15151 5596 15976 5624
rect 19889 5627 19947 5633
rect 15151 5593 15163 5596
rect 15105 5587 15163 5593
rect 19889 5593 19901 5627
rect 19935 5593 19947 5627
rect 19889 5587 19947 5593
rect 20806 5584 20812 5636
rect 20864 5624 20870 5636
rect 21468 5624 21496 5655
rect 23290 5652 23296 5704
rect 23348 5692 23354 5704
rect 24029 5695 24087 5701
rect 24029 5692 24041 5695
rect 23348 5664 24041 5692
rect 23348 5652 23354 5664
rect 24029 5661 24041 5664
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5692 24271 5695
rect 24670 5692 24676 5704
rect 24259 5664 24676 5692
rect 24259 5661 24271 5664
rect 24213 5655 24271 5661
rect 20864 5596 21496 5624
rect 22373 5627 22431 5633
rect 20864 5584 20870 5596
rect 22373 5593 22385 5627
rect 22419 5624 22431 5627
rect 22462 5624 22468 5636
rect 22419 5596 22468 5624
rect 22419 5593 22431 5596
rect 22373 5587 22431 5593
rect 22462 5584 22468 5596
rect 22520 5624 22526 5636
rect 23569 5627 23627 5633
rect 23569 5624 23581 5627
rect 22520 5596 23581 5624
rect 22520 5584 22526 5596
rect 23569 5593 23581 5596
rect 23615 5593 23627 5627
rect 24044 5624 24072 5655
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 24949 5627 25007 5633
rect 24949 5624 24961 5627
rect 24044 5596 24961 5624
rect 23569 5587 23627 5593
rect 24949 5593 24961 5596
rect 24995 5593 25007 5627
rect 24949 5587 25007 5593
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 13538 5556 13544 5568
rect 12584 5528 13544 5556
rect 12584 5516 12590 5528
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 16945 5559 17003 5565
rect 16945 5525 16957 5559
rect 16991 5556 17003 5559
rect 17310 5556 17316 5568
rect 16991 5528 17316 5556
rect 16991 5525 17003 5528
rect 16945 5519 17003 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 20346 5556 20352 5568
rect 20307 5528 20352 5556
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 20901 5559 20959 5565
rect 20901 5556 20913 5559
rect 20772 5528 20913 5556
rect 20772 5516 20778 5528
rect 20901 5525 20913 5528
rect 20947 5525 20959 5559
rect 20901 5519 20959 5525
rect 22649 5559 22707 5565
rect 22649 5525 22661 5559
rect 22695 5556 22707 5559
rect 22922 5556 22928 5568
rect 22695 5528 22928 5556
rect 22695 5525 22707 5528
rect 22649 5519 22707 5525
rect 22922 5516 22928 5528
rect 22980 5516 22986 5568
rect 23106 5556 23112 5568
rect 23067 5528 23112 5556
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 23474 5556 23480 5568
rect 23387 5528 23480 5556
rect 23474 5516 23480 5528
rect 23532 5556 23538 5568
rect 24670 5556 24676 5568
rect 23532 5528 24676 5556
rect 23532 5516 23538 5528
rect 24670 5516 24676 5528
rect 24728 5516 24734 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 15654 5312 15660 5364
rect 15712 5352 15718 5364
rect 15933 5355 15991 5361
rect 15933 5352 15945 5355
rect 15712 5324 15945 5352
rect 15712 5312 15718 5324
rect 15933 5321 15945 5324
rect 15979 5321 15991 5355
rect 19518 5352 19524 5364
rect 19479 5324 19524 5352
rect 15933 5315 15991 5321
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 19889 5355 19947 5361
rect 19889 5321 19901 5355
rect 19935 5352 19947 5355
rect 19978 5352 19984 5364
rect 19935 5324 19984 5352
rect 19935 5321 19947 5324
rect 19889 5315 19947 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20864 5324 21005 5352
rect 20864 5312 20870 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 20993 5315 21051 5321
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 21818 5312 21824 5364
rect 21876 5352 21882 5364
rect 22005 5355 22063 5361
rect 22005 5352 22017 5355
rect 21876 5324 22017 5352
rect 21876 5312 21882 5324
rect 22005 5321 22017 5324
rect 22051 5321 22063 5355
rect 23014 5352 23020 5364
rect 22975 5324 23020 5352
rect 22005 5315 22063 5321
rect 23014 5312 23020 5324
rect 23072 5312 23078 5364
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 23164 5324 24716 5352
rect 23164 5312 23170 5324
rect 11885 5287 11943 5293
rect 11885 5253 11897 5287
rect 11931 5284 11943 5287
rect 11931 5256 13032 5284
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 11330 5216 11336 5228
rect 11291 5188 11336 5216
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13004 5225 13032 5256
rect 22738 5244 22744 5296
rect 22796 5284 22802 5296
rect 23385 5287 23443 5293
rect 23385 5284 23397 5287
rect 22796 5256 23397 5284
rect 22796 5244 22802 5256
rect 23385 5253 23397 5256
rect 23431 5284 23443 5287
rect 24688 5284 24716 5324
rect 24854 5312 24860 5364
rect 24912 5352 24918 5364
rect 25685 5355 25743 5361
rect 25685 5352 25697 5355
rect 24912 5324 25697 5352
rect 24912 5312 24918 5324
rect 25685 5321 25697 5324
rect 25731 5321 25743 5355
rect 25685 5315 25743 5321
rect 25133 5287 25191 5293
rect 25133 5284 25145 5287
rect 23431 5256 23796 5284
rect 24688 5256 25145 5284
rect 23431 5253 23443 5256
rect 23385 5247 23443 5253
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13630 5216 13636 5228
rect 13035 5188 13636 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 18966 5216 18972 5228
rect 18927 5188 18972 5216
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 20346 5176 20352 5228
rect 20404 5216 20410 5228
rect 20530 5216 20536 5228
rect 20404 5188 20536 5216
rect 20404 5176 20410 5188
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 22462 5216 22468 5228
rect 22423 5188 22468 5216
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5216 22707 5219
rect 22833 5219 22891 5225
rect 22833 5216 22845 5219
rect 22695 5188 22845 5216
rect 22695 5185 22707 5188
rect 22649 5179 22707 5185
rect 22833 5185 22845 5188
rect 22879 5216 22891 5219
rect 23106 5216 23112 5228
rect 22879 5188 23112 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 23106 5176 23112 5188
rect 23164 5176 23170 5228
rect 23768 5225 23796 5256
rect 25133 5253 25145 5256
rect 25179 5253 25191 5287
rect 25133 5247 25191 5253
rect 23753 5219 23811 5225
rect 23753 5185 23765 5219
rect 23799 5185 23811 5219
rect 23753 5179 23811 5185
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 13170 5148 13176 5160
rect 12851 5120 13176 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5148 13967 5151
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13955 5120 14013 5148
rect 13955 5117 13967 5120
rect 13909 5111 13967 5117
rect 14001 5117 14013 5120
rect 14047 5148 14059 5151
rect 14090 5148 14096 5160
rect 14047 5120 14096 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 16758 5148 16764 5160
rect 16719 5120 16764 5148
rect 16758 5108 16764 5120
rect 16816 5148 16822 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 16816 5120 17325 5148
rect 16816 5108 16822 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5148 18383 5151
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 18371 5120 18797 5148
rect 18371 5117 18383 5120
rect 18325 5111 18383 5117
rect 18785 5117 18797 5120
rect 18831 5148 18843 5151
rect 19334 5148 19340 5160
rect 18831 5120 19340 5148
rect 18831 5117 18843 5120
rect 18785 5111 18843 5117
rect 19334 5108 19340 5120
rect 19392 5108 19398 5160
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20441 5151 20499 5157
rect 20441 5148 20453 5151
rect 20036 5120 20453 5148
rect 20036 5108 20042 5120
rect 20441 5117 20453 5120
rect 20487 5117 20499 5151
rect 22370 5148 22376 5160
rect 22283 5120 22376 5148
rect 20441 5111 20499 5117
rect 22370 5108 22376 5120
rect 22428 5148 22434 5160
rect 23566 5148 23572 5160
rect 22428 5120 23572 5148
rect 22428 5108 22434 5120
rect 23566 5108 23572 5120
rect 23624 5108 23630 5160
rect 13541 5083 13599 5089
rect 13541 5049 13553 5083
rect 13587 5080 13599 5083
rect 14246 5083 14304 5089
rect 14246 5080 14258 5083
rect 13587 5052 14258 5080
rect 13587 5049 13599 5052
rect 13541 5043 13599 5049
rect 14246 5049 14258 5052
rect 14292 5080 14304 5083
rect 15102 5080 15108 5092
rect 14292 5052 15108 5080
rect 14292 5049 14304 5052
rect 14246 5043 14304 5049
rect 15102 5040 15108 5052
rect 15160 5040 15166 5092
rect 18877 5083 18935 5089
rect 18877 5080 18889 5083
rect 17788 5052 18889 5080
rect 17788 5024 17816 5052
rect 18877 5049 18889 5052
rect 18923 5049 18935 5083
rect 18877 5043 18935 5049
rect 19518 5040 19524 5092
rect 19576 5080 19582 5092
rect 21913 5083 21971 5089
rect 19576 5052 20484 5080
rect 19576 5040 19582 5052
rect 12158 5012 12164 5024
rect 12119 4984 12164 5012
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 12400 4984 12449 5012
rect 12400 4972 12406 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 12437 4975 12495 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16942 5012 16948 5024
rect 16903 4984 16948 5012
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20456 5012 20484 5052
rect 21913 5049 21925 5083
rect 21959 5080 21971 5083
rect 22833 5083 22891 5089
rect 22833 5080 22845 5083
rect 21959 5052 22845 5080
rect 21959 5049 21971 5052
rect 21913 5043 21971 5049
rect 22833 5049 22845 5052
rect 22879 5049 22891 5083
rect 22833 5043 22891 5049
rect 24020 5083 24078 5089
rect 24020 5049 24032 5083
rect 24066 5080 24078 5083
rect 24670 5080 24676 5092
rect 24066 5052 24676 5080
rect 24066 5049 24078 5052
rect 24020 5043 24078 5049
rect 24670 5040 24676 5052
rect 24728 5040 24734 5092
rect 24762 5012 24768 5024
rect 20456 4984 24768 5012
rect 24762 4972 24768 4984
rect 24820 4972 24826 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 13170 4808 13176 4820
rect 11839 4780 13176 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 15930 4808 15936 4820
rect 15436 4780 15936 4808
rect 15436 4768 15442 4780
rect 15930 4768 15936 4780
rect 15988 4808 15994 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 15988 4780 16129 4808
rect 15988 4768 15994 4780
rect 16117 4777 16129 4780
rect 16163 4777 16175 4811
rect 16117 4771 16175 4777
rect 16482 4768 16488 4820
rect 16540 4808 16546 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16540 4780 16681 4808
rect 16540 4768 16546 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 16669 4771 16727 4777
rect 17037 4811 17095 4817
rect 17037 4777 17049 4811
rect 17083 4808 17095 4811
rect 17310 4808 17316 4820
rect 17083 4780 17316 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 17310 4768 17316 4780
rect 17368 4808 17374 4820
rect 17862 4808 17868 4820
rect 17368 4780 17868 4808
rect 17368 4768 17374 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18322 4808 18328 4820
rect 18187 4780 18328 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 18785 4811 18843 4817
rect 18785 4777 18797 4811
rect 18831 4808 18843 4811
rect 18966 4808 18972 4820
rect 18831 4780 18972 4808
rect 18831 4777 18843 4780
rect 18785 4771 18843 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19242 4808 19248 4820
rect 19203 4780 19248 4808
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 21266 4808 21272 4820
rect 20763 4780 21272 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 22925 4811 22983 4817
rect 22925 4777 22937 4811
rect 22971 4808 22983 4811
rect 23474 4808 23480 4820
rect 22971 4780 23480 4808
rect 22971 4777 22983 4780
rect 22925 4771 22983 4777
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 12161 4743 12219 4749
rect 12161 4709 12173 4743
rect 12207 4740 12219 4743
rect 12250 4740 12256 4752
rect 12207 4712 12256 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 16390 4700 16396 4752
rect 16448 4740 16454 4752
rect 17126 4740 17132 4752
rect 16448 4712 17132 4740
rect 16448 4700 16454 4712
rect 17126 4700 17132 4712
rect 17184 4700 17190 4752
rect 18233 4743 18291 4749
rect 18233 4709 18245 4743
rect 18279 4740 18291 4743
rect 20257 4743 20315 4749
rect 20257 4740 20269 4743
rect 18279 4712 20269 4740
rect 18279 4709 18291 4712
rect 18233 4703 18291 4709
rect 20257 4709 20269 4712
rect 20303 4740 20315 4743
rect 20346 4740 20352 4752
rect 20303 4712 20352 4740
rect 20303 4709 20315 4712
rect 20257 4703 20315 4709
rect 20346 4700 20352 4712
rect 20404 4700 20410 4752
rect 20530 4700 20536 4752
rect 20588 4740 20594 4752
rect 20990 4740 20996 4752
rect 20588 4712 20996 4740
rect 20588 4700 20594 4712
rect 20990 4700 20996 4712
rect 21048 4740 21054 4752
rect 21146 4743 21204 4749
rect 21146 4740 21158 4743
rect 21048 4712 21158 4740
rect 21048 4700 21054 4712
rect 21146 4709 21158 4712
rect 21192 4709 21204 4743
rect 21146 4703 21204 4709
rect 12526 4681 12532 4684
rect 12520 4672 12532 4681
rect 12487 4644 12532 4672
rect 12520 4635 12532 4644
rect 12526 4632 12532 4635
rect 12584 4632 12590 4684
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 15028 4644 15577 4672
rect 12250 4604 12256 4616
rect 12211 4576 12256 4604
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 13446 4468 13452 4480
rect 13228 4440 13452 4468
rect 13228 4428 13234 4440
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 15028 4477 15056 4644
rect 15565 4641 15577 4644
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 16577 4675 16635 4681
rect 16577 4641 16589 4675
rect 16623 4672 16635 4675
rect 17586 4672 17592 4684
rect 16623 4644 17592 4672
rect 16623 4641 16635 4644
rect 16577 4635 16635 4641
rect 17586 4632 17592 4644
rect 17644 4632 17650 4684
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 19978 4672 19984 4684
rect 19659 4644 19984 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 23641 4675 23699 4681
rect 23641 4672 23653 4675
rect 23216 4644 23653 4672
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4604 17371 4607
rect 17402 4604 17408 4616
rect 17359 4576 17408 4604
rect 17359 4573 17371 4576
rect 17313 4567 17371 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19886 4604 19892 4616
rect 19847 4576 19892 4604
rect 19705 4567 19763 4573
rect 19153 4539 19211 4545
rect 19153 4505 19165 4539
rect 19199 4536 19211 4539
rect 19720 4536 19748 4567
rect 19886 4564 19892 4576
rect 19944 4564 19950 4616
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20864 4576 20913 4604
rect 20864 4564 20870 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 20438 4536 20444 4548
rect 19199 4508 20444 4536
rect 19199 4505 19211 4508
rect 19153 4499 19211 4505
rect 20438 4496 20444 4508
rect 20496 4496 20502 4548
rect 23216 4545 23244 4644
rect 23641 4641 23653 4644
rect 23687 4641 23699 4675
rect 23641 4635 23699 4641
rect 23385 4607 23443 4613
rect 23385 4573 23397 4607
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 23201 4539 23259 4545
rect 23201 4536 23213 4539
rect 22296 4508 23213 4536
rect 22296 4480 22324 4508
rect 23201 4505 23213 4508
rect 23247 4505 23259 4539
rect 23201 4499 23259 4505
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14884 4440 15025 4468
rect 14884 4428 14890 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 15749 4471 15807 4477
rect 15749 4437 15761 4471
rect 15795 4468 15807 4471
rect 17126 4468 17132 4480
rect 15795 4440 17132 4468
rect 15795 4437 15807 4440
rect 15749 4431 15807 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 17586 4428 17592 4480
rect 17644 4468 17650 4480
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17644 4440 17693 4468
rect 17644 4428 17650 4440
rect 17681 4437 17693 4440
rect 17727 4437 17739 4471
rect 22278 4468 22284 4480
rect 22239 4440 22284 4468
rect 17681 4431 17739 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22738 4428 22744 4480
rect 22796 4468 22802 4480
rect 23400 4468 23428 4567
rect 24762 4468 24768 4480
rect 22796 4440 23428 4468
rect 24723 4440 24768 4468
rect 22796 4428 22802 4440
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12526 4264 12532 4276
rect 12299 4236 12532 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 17221 4267 17279 4273
rect 17221 4233 17233 4267
rect 17267 4264 17279 4267
rect 17402 4264 17408 4276
rect 17267 4236 17408 4264
rect 17267 4233 17279 4236
rect 17221 4227 17279 4233
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 19886 4264 19892 4276
rect 19628 4236 19892 4264
rect 14734 4156 14740 4208
rect 14792 4196 14798 4208
rect 19628 4196 19656 4236
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 20990 4264 20996 4276
rect 20951 4236 20996 4264
rect 20990 4224 20996 4236
rect 21048 4264 21054 4276
rect 21450 4264 21456 4276
rect 21048 4236 21456 4264
rect 21048 4224 21054 4236
rect 21450 4224 21456 4236
rect 21508 4264 21514 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21508 4236 21925 4264
rect 21508 4224 21514 4236
rect 21913 4233 21925 4236
rect 21959 4233 21971 4267
rect 21913 4227 21971 4233
rect 22738 4224 22744 4276
rect 22796 4264 22802 4276
rect 23017 4267 23075 4273
rect 23017 4264 23029 4267
rect 22796 4236 23029 4264
rect 22796 4224 22802 4236
rect 23017 4233 23029 4236
rect 23063 4264 23075 4267
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 23063 4236 23397 4264
rect 23063 4233 23075 4236
rect 23017 4227 23075 4233
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 23385 4227 23443 4233
rect 14792 4168 15148 4196
rect 14792 4156 14798 4168
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 8202 4128 8208 4140
rect 7800 4100 8208 4128
rect 7800 4088 7806 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12986 4128 12992 4140
rect 12584 4100 12992 4128
rect 12584 4088 12590 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 15120 4128 15148 4168
rect 19352 4168 19656 4196
rect 16577 4131 16635 4137
rect 16577 4128 16589 4131
rect 15120 4100 16589 4128
rect 16577 4097 16589 4100
rect 16623 4097 16635 4131
rect 16577 4091 16635 4097
rect 16761 4131 16819 4137
rect 16761 4097 16773 4131
rect 16807 4128 16819 4131
rect 16942 4128 16948 4140
rect 16807 4100 16948 4128
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11379 4032 11897 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11885 4029 11897 4032
rect 11931 4060 11943 4063
rect 12342 4060 12348 4072
rect 11931 4032 12348 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 13446 4060 13452 4072
rect 13403 4032 13452 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13630 4069 13636 4072
rect 13624 4060 13636 4069
rect 13591 4032 13636 4060
rect 13624 4023 13636 4032
rect 13630 4020 13636 4023
rect 13688 4020 13694 4072
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 16390 4060 16396 4072
rect 15703 4032 16396 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16592 4060 16620 4091
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 17828 4100 18092 4128
rect 17828 4088 17834 4100
rect 18064 4060 18092 4100
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 18380 4100 18521 4128
rect 18380 4088 18386 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 18874 4128 18880 4140
rect 18739 4100 18880 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19352 4128 19380 4168
rect 19199 4100 19380 4128
rect 23400 4128 23428 4227
rect 24670 4224 24676 4276
rect 24728 4264 24734 4276
rect 25041 4267 25099 4273
rect 25041 4264 25053 4267
rect 24728 4236 25053 4264
rect 24728 4224 24734 4236
rect 25041 4233 25053 4236
rect 25087 4233 25099 4267
rect 25041 4227 25099 4233
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23400 4100 23673 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 16592 4032 18000 4060
rect 18064 4032 18429 4060
rect 16485 3995 16543 4001
rect 16485 3992 16497 3995
rect 15948 3964 16497 3992
rect 15948 3936 15976 3964
rect 16485 3961 16497 3964
rect 16531 3961 16543 3995
rect 16485 3955 16543 3961
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12713 3927 12771 3933
rect 12713 3924 12725 3927
rect 12308 3896 12725 3924
rect 12308 3884 12314 3896
rect 12713 3893 12725 3896
rect 12759 3924 12771 3927
rect 13265 3927 13323 3933
rect 13265 3924 13277 3927
rect 12759 3896 13277 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 13265 3893 13277 3896
rect 13311 3924 13323 3927
rect 13446 3924 13452 3936
rect 13311 3896 13452 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13446 3884 13452 3896
rect 13504 3924 13510 3936
rect 14090 3924 14096 3936
rect 13504 3896 14096 3924
rect 13504 3884 13510 3896
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 14826 3924 14832 3936
rect 14783 3896 14832 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15930 3924 15936 3936
rect 15891 3896 15936 3924
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 17972 3924 18000 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 19337 4063 19395 4069
rect 19337 4029 19349 4063
rect 19383 4060 19395 4063
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 19383 4032 19625 4060
rect 19383 4029 19395 4032
rect 19337 4023 19395 4029
rect 19613 4029 19625 4032
rect 19659 4060 19671 4063
rect 20806 4060 20812 4072
rect 19659 4032 20812 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 20806 4020 20812 4032
rect 20864 4060 20870 4072
rect 21545 4063 21603 4069
rect 21545 4060 21557 4063
rect 20864 4032 21557 4060
rect 20864 4020 20870 4032
rect 21545 4029 21557 4032
rect 21591 4029 21603 4063
rect 21545 4023 21603 4029
rect 18966 3952 18972 4004
rect 19024 3992 19030 4004
rect 19858 3995 19916 4001
rect 19858 3992 19870 3995
rect 19024 3964 19870 3992
rect 19024 3952 19030 3964
rect 19858 3961 19870 3964
rect 19904 3992 19916 3995
rect 20070 3992 20076 4004
rect 19904 3964 20076 3992
rect 19904 3961 19916 3964
rect 19858 3955 19916 3961
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 21560 3992 21588 4023
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 22649 4063 22707 4069
rect 22649 4060 22661 4063
rect 22152 4032 22661 4060
rect 22152 4020 22158 4032
rect 22649 4029 22661 4032
rect 22695 4029 22707 4063
rect 22649 4023 22707 4029
rect 22738 3992 22744 4004
rect 21560 3964 22744 3992
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 23842 3952 23848 4004
rect 23900 4001 23906 4004
rect 23900 3995 23964 4001
rect 23900 3961 23918 3995
rect 23952 3961 23964 3995
rect 23900 3955 23964 3961
rect 23900 3952 23906 3955
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17972 3896 18061 3924
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 19337 3927 19395 3933
rect 19337 3924 19349 3927
rect 18380 3896 19349 3924
rect 18380 3884 18386 3896
rect 19337 3893 19349 3896
rect 19383 3924 19395 3927
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 19383 3896 19441 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 22278 3924 22284 3936
rect 22239 3896 22284 3924
rect 19429 3887 19487 3893
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 11698 3720 11704 3732
rect 11659 3692 11704 3720
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 13449 3723 13507 3729
rect 13449 3689 13461 3723
rect 13495 3720 13507 3723
rect 13630 3720 13636 3732
rect 13495 3692 13636 3720
rect 13495 3689 13507 3692
rect 13449 3683 13507 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14550 3720 14556 3732
rect 14240 3692 14556 3720
rect 14240 3680 14246 3692
rect 14550 3680 14556 3692
rect 14608 3720 14614 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14608 3692 14657 3720
rect 14608 3680 14614 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 15102 3720 15108 3732
rect 14884 3692 15108 3720
rect 14884 3680 14890 3692
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 19337 3723 19395 3729
rect 19337 3689 19349 3723
rect 19383 3720 19395 3723
rect 19426 3720 19432 3732
rect 19383 3692 19432 3720
rect 19383 3689 19395 3692
rect 19337 3683 19395 3689
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 19978 3680 19984 3732
rect 20036 3720 20042 3732
rect 20349 3723 20407 3729
rect 20349 3720 20361 3723
rect 20036 3692 20361 3720
rect 20036 3680 20042 3692
rect 20349 3689 20361 3692
rect 20395 3689 20407 3723
rect 20349 3683 20407 3689
rect 20438 3680 20444 3732
rect 20496 3720 20502 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20496 3692 20913 3720
rect 20496 3680 20502 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 21358 3720 21364 3732
rect 21319 3692 21364 3720
rect 20901 3683 20959 3689
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22370 3720 22376 3732
rect 22143 3692 22376 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 22554 3720 22560 3732
rect 22515 3692 22560 3720
rect 22554 3680 22560 3692
rect 22612 3680 22618 3732
rect 23290 3720 23296 3732
rect 23251 3692 23296 3720
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 23750 3720 23756 3732
rect 23711 3692 23756 3720
rect 23750 3680 23756 3692
rect 23808 3680 23814 3732
rect 24854 3720 24860 3732
rect 24815 3692 24860 3720
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 25222 3720 25228 3732
rect 25183 3692 25228 3720
rect 25222 3680 25228 3692
rect 25280 3680 25286 3732
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 25372 3692 25417 3720
rect 25372 3680 25378 3692
rect 14001 3655 14059 3661
rect 14001 3621 14013 3655
rect 14047 3652 14059 3655
rect 14090 3652 14096 3664
rect 14047 3624 14096 3652
rect 14047 3621 14059 3624
rect 14001 3615 14059 3621
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 16209 3655 16267 3661
rect 16209 3621 16221 3655
rect 16255 3652 16267 3655
rect 16752 3655 16810 3661
rect 16752 3652 16764 3655
rect 16255 3624 16764 3652
rect 16255 3621 16267 3624
rect 16209 3615 16267 3621
rect 16752 3621 16764 3624
rect 16798 3652 16810 3655
rect 16942 3652 16948 3664
rect 16798 3624 16948 3652
rect 16798 3621 16810 3624
rect 16752 3615 16810 3621
rect 16942 3612 16948 3624
rect 17000 3612 17006 3664
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3584 10563 3587
rect 10778 3584 10784 3596
rect 10551 3556 10784 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3584 11575 3587
rect 12250 3584 12256 3596
rect 11563 3556 12256 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3584 12587 3587
rect 12710 3584 12716 3596
rect 12575 3556 12716 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 15378 3584 15384 3596
rect 15339 3556 15384 3584
rect 15378 3544 15384 3556
rect 15436 3584 15442 3596
rect 15654 3584 15660 3596
rect 15436 3556 15660 3584
rect 15436 3544 15442 3556
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 19444 3584 19472 3680
rect 20070 3652 20076 3664
rect 20031 3624 20076 3652
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 23198 3612 23204 3664
rect 23256 3652 23262 3664
rect 23661 3655 23719 3661
rect 23661 3652 23673 3655
rect 23256 3624 23673 3652
rect 23256 3612 23262 3624
rect 23661 3621 23673 3624
rect 23707 3621 23719 3655
rect 23661 3615 23719 3621
rect 19978 3584 19984 3596
rect 19444 3556 19984 3584
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13906 3516 13912 3528
rect 13136 3488 13912 3516
rect 13136 3476 13142 3488
rect 13906 3476 13912 3488
rect 13964 3516 13970 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13964 3488 14105 3516
rect 13964 3476 13970 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14826 3516 14832 3528
rect 14323 3488 14832 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 16390 3476 16396 3528
rect 16448 3516 16454 3528
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 16448 3488 16497 3516
rect 16448 3476 16454 3488
rect 16485 3485 16497 3488
rect 16531 3485 16543 3519
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 16485 3479 16543 3485
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 18874 3448 18880 3460
rect 18196 3420 18880 3448
rect 18196 3408 18202 3420
rect 18874 3408 18880 3420
rect 18932 3448 18938 3460
rect 19536 3448 19564 3479
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 23937 3519 23995 3525
rect 21508 3488 21553 3516
rect 21508 3476 21514 3488
rect 23937 3485 23949 3519
rect 23983 3485 23995 3519
rect 25498 3516 25504 3528
rect 25459 3488 25504 3516
rect 23937 3479 23995 3485
rect 18932 3420 19564 3448
rect 18932 3408 18938 3420
rect 23842 3408 23848 3460
rect 23900 3448 23906 3460
rect 23952 3448 23980 3479
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 24397 3451 24455 3457
rect 24397 3448 24409 3451
rect 23900 3420 24409 3448
rect 23900 3408 23906 3420
rect 24397 3417 24409 3420
rect 24443 3448 24455 3451
rect 24762 3448 24768 3460
rect 24443 3420 24768 3448
rect 24443 3417 24455 3420
rect 24397 3411 24455 3417
rect 24762 3408 24768 3420
rect 24820 3448 24826 3460
rect 25516 3448 25544 3476
rect 24820 3420 25544 3448
rect 24820 3408 24826 3420
rect 10686 3380 10692 3392
rect 10647 3352 10692 3380
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 12713 3383 12771 3389
rect 12713 3349 12725 3383
rect 12759 3380 12771 3383
rect 13538 3380 13544 3392
rect 12759 3352 13544 3380
rect 12759 3349 12771 3352
rect 12713 3343 12771 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13722 3380 13728 3392
rect 13679 3352 13728 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 15562 3380 15568 3392
rect 15523 3352 15568 3380
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 16724 3352 17877 3380
rect 16724 3340 16730 3352
rect 17865 3349 17877 3352
rect 17911 3380 17923 3383
rect 18414 3380 18420 3392
rect 17911 3352 18420 3380
rect 17911 3349 17923 3352
rect 17865 3343 17923 3349
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 18966 3380 18972 3392
rect 18927 3352 18972 3380
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12250 3176 12256 3188
rect 12211 3148 12256 3176
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12768 3148 12909 3176
rect 12768 3136 12774 3148
rect 12897 3145 12909 3148
rect 12943 3145 12955 3179
rect 13354 3176 13360 3188
rect 13315 3148 13360 3176
rect 12897 3139 12955 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13906 3136 13912 3188
rect 13964 3176 13970 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 13964 3148 14381 3176
rect 13964 3136 13970 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 15933 3179 15991 3185
rect 14369 3139 14427 3145
rect 14568 3148 15700 3176
rect 10413 3111 10471 3117
rect 10413 3077 10425 3111
rect 10459 3108 10471 3111
rect 14090 3108 14096 3120
rect 10459 3080 11284 3108
rect 14003 3080 14096 3108
rect 10459 3077 10471 3080
rect 10413 3071 10471 3077
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 11146 2972 11152 2984
rect 10275 2944 11152 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11256 2981 11284 3080
rect 14090 3068 14096 3080
rect 14148 3108 14154 3120
rect 14568 3108 14596 3148
rect 14148 3080 14596 3108
rect 15672 3108 15700 3148
rect 15933 3145 15945 3179
rect 15979 3176 15991 3179
rect 16942 3176 16948 3188
rect 15979 3148 16948 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17310 3176 17316 3188
rect 17271 3148 17316 3176
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 19705 3179 19763 3185
rect 19705 3145 19717 3179
rect 19751 3176 19763 3179
rect 20070 3176 20076 3188
rect 19751 3148 20076 3176
rect 19751 3145 19763 3148
rect 19705 3139 19763 3145
rect 20070 3136 20076 3148
rect 20128 3176 20134 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 20128 3148 20269 3176
rect 20128 3136 20134 3148
rect 20257 3145 20269 3148
rect 20303 3145 20315 3179
rect 20257 3139 20315 3145
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3176 20867 3179
rect 21266 3176 21272 3188
rect 20855 3148 21272 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 16758 3108 16764 3120
rect 15672 3080 16764 3108
rect 14148 3068 14154 3080
rect 16758 3068 16764 3080
rect 16816 3068 16822 3120
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 14550 3040 14556 3052
rect 12492 3012 12537 3040
rect 14511 3012 14556 3040
rect 12492 3000 12498 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 20272 3040 20300 3139
rect 21266 3136 21272 3148
rect 21324 3176 21330 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 21324 3148 22201 3176
rect 21324 3136 21330 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 22189 3139 22247 3145
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 23256 3148 23305 3176
rect 23256 3136 23262 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23293 3139 23351 3145
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3108 20775 3111
rect 21082 3108 21088 3120
rect 20763 3080 21088 3108
rect 20763 3077 20775 3080
rect 20717 3071 20775 3077
rect 21082 3068 21088 3080
rect 21140 3068 21146 3120
rect 21450 3068 21456 3120
rect 21508 3108 21514 3120
rect 21821 3111 21879 3117
rect 21821 3108 21833 3111
rect 21508 3080 21833 3108
rect 21508 3068 21514 3080
rect 21821 3077 21833 3080
rect 21867 3077 21879 3111
rect 23308 3108 23336 3139
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 23845 3179 23903 3185
rect 23845 3176 23857 3179
rect 23808 3148 23857 3176
rect 23808 3136 23814 3148
rect 23845 3145 23857 3148
rect 23891 3145 23903 3179
rect 23845 3139 23903 3145
rect 25225 3179 25283 3185
rect 25225 3145 25237 3179
rect 25271 3176 25283 3179
rect 25314 3176 25320 3188
rect 25271 3148 25320 3176
rect 25271 3145 25283 3148
rect 25225 3139 25283 3145
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 25498 3136 25504 3188
rect 25556 3176 25562 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25556 3148 25881 3176
rect 25556 3136 25562 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 25869 3139 25927 3145
rect 24397 3111 24455 3117
rect 24397 3108 24409 3111
rect 23308 3080 24409 3108
rect 21821 3071 21879 3077
rect 24397 3077 24409 3080
rect 24443 3077 24455 3111
rect 24397 3071 24455 3077
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 20272 3012 21373 3040
rect 21361 3009 21373 3012
rect 21407 3009 21419 3043
rect 21361 3003 21419 3009
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11287 2944 11805 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 13354 2932 13360 2984
rect 13412 2972 13418 2984
rect 13449 2975 13507 2981
rect 13449 2972 13461 2975
rect 13412 2944 13461 2972
rect 13412 2932 13418 2944
rect 13449 2941 13461 2944
rect 13495 2941 13507 2975
rect 13449 2935 13507 2941
rect 14568 2904 14596 3000
rect 14826 2981 14832 2984
rect 14820 2972 14832 2981
rect 14787 2944 14832 2972
rect 14820 2935 14832 2944
rect 14826 2932 14832 2935
rect 14884 2932 14890 2984
rect 18322 2972 18328 2984
rect 17788 2944 18328 2972
rect 16390 2904 16396 2916
rect 14568 2876 16396 2904
rect 16390 2864 16396 2876
rect 16448 2904 16454 2916
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 16448 2876 16497 2904
rect 16448 2864 16454 2876
rect 16485 2873 16497 2876
rect 16531 2904 16543 2907
rect 17586 2904 17592 2916
rect 16531 2876 17592 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 17586 2864 17592 2876
rect 17644 2904 17650 2916
rect 17788 2913 17816 2944
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 18581 2975 18639 2981
rect 18581 2972 18593 2975
rect 18472 2944 18593 2972
rect 18472 2932 18478 2944
rect 18581 2941 18593 2944
rect 18627 2941 18639 2975
rect 21174 2972 21180 2984
rect 21135 2944 21180 2972
rect 18581 2935 18639 2941
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 22554 2972 22560 2984
rect 22511 2944 22560 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24412 2972 24440 3071
rect 25222 3000 25228 3052
rect 25280 3040 25286 3052
rect 25501 3043 25559 3049
rect 25501 3040 25513 3043
rect 25280 3012 25513 3040
rect 25280 3000 25286 3012
rect 25501 3009 25513 3012
rect 25547 3009 25559 3043
rect 25501 3003 25559 3009
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 24412 2944 24593 2972
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 17773 2907 17831 2913
rect 17773 2904 17785 2907
rect 17644 2876 17785 2904
rect 17644 2864 17650 2876
rect 17773 2873 17785 2876
rect 17819 2873 17831 2907
rect 17773 2867 17831 2873
rect 21082 2864 21088 2916
rect 21140 2904 21146 2916
rect 21266 2904 21272 2916
rect 21140 2876 21272 2904
rect 21140 2864 21146 2876
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 13630 2836 13636 2848
rect 13591 2808 13636 2836
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 14366 2796 14372 2848
rect 14424 2836 14430 2848
rect 15470 2836 15476 2848
rect 14424 2808 15476 2836
rect 14424 2796 14430 2808
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 16942 2836 16948 2848
rect 16903 2808 16948 2836
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 22649 2839 22707 2845
rect 22649 2805 22661 2839
rect 22695 2836 22707 2839
rect 23198 2836 23204 2848
rect 22695 2808 23204 2836
rect 22695 2805 22707 2808
rect 22649 2799 22707 2805
rect 23198 2796 23204 2808
rect 23256 2796 23262 2848
rect 24762 2836 24768 2848
rect 24723 2808 24768 2836
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 5994 2632 6000 2644
rect 5767 2604 6000 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 8297 2635 8355 2641
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 8386 2632 8392 2644
rect 8343 2604 8392 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 13814 2632 13820 2644
rect 13775 2604 13820 2632
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 14826 2632 14832 2644
rect 14231 2604 14832 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 17000 2604 17693 2632
rect 17000 2592 17006 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 17681 2595 17739 2601
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 12492 2536 12537 2564
rect 12492 2524 12498 2536
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 2958 2496 2964 2508
rect 2823 2468 2964 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 2958 2456 2964 2468
rect 3016 2496 3022 2508
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 3016 2468 3341 2496
rect 3016 2456 3022 2468
rect 3329 2465 3341 2468
rect 3375 2465 3387 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 3329 2459 3387 2465
rect 5534 2456 5540 2468
rect 5592 2496 5598 2508
rect 6089 2499 6147 2505
rect 6089 2496 6101 2499
rect 5592 2468 6101 2496
rect 5592 2456 5598 2468
rect 6089 2465 6101 2468
rect 6135 2465 6147 2499
rect 6089 2459 6147 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8386 2496 8392 2508
rect 8159 2468 8392 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10686 2496 10692 2508
rect 10367 2468 10692 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 10686 2456 10692 2468
rect 10744 2496 10750 2508
rect 10873 2499 10931 2505
rect 10873 2496 10885 2499
rect 10744 2468 10885 2496
rect 10744 2456 10750 2468
rect 10873 2465 10885 2468
rect 10919 2465 10931 2499
rect 10873 2459 10931 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11514 2496 11520 2508
rect 11471 2468 11520 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11514 2456 11520 2468
rect 11572 2496 11578 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11572 2468 11989 2496
rect 11572 2456 11578 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13832 2496 13860 2592
rect 17696 2564 17724 2595
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19797 2635 19855 2641
rect 19797 2601 19809 2635
rect 19843 2632 19855 2635
rect 19978 2632 19984 2644
rect 19843 2604 19984 2632
rect 19843 2601 19855 2604
rect 19797 2595 19855 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20901 2635 20959 2641
rect 20901 2601 20913 2635
rect 20947 2632 20959 2635
rect 21174 2632 21180 2644
rect 20947 2604 21180 2632
rect 20947 2601 20959 2604
rect 20901 2595 20959 2601
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 21358 2632 21364 2644
rect 21319 2604 21364 2632
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 23842 2632 23848 2644
rect 23803 2604 23848 2632
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 17696 2536 18920 2564
rect 13219 2468 13860 2496
rect 14277 2499 14335 2505
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14366 2496 14372 2508
rect 14323 2468 14372 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14366 2456 14372 2468
rect 14424 2496 14430 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14424 2468 14841 2496
rect 14424 2456 14430 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 16114 2496 16120 2508
rect 15988 2468 16120 2496
rect 15988 2456 15994 2468
rect 16114 2456 16120 2468
rect 16172 2496 16178 2508
rect 16301 2499 16359 2505
rect 16301 2496 16313 2499
rect 16172 2468 16313 2496
rect 16172 2456 16178 2468
rect 16301 2465 16313 2468
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 18693 2499 18751 2505
rect 18693 2496 18705 2499
rect 17083 2468 18705 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 16390 2428 16396 2440
rect 13127 2400 16396 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 16482 2388 16488 2440
rect 16540 2428 16546 2440
rect 16540 2400 16633 2428
rect 16540 2388 16546 2400
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 4062 2360 4068 2372
rect 3007 2332 4068 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 15378 2320 15384 2372
rect 15436 2360 15442 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 15436 2332 15945 2360
rect 15436 2320 15442 2332
rect 15933 2329 15945 2332
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 10502 2292 10508 2304
rect 10463 2264 10508 2292
rect 8665 2255 8723 2261
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2292 15347 2295
rect 16500 2292 16528 2388
rect 18322 2360 18328 2372
rect 18283 2332 18328 2360
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 18616 2360 18644 2468
rect 18693 2465 18705 2468
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 18782 2428 18788 2440
rect 18743 2400 18788 2428
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 18892 2437 18920 2536
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 20162 2496 20168 2508
rect 19935 2468 20168 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20162 2456 20168 2468
rect 20220 2496 20226 2508
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 20220 2468 20453 2496
rect 20220 2456 20226 2468
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 21726 2496 21732 2508
rect 21687 2468 21732 2496
rect 20441 2459 20499 2465
rect 21726 2456 21732 2468
rect 21784 2496 21790 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 21784 2468 22293 2496
rect 21784 2456 21790 2468
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22830 2496 22836 2508
rect 22791 2468 22836 2496
rect 22281 2459 22339 2465
rect 22830 2456 22836 2468
rect 22888 2496 22894 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22888 2468 23397 2496
rect 22888 2456 22894 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 23385 2459 23443 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23992 2468 24593 2496
rect 23992 2456 23998 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 18966 2360 18972 2372
rect 18616 2332 18972 2360
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 23017 2363 23075 2369
rect 23017 2329 23029 2363
rect 23063 2360 23075 2363
rect 24670 2360 24676 2372
rect 23063 2332 24676 2360
rect 23063 2329 23075 2332
rect 23017 2323 23075 2329
rect 24670 2320 24676 2332
rect 24728 2320 24734 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 26142 2360 26148 2372
rect 24811 2332 26148 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 26142 2320 26148 2332
rect 26200 2320 26206 2372
rect 15335 2264 16528 2292
rect 15335 2261 15347 2264
rect 15289 2255 15347 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17313 2295 17371 2301
rect 17313 2292 17325 2295
rect 17276 2264 17325 2292
rect 17276 2252 17282 2264
rect 17313 2261 17325 2264
rect 17359 2292 17371 2295
rect 18782 2292 18788 2304
rect 17359 2264 18788 2292
rect 17359 2261 17371 2264
rect 17313 2255 17371 2261
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 19334 2292 19340 2304
rect 19295 2264 19340 2292
rect 19334 2252 19340 2264
rect 19392 2252 19398 2304
rect 20070 2292 20076 2304
rect 20031 2264 20076 2292
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 21910 2292 21916 2304
rect 21871 2264 21916 2292
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 13906 552 13912 604
rect 13964 592 13970 604
rect 14366 592 14372 604
rect 13964 564 14372 592
rect 13964 552 13970 564
rect 14366 552 14372 564
rect 14424 552 14430 604
rect 17126 552 17132 604
rect 17184 592 17190 604
rect 17310 592 17316 604
rect 17184 564 17316 592
rect 17184 552 17190 564
rect 17310 552 17316 564
rect 17368 552 17374 604
rect 22922 552 22928 604
rect 22980 592 22986 604
rect 23474 592 23480 604
rect 22980 564 23480 592
rect 22980 552 22986 564
rect 23474 552 23480 564
rect 23532 552 23538 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 15936 25440 15988 25492
rect 17960 25440 18012 25492
rect 20076 25440 20128 25492
rect 22744 25440 22796 25492
rect 14372 25304 14424 25356
rect 16948 25304 17000 25356
rect 19432 25347 19484 25356
rect 19432 25313 19441 25347
rect 19441 25313 19475 25347
rect 19475 25313 19484 25347
rect 19432 25304 19484 25313
rect 22008 25347 22060 25356
rect 22008 25313 22017 25347
rect 22017 25313 22051 25347
rect 22051 25313 22060 25347
rect 22008 25304 22060 25313
rect 17592 25236 17644 25288
rect 17316 25168 17368 25220
rect 16396 25100 16448 25152
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 21640 25100 21692 25152
rect 24676 25100 24728 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 18972 24896 19024 24948
rect 23572 24896 23624 24948
rect 16396 24828 16448 24880
rect 21732 24828 21784 24880
rect 22008 24871 22060 24880
rect 22008 24837 22017 24871
rect 22017 24837 22051 24871
rect 22051 24837 22060 24871
rect 22008 24828 22060 24837
rect 19524 24760 19576 24812
rect 12900 24692 12952 24744
rect 14280 24735 14332 24744
rect 14280 24701 14289 24735
rect 14289 24701 14323 24735
rect 14323 24701 14332 24735
rect 14280 24692 14332 24701
rect 18144 24692 18196 24744
rect 21548 24692 21600 24744
rect 14372 24624 14424 24676
rect 15200 24667 15252 24676
rect 15200 24633 15209 24667
rect 15209 24633 15243 24667
rect 15243 24633 15252 24667
rect 15200 24624 15252 24633
rect 17500 24624 17552 24676
rect 19432 24624 19484 24676
rect 20168 24624 20220 24676
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 14464 24599 14516 24608
rect 14464 24565 14473 24599
rect 14473 24565 14507 24599
rect 14507 24565 14516 24599
rect 14464 24556 14516 24565
rect 15384 24599 15436 24608
rect 15384 24565 15393 24599
rect 15393 24565 15427 24599
rect 15427 24565 15436 24599
rect 15384 24556 15436 24565
rect 15752 24599 15804 24608
rect 15752 24565 15761 24599
rect 15761 24565 15795 24599
rect 15795 24565 15804 24599
rect 15752 24556 15804 24565
rect 16948 24556 17000 24608
rect 18144 24556 18196 24608
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 22100 24624 22152 24676
rect 21824 24556 21876 24608
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 23664 24599 23716 24608
rect 23664 24565 23673 24599
rect 23673 24565 23707 24599
rect 23707 24565 23716 24599
rect 23664 24556 23716 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 15384 24352 15436 24404
rect 16304 24395 16356 24404
rect 16304 24361 16313 24395
rect 16313 24361 16347 24395
rect 16347 24361 16356 24395
rect 16304 24352 16356 24361
rect 20628 24352 20680 24404
rect 21456 24395 21508 24404
rect 21456 24361 21465 24395
rect 21465 24361 21499 24395
rect 21499 24361 21508 24395
rect 21456 24352 21508 24361
rect 21916 24395 21968 24404
rect 21916 24361 21925 24395
rect 21925 24361 21959 24395
rect 21959 24361 21968 24395
rect 21916 24352 21968 24361
rect 22560 24395 22612 24404
rect 22560 24361 22569 24395
rect 22569 24361 22603 24395
rect 22603 24361 22612 24395
rect 22560 24352 22612 24361
rect 23756 24352 23808 24404
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 10140 24284 10192 24336
rect 15568 24284 15620 24336
rect 15752 24284 15804 24336
rect 12072 24216 12124 24268
rect 13728 24259 13780 24268
rect 13728 24225 13737 24259
rect 13737 24225 13771 24259
rect 13771 24225 13780 24259
rect 13728 24216 13780 24225
rect 16672 24216 16724 24268
rect 18052 24216 18104 24268
rect 18328 24216 18380 24268
rect 21088 24216 21140 24268
rect 22376 24259 22428 24268
rect 22376 24225 22385 24259
rect 22385 24225 22419 24259
rect 22419 24225 22428 24259
rect 22376 24216 22428 24225
rect 23112 24216 23164 24268
rect 24216 24216 24268 24268
rect 11796 24148 11848 24200
rect 12716 24148 12768 24200
rect 13636 24148 13688 24200
rect 14004 24191 14056 24200
rect 14004 24157 14013 24191
rect 14013 24157 14047 24191
rect 14047 24157 14056 24191
rect 14004 24148 14056 24157
rect 16120 24148 16172 24200
rect 16488 24148 16540 24200
rect 18420 24191 18472 24200
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 12348 24012 12400 24064
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 17684 24080 17736 24132
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 15752 24012 15804 24064
rect 17776 24055 17828 24064
rect 17776 24021 17785 24055
rect 17785 24021 17819 24055
rect 17819 24021 17828 24055
rect 17776 24012 17828 24021
rect 18880 24055 18932 24064
rect 18880 24021 18889 24055
rect 18889 24021 18923 24055
rect 18923 24021 18932 24055
rect 18880 24012 18932 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 11428 23851 11480 23860
rect 11428 23817 11437 23851
rect 11437 23817 11471 23851
rect 11471 23817 11480 23851
rect 11428 23808 11480 23817
rect 11796 23851 11848 23860
rect 11796 23817 11805 23851
rect 11805 23817 11839 23851
rect 11839 23817 11848 23851
rect 11796 23808 11848 23817
rect 13728 23808 13780 23860
rect 16120 23808 16172 23860
rect 16304 23851 16356 23860
rect 16304 23817 16313 23851
rect 16313 23817 16347 23851
rect 16347 23817 16356 23851
rect 16304 23808 16356 23817
rect 17040 23851 17092 23860
rect 17040 23817 17049 23851
rect 17049 23817 17083 23851
rect 17083 23817 17092 23851
rect 17040 23808 17092 23817
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 15752 23672 15804 23724
rect 18880 23715 18932 23724
rect 18880 23681 18889 23715
rect 18889 23681 18923 23715
rect 18923 23681 18932 23715
rect 18880 23672 18932 23681
rect 21732 23672 21784 23724
rect 24216 23672 24268 23724
rect 11336 23604 11388 23656
rect 12256 23604 12308 23656
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 12716 23647 12768 23656
rect 12716 23613 12750 23647
rect 12750 23613 12768 23647
rect 12716 23604 12768 23613
rect 16212 23604 16264 23656
rect 18420 23579 18472 23588
rect 18420 23545 18429 23579
rect 18429 23545 18463 23579
rect 18463 23545 18472 23579
rect 18420 23536 18472 23545
rect 19248 23536 19300 23588
rect 21640 23604 21692 23656
rect 21916 23536 21968 23588
rect 22928 23536 22980 23588
rect 8392 23468 8444 23520
rect 9588 23468 9640 23520
rect 12072 23468 12124 23520
rect 13452 23468 13504 23520
rect 14004 23468 14056 23520
rect 15292 23511 15344 23520
rect 15292 23477 15301 23511
rect 15301 23477 15335 23511
rect 15335 23477 15344 23511
rect 15292 23468 15344 23477
rect 16672 23511 16724 23520
rect 16672 23477 16681 23511
rect 16681 23477 16715 23511
rect 16715 23477 16724 23511
rect 16672 23468 16724 23477
rect 18328 23468 18380 23520
rect 20628 23468 20680 23520
rect 20812 23511 20864 23520
rect 20812 23477 20821 23511
rect 20821 23477 20855 23511
rect 20855 23477 20864 23511
rect 20812 23468 20864 23477
rect 21088 23468 21140 23520
rect 21364 23511 21416 23520
rect 21364 23477 21373 23511
rect 21373 23477 21407 23511
rect 21407 23477 21416 23511
rect 21364 23468 21416 23477
rect 22376 23511 22428 23520
rect 22376 23477 22385 23511
rect 22385 23477 22419 23511
rect 22419 23477 22428 23511
rect 22376 23468 22428 23477
rect 23112 23468 23164 23520
rect 24124 23468 24176 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 13360 23264 13412 23316
rect 15752 23264 15804 23316
rect 16580 23264 16632 23316
rect 17408 23264 17460 23316
rect 17684 23307 17736 23316
rect 17684 23273 17693 23307
rect 17693 23273 17727 23307
rect 17727 23273 17736 23307
rect 17684 23264 17736 23273
rect 18144 23307 18196 23316
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 19340 23264 19392 23316
rect 21640 23264 21692 23316
rect 23388 23307 23440 23316
rect 23388 23273 23397 23307
rect 23397 23273 23431 23307
rect 23431 23273 23440 23307
rect 23388 23264 23440 23273
rect 23664 23264 23716 23316
rect 24032 23307 24084 23316
rect 24032 23273 24041 23307
rect 24041 23273 24075 23307
rect 24075 23273 24084 23307
rect 24032 23264 24084 23273
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 12440 23196 12492 23248
rect 10876 23171 10928 23180
rect 10876 23137 10910 23171
rect 10910 23137 10928 23171
rect 16396 23196 16448 23248
rect 10876 23128 10928 23137
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 15844 23128 15896 23180
rect 18880 23196 18932 23248
rect 13820 23060 13872 23112
rect 14188 23103 14240 23112
rect 14188 23069 14197 23103
rect 14197 23069 14231 23103
rect 14231 23069 14240 23103
rect 14188 23060 14240 23069
rect 17408 23060 17460 23112
rect 20996 23128 21048 23180
rect 24676 23128 24728 23180
rect 20720 23060 20772 23112
rect 23020 23060 23072 23112
rect 23940 23060 23992 23112
rect 20904 23035 20956 23044
rect 20904 23001 20913 23035
rect 20913 23001 20947 23035
rect 20947 23001 20956 23035
rect 20904 22992 20956 23001
rect 11980 22967 12032 22976
rect 11980 22933 11989 22967
rect 11989 22933 12023 22967
rect 12023 22933 12032 22967
rect 11980 22924 12032 22933
rect 13084 22967 13136 22976
rect 13084 22933 13093 22967
rect 13093 22933 13127 22967
rect 13127 22933 13136 22967
rect 13084 22924 13136 22933
rect 14832 22924 14884 22976
rect 15292 22924 15344 22976
rect 21732 22924 21784 22976
rect 21916 22967 21968 22976
rect 21916 22933 21925 22967
rect 21925 22933 21959 22967
rect 21959 22933 21968 22967
rect 21916 22924 21968 22933
rect 22468 22924 22520 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10876 22720 10928 22772
rect 13820 22763 13872 22772
rect 13820 22729 13829 22763
rect 13829 22729 13863 22763
rect 13863 22729 13872 22763
rect 13820 22720 13872 22729
rect 15844 22720 15896 22772
rect 16396 22763 16448 22772
rect 16396 22729 16405 22763
rect 16405 22729 16439 22763
rect 16439 22729 16448 22763
rect 16396 22720 16448 22729
rect 16488 22720 16540 22772
rect 17040 22763 17092 22772
rect 17040 22729 17049 22763
rect 17049 22729 17083 22763
rect 17083 22729 17092 22763
rect 17040 22720 17092 22729
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 18052 22763 18104 22772
rect 18052 22729 18061 22763
rect 18061 22729 18095 22763
rect 18095 22729 18104 22763
rect 18052 22720 18104 22729
rect 18880 22720 18932 22772
rect 10600 22584 10652 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 15752 22584 15804 22636
rect 16396 22516 16448 22568
rect 17408 22652 17460 22704
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 21916 22720 21968 22772
rect 23020 22763 23072 22772
rect 23020 22729 23029 22763
rect 23029 22729 23063 22763
rect 23063 22729 23072 22763
rect 23020 22720 23072 22729
rect 23388 22720 23440 22772
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 16764 22516 16816 22568
rect 17500 22516 17552 22568
rect 18144 22516 18196 22568
rect 20904 22516 20956 22568
rect 23296 22584 23348 22636
rect 23388 22584 23440 22636
rect 23940 22584 23992 22636
rect 24032 22559 24084 22568
rect 24032 22525 24041 22559
rect 24041 22525 24075 22559
rect 24075 22525 24084 22559
rect 24032 22516 24084 22525
rect 13452 22448 13504 22500
rect 20260 22448 20312 22500
rect 21732 22448 21784 22500
rect 23112 22448 23164 22500
rect 14924 22423 14976 22432
rect 14924 22389 14933 22423
rect 14933 22389 14967 22423
rect 14967 22389 14976 22423
rect 14924 22380 14976 22389
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 15384 22423 15436 22432
rect 15384 22389 15393 22423
rect 15393 22389 15427 22423
rect 15427 22389 15436 22423
rect 15384 22380 15436 22389
rect 23296 22380 23348 22432
rect 23664 22423 23716 22432
rect 23664 22389 23673 22423
rect 23673 22389 23707 22423
rect 23707 22389 23716 22423
rect 23664 22380 23716 22389
rect 23756 22380 23808 22432
rect 24216 22380 24268 22432
rect 24676 22423 24728 22432
rect 24676 22389 24685 22423
rect 24685 22389 24719 22423
rect 24719 22389 24728 22423
rect 24676 22380 24728 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 13544 22176 13596 22228
rect 16672 22176 16724 22228
rect 18512 22176 18564 22228
rect 18972 22219 19024 22228
rect 18972 22185 18981 22219
rect 18981 22185 19015 22219
rect 19015 22185 19024 22219
rect 18972 22176 19024 22185
rect 19156 22176 19208 22228
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 20720 22219 20772 22228
rect 20720 22185 20729 22219
rect 20729 22185 20763 22219
rect 20763 22185 20772 22219
rect 20720 22176 20772 22185
rect 21640 22219 21692 22228
rect 21640 22185 21649 22219
rect 21649 22185 21683 22219
rect 21683 22185 21692 22219
rect 21640 22176 21692 22185
rect 23388 22176 23440 22228
rect 13820 22108 13872 22160
rect 14924 22108 14976 22160
rect 12440 22040 12492 22092
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 13544 22040 13596 22092
rect 13452 22015 13504 22024
rect 13452 21981 13461 22015
rect 13461 21981 13495 22015
rect 13495 21981 13504 22015
rect 13452 21972 13504 21981
rect 14648 21972 14700 22024
rect 17316 22083 17368 22092
rect 17316 22049 17325 22083
rect 17325 22049 17359 22083
rect 17359 22049 17368 22083
rect 17316 22040 17368 22049
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 16304 21972 16356 22024
rect 16580 21972 16632 22024
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 16856 21904 16908 21956
rect 18144 21972 18196 22024
rect 19248 22040 19300 22092
rect 21272 22040 21324 22092
rect 22100 22083 22152 22092
rect 22100 22049 22109 22083
rect 22109 22049 22143 22083
rect 22143 22049 22152 22083
rect 23664 22108 23716 22160
rect 23388 22083 23440 22092
rect 22100 22040 22152 22049
rect 18696 21904 18748 21956
rect 21180 21972 21232 22024
rect 21916 21972 21968 22024
rect 22376 21972 22428 22024
rect 23388 22049 23422 22083
rect 23422 22049 23440 22083
rect 23388 22040 23440 22049
rect 24124 22040 24176 22092
rect 24584 22040 24636 22092
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 11980 21836 12032 21888
rect 12164 21879 12216 21888
rect 12164 21845 12173 21879
rect 12173 21845 12207 21879
rect 12207 21845 12216 21879
rect 12164 21836 12216 21845
rect 15292 21836 15344 21888
rect 17132 21836 17184 21888
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 21916 21836 21968 21888
rect 23296 21836 23348 21888
rect 24216 21836 24268 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10600 21675 10652 21684
rect 10600 21641 10609 21675
rect 10609 21641 10643 21675
rect 10643 21641 10652 21675
rect 10600 21632 10652 21641
rect 13452 21675 13504 21684
rect 13452 21641 13461 21675
rect 13461 21641 13495 21675
rect 13495 21641 13504 21675
rect 13452 21632 13504 21641
rect 14648 21632 14700 21684
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 16304 21675 16356 21684
rect 16304 21641 16313 21675
rect 16313 21641 16347 21675
rect 16347 21641 16356 21675
rect 16304 21632 16356 21641
rect 16856 21675 16908 21684
rect 16856 21641 16865 21675
rect 16865 21641 16899 21675
rect 16899 21641 16908 21675
rect 16856 21632 16908 21641
rect 17408 21675 17460 21684
rect 17408 21641 17417 21675
rect 17417 21641 17451 21675
rect 17451 21641 17460 21675
rect 17408 21632 17460 21641
rect 18880 21675 18932 21684
rect 18880 21641 18889 21675
rect 18889 21641 18923 21675
rect 18923 21641 18932 21675
rect 18880 21632 18932 21641
rect 20260 21632 20312 21684
rect 22100 21632 22152 21684
rect 11980 21496 12032 21548
rect 14004 21496 14056 21548
rect 16028 21496 16080 21548
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 23756 21496 23808 21548
rect 12164 21428 12216 21480
rect 12716 21428 12768 21480
rect 14372 21428 14424 21480
rect 14740 21428 14792 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 19616 21428 19668 21480
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 12532 21360 12584 21412
rect 10784 21335 10836 21344
rect 10784 21301 10793 21335
rect 10793 21301 10827 21335
rect 10827 21301 10836 21335
rect 10784 21292 10836 21301
rect 11060 21292 11112 21344
rect 11244 21292 11296 21344
rect 12624 21292 12676 21344
rect 12716 21292 12768 21344
rect 13728 21292 13780 21344
rect 14924 21335 14976 21344
rect 14924 21301 14933 21335
rect 14933 21301 14967 21335
rect 14967 21301 14976 21335
rect 14924 21292 14976 21301
rect 17224 21292 17276 21344
rect 17316 21292 17368 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18144 21292 18196 21344
rect 21272 21292 21324 21344
rect 21824 21292 21876 21344
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 23848 21292 23900 21344
rect 24216 21428 24268 21480
rect 25504 21335 25556 21344
rect 25504 21301 25513 21335
rect 25513 21301 25547 21335
rect 25547 21301 25556 21335
rect 25504 21292 25556 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 13820 21131 13872 21140
rect 13820 21097 13829 21131
rect 13829 21097 13863 21131
rect 13863 21097 13872 21131
rect 13820 21088 13872 21097
rect 14832 21088 14884 21140
rect 15292 21088 15344 21140
rect 17132 21131 17184 21140
rect 17132 21097 17141 21131
rect 17141 21097 17175 21131
rect 17175 21097 17184 21131
rect 17132 21088 17184 21097
rect 22100 21088 22152 21140
rect 23388 21088 23440 21140
rect 23756 21131 23808 21140
rect 23756 21097 23765 21131
rect 23765 21097 23799 21131
rect 23799 21097 23808 21131
rect 23756 21088 23808 21097
rect 11980 21020 12032 21072
rect 19156 21020 19208 21072
rect 22928 21020 22980 21072
rect 23572 21020 23624 21072
rect 1952 20952 2004 21004
rect 15660 20952 15712 21004
rect 18604 20952 18656 21004
rect 19248 20995 19300 21004
rect 19248 20961 19257 20995
rect 19257 20961 19291 20995
rect 19291 20961 19300 20995
rect 19248 20952 19300 20961
rect 22100 20995 22152 21004
rect 22100 20961 22134 20995
rect 22134 20961 22152 20995
rect 22100 20952 22152 20961
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 15292 20884 15344 20936
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 17868 20927 17920 20936
rect 17868 20893 17877 20927
rect 17877 20893 17911 20927
rect 17911 20893 17920 20927
rect 17868 20884 17920 20893
rect 20260 20884 20312 20936
rect 21824 20927 21876 20936
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 23756 20884 23808 20936
rect 1584 20859 1636 20868
rect 1584 20825 1593 20859
rect 1593 20825 1627 20859
rect 1627 20825 1636 20859
rect 1584 20816 1636 20825
rect 25504 20884 25556 20936
rect 25136 20816 25188 20868
rect 11060 20748 11112 20800
rect 11704 20748 11756 20800
rect 13176 20748 13228 20800
rect 15752 20748 15804 20800
rect 17960 20748 18012 20800
rect 20444 20748 20496 20800
rect 24124 20791 24176 20800
rect 24124 20757 24133 20791
rect 24133 20757 24167 20791
rect 24167 20757 24176 20791
rect 24124 20748 24176 20757
rect 24216 20748 24268 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 11980 20544 12032 20596
rect 12532 20544 12584 20596
rect 16028 20544 16080 20596
rect 17868 20544 17920 20596
rect 19524 20544 19576 20596
rect 20260 20544 20312 20596
rect 22100 20544 22152 20596
rect 23572 20544 23624 20596
rect 24032 20544 24084 20596
rect 25320 20544 25372 20596
rect 25504 20587 25556 20596
rect 25504 20553 25513 20587
rect 25513 20553 25547 20587
rect 25547 20553 25556 20587
rect 25504 20544 25556 20553
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 13176 20408 13228 20460
rect 20720 20408 20772 20460
rect 25044 20408 25096 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 15476 20340 15528 20392
rect 18880 20340 18932 20392
rect 21640 20340 21692 20392
rect 24124 20340 24176 20392
rect 13268 20272 13320 20324
rect 18696 20272 18748 20324
rect 24860 20272 24912 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 10968 20204 11020 20256
rect 11336 20247 11388 20256
rect 11336 20213 11345 20247
rect 11345 20213 11379 20247
rect 11379 20213 11388 20247
rect 11336 20204 11388 20213
rect 11428 20204 11480 20256
rect 11888 20247 11940 20256
rect 11888 20213 11897 20247
rect 11897 20213 11931 20247
rect 11931 20213 11940 20247
rect 11888 20204 11940 20213
rect 13176 20204 13228 20256
rect 14188 20247 14240 20256
rect 14188 20213 14197 20247
rect 14197 20213 14231 20247
rect 14231 20213 14240 20247
rect 14188 20204 14240 20213
rect 14372 20204 14424 20256
rect 15292 20204 15344 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 21824 20247 21876 20256
rect 21824 20213 21833 20247
rect 21833 20213 21867 20247
rect 21867 20213 21876 20247
rect 21824 20204 21876 20213
rect 23940 20247 23992 20256
rect 23940 20213 23949 20247
rect 23949 20213 23983 20247
rect 23983 20213 23992 20247
rect 23940 20204 23992 20213
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 25136 20247 25188 20256
rect 25136 20213 25145 20247
rect 25145 20213 25179 20247
rect 25179 20213 25188 20247
rect 25136 20204 25188 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 11336 20000 11388 20052
rect 12532 20000 12584 20052
rect 14004 20000 14056 20052
rect 17868 20000 17920 20052
rect 18052 20043 18104 20052
rect 18052 20009 18061 20043
rect 18061 20009 18095 20043
rect 18095 20009 18104 20043
rect 18052 20000 18104 20009
rect 19248 20000 19300 20052
rect 20904 20000 20956 20052
rect 22100 20000 22152 20052
rect 24124 20000 24176 20052
rect 9864 19864 9916 19916
rect 11428 19932 11480 19984
rect 13176 19932 13228 19984
rect 16028 19932 16080 19984
rect 19524 19932 19576 19984
rect 20536 19932 20588 19984
rect 25044 19932 25096 19984
rect 10324 19864 10376 19916
rect 11244 19864 11296 19916
rect 11888 19864 11940 19916
rect 13544 19864 13596 19916
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 20076 19864 20128 19916
rect 20628 19864 20680 19916
rect 20996 19864 21048 19916
rect 23848 19864 23900 19916
rect 19248 19796 19300 19848
rect 19432 19796 19484 19848
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 1400 19660 1452 19712
rect 11612 19703 11664 19712
rect 11612 19669 11621 19703
rect 11621 19669 11655 19703
rect 11655 19669 11664 19703
rect 11612 19660 11664 19669
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 16856 19703 16908 19712
rect 16856 19669 16865 19703
rect 16865 19669 16899 19703
rect 16899 19669 16908 19703
rect 16856 19660 16908 19669
rect 25320 19703 25372 19712
rect 25320 19669 25329 19703
rect 25329 19669 25363 19703
rect 25363 19669 25372 19703
rect 25320 19660 25372 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 10324 19456 10376 19508
rect 13544 19499 13596 19508
rect 13544 19465 13553 19499
rect 13553 19465 13587 19499
rect 13587 19465 13596 19499
rect 13544 19456 13596 19465
rect 9864 19431 9916 19440
rect 9864 19397 9873 19431
rect 9873 19397 9907 19431
rect 9907 19397 9916 19431
rect 9864 19388 9916 19397
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 11612 19320 11664 19372
rect 9680 19252 9732 19304
rect 13176 19320 13228 19372
rect 15660 19456 15712 19508
rect 16028 19456 16080 19508
rect 18604 19456 18656 19508
rect 21272 19499 21324 19508
rect 21272 19465 21281 19499
rect 21281 19465 21315 19499
rect 21315 19465 21324 19499
rect 21272 19456 21324 19465
rect 22100 19456 22152 19508
rect 15476 19388 15528 19440
rect 16120 19431 16172 19440
rect 16120 19397 16129 19431
rect 16129 19397 16163 19431
rect 16163 19397 16172 19431
rect 16120 19388 16172 19397
rect 20904 19431 20956 19440
rect 20904 19397 20913 19431
rect 20913 19397 20947 19431
rect 20947 19397 20956 19431
rect 20904 19388 20956 19397
rect 21824 19388 21876 19440
rect 16028 19320 16080 19372
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 12532 19252 12584 19304
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 18052 19252 18104 19304
rect 14648 19184 14700 19236
rect 10692 19116 10744 19168
rect 10876 19116 10928 19168
rect 12716 19116 12768 19168
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 14188 19116 14240 19168
rect 17776 19184 17828 19236
rect 16948 19116 17000 19168
rect 18696 19116 18748 19168
rect 19156 19159 19208 19168
rect 19156 19125 19165 19159
rect 19165 19125 19199 19159
rect 19199 19125 19208 19159
rect 20996 19320 21048 19372
rect 22928 19388 22980 19440
rect 24860 19456 24912 19508
rect 25044 19499 25096 19508
rect 25044 19465 25053 19499
rect 25053 19465 25087 19499
rect 25087 19465 25096 19499
rect 25044 19456 25096 19465
rect 23940 19388 23992 19440
rect 24308 19388 24360 19440
rect 24584 19363 24636 19372
rect 20076 19295 20128 19304
rect 20076 19261 20085 19295
rect 20085 19261 20119 19295
rect 20119 19261 20128 19295
rect 20076 19252 20128 19261
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 25320 19320 25372 19372
rect 24124 19252 24176 19304
rect 25504 19295 25556 19304
rect 25504 19261 25513 19295
rect 25513 19261 25547 19295
rect 25547 19261 25556 19295
rect 25504 19252 25556 19261
rect 23848 19184 23900 19236
rect 24216 19184 24268 19236
rect 19156 19116 19208 19125
rect 19432 19116 19484 19168
rect 19984 19116 20036 19168
rect 20076 19116 20128 19168
rect 21640 19159 21692 19168
rect 21640 19125 21649 19159
rect 21649 19125 21683 19159
rect 21683 19125 21692 19159
rect 21640 19116 21692 19125
rect 22744 19159 22796 19168
rect 22744 19125 22753 19159
rect 22753 19125 22787 19159
rect 22787 19125 22796 19159
rect 22744 19116 22796 19125
rect 23940 19159 23992 19168
rect 23940 19125 23949 19159
rect 23949 19125 23983 19159
rect 23983 19125 23992 19159
rect 23940 19116 23992 19125
rect 25688 19159 25740 19168
rect 25688 19125 25697 19159
rect 25697 19125 25731 19159
rect 25731 19125 25740 19159
rect 25688 19116 25740 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 12808 18955 12860 18964
rect 12808 18921 12817 18955
rect 12817 18921 12851 18955
rect 12851 18921 12860 18955
rect 12808 18912 12860 18921
rect 13176 18955 13228 18964
rect 13176 18921 13185 18955
rect 13185 18921 13219 18955
rect 13219 18921 13228 18955
rect 13176 18912 13228 18921
rect 13728 18912 13780 18964
rect 13912 18912 13964 18964
rect 14648 18955 14700 18964
rect 14648 18921 14657 18955
rect 14657 18921 14691 18955
rect 14691 18921 14700 18955
rect 14648 18912 14700 18921
rect 16672 18912 16724 18964
rect 19156 18912 19208 18964
rect 19524 18955 19576 18964
rect 19524 18921 19533 18955
rect 19533 18921 19567 18955
rect 19567 18921 19576 18955
rect 19524 18912 19576 18921
rect 19984 18912 20036 18964
rect 21640 18912 21692 18964
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 13820 18844 13872 18896
rect 15752 18887 15804 18896
rect 15752 18853 15761 18887
rect 15761 18853 15795 18887
rect 15795 18853 15804 18887
rect 15752 18844 15804 18853
rect 19432 18844 19484 18896
rect 20076 18844 20128 18896
rect 21548 18887 21600 18896
rect 21548 18853 21557 18887
rect 21557 18853 21591 18887
rect 21591 18853 21600 18887
rect 21548 18844 21600 18853
rect 24308 18912 24360 18964
rect 24216 18844 24268 18896
rect 24584 18844 24636 18896
rect 10324 18776 10376 18828
rect 10968 18819 11020 18828
rect 10968 18785 10991 18819
rect 10991 18785 11020 18819
rect 10968 18776 11020 18785
rect 14004 18776 14056 18828
rect 15292 18776 15344 18828
rect 16580 18776 16632 18828
rect 17684 18776 17736 18828
rect 19248 18776 19300 18828
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 22560 18776 22612 18828
rect 23020 18776 23072 18828
rect 23480 18776 23532 18828
rect 10600 18708 10652 18760
rect 13820 18708 13872 18760
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 16120 18708 16172 18760
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 21180 18708 21232 18760
rect 21456 18708 21508 18760
rect 20996 18640 21048 18692
rect 22744 18708 22796 18760
rect 23388 18708 23440 18760
rect 23848 18751 23900 18760
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 10876 18572 10928 18624
rect 11428 18572 11480 18624
rect 14832 18572 14884 18624
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 25228 18615 25280 18624
rect 25228 18581 25237 18615
rect 25237 18581 25271 18615
rect 25271 18581 25280 18615
rect 25228 18572 25280 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 13912 18368 13964 18420
rect 14648 18368 14700 18420
rect 15844 18368 15896 18420
rect 16028 18368 16080 18420
rect 16856 18368 16908 18420
rect 17684 18411 17736 18420
rect 17684 18377 17693 18411
rect 17693 18377 17727 18411
rect 17727 18377 17736 18411
rect 17684 18368 17736 18377
rect 20444 18368 20496 18420
rect 22744 18368 22796 18420
rect 23204 18368 23256 18420
rect 10692 18232 10744 18284
rect 16580 18300 16632 18352
rect 17132 18300 17184 18352
rect 11428 18275 11480 18284
rect 11428 18241 11437 18275
rect 11437 18241 11471 18275
rect 11471 18241 11480 18275
rect 11428 18232 11480 18241
rect 13636 18232 13688 18284
rect 14004 18232 14056 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23848 18368 23900 18420
rect 24676 18232 24728 18284
rect 25228 18368 25280 18420
rect 12808 18164 12860 18216
rect 14372 18207 14424 18216
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 16580 18164 16632 18216
rect 21180 18207 21232 18216
rect 21180 18173 21189 18207
rect 21189 18173 21223 18207
rect 21223 18173 21232 18207
rect 21180 18164 21232 18173
rect 23664 18164 23716 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 12440 18096 12492 18148
rect 13268 18139 13320 18148
rect 13268 18105 13277 18139
rect 13277 18105 13311 18139
rect 13311 18105 13320 18139
rect 13268 18096 13320 18105
rect 14188 18096 14240 18148
rect 14832 18096 14884 18148
rect 19064 18096 19116 18148
rect 20720 18096 20772 18148
rect 22192 18096 22244 18148
rect 23204 18096 23256 18148
rect 23572 18096 23624 18148
rect 10968 18028 11020 18080
rect 11152 18071 11204 18080
rect 11152 18037 11161 18071
rect 11161 18037 11195 18071
rect 11195 18037 11204 18071
rect 11152 18028 11204 18037
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 17224 18028 17276 18080
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 23664 18071 23716 18080
rect 23664 18037 23673 18071
rect 23673 18037 23707 18071
rect 23707 18037 23716 18071
rect 23664 18028 23716 18037
rect 25412 18071 25464 18080
rect 25412 18037 25421 18071
rect 25421 18037 25455 18071
rect 25455 18037 25464 18071
rect 25412 18028 25464 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 13728 17867 13780 17876
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 20076 17824 20128 17876
rect 20352 17867 20404 17876
rect 20352 17833 20361 17867
rect 20361 17833 20395 17867
rect 20395 17833 20404 17867
rect 20352 17824 20404 17833
rect 21548 17824 21600 17876
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 24216 17867 24268 17876
rect 24216 17833 24225 17867
rect 24225 17833 24259 17867
rect 24259 17833 24268 17867
rect 24216 17824 24268 17833
rect 11428 17756 11480 17808
rect 14556 17756 14608 17808
rect 15660 17799 15712 17808
rect 15660 17765 15669 17799
rect 15669 17765 15703 17799
rect 15703 17765 15712 17799
rect 15660 17756 15712 17765
rect 17408 17756 17460 17808
rect 22468 17756 22520 17808
rect 23204 17756 23256 17808
rect 23296 17756 23348 17808
rect 10692 17688 10744 17740
rect 11796 17688 11848 17740
rect 17040 17688 17092 17740
rect 19800 17731 19852 17740
rect 19800 17697 19809 17731
rect 19809 17697 19843 17731
rect 19843 17697 19852 17731
rect 19800 17688 19852 17697
rect 20720 17688 20772 17740
rect 23572 17731 23624 17740
rect 23572 17697 23581 17731
rect 23581 17697 23615 17731
rect 23615 17697 23624 17731
rect 23572 17688 23624 17697
rect 25596 17688 25648 17740
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 14556 17620 14608 17672
rect 21640 17620 21692 17672
rect 23296 17620 23348 17672
rect 16028 17552 16080 17604
rect 22192 17552 22244 17604
rect 23204 17595 23256 17604
rect 23204 17561 23213 17595
rect 23213 17561 23247 17595
rect 23247 17561 23256 17595
rect 23204 17552 23256 17561
rect 23940 17552 23992 17604
rect 24584 17552 24636 17604
rect 12716 17484 12768 17536
rect 14188 17484 14240 17536
rect 14372 17484 14424 17536
rect 14832 17484 14884 17536
rect 15384 17484 15436 17536
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 13820 17323 13872 17332
rect 11244 17144 11296 17196
rect 11428 17187 11480 17196
rect 11428 17153 11437 17187
rect 11437 17153 11471 17187
rect 11471 17153 11480 17187
rect 11428 17144 11480 17153
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 14648 17280 14700 17332
rect 16028 17280 16080 17332
rect 17040 17323 17092 17332
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 20444 17280 20496 17332
rect 20996 17280 21048 17332
rect 21824 17280 21876 17332
rect 22284 17280 22336 17332
rect 22468 17323 22520 17332
rect 22468 17289 22477 17323
rect 22477 17289 22511 17323
rect 22511 17289 22520 17323
rect 22468 17280 22520 17289
rect 23296 17280 23348 17332
rect 25596 17323 25648 17332
rect 25596 17289 25605 17323
rect 25605 17289 25639 17323
rect 25639 17289 25648 17323
rect 25596 17280 25648 17289
rect 16120 17212 16172 17264
rect 16396 17212 16448 17264
rect 20904 17212 20956 17264
rect 20720 17144 20772 17196
rect 21640 17187 21692 17196
rect 21640 17153 21649 17187
rect 21649 17153 21683 17187
rect 21683 17153 21692 17187
rect 21640 17144 21692 17153
rect 11336 17008 11388 17060
rect 12716 17119 12768 17128
rect 12716 17085 12750 17119
rect 12750 17085 12768 17119
rect 12716 17076 12768 17085
rect 14832 17051 14884 17060
rect 14832 17017 14841 17051
rect 14841 17017 14875 17051
rect 14875 17017 14884 17051
rect 15016 17076 15068 17128
rect 20812 17076 20864 17128
rect 22100 17076 22152 17128
rect 24676 17076 24728 17128
rect 14832 17008 14884 17017
rect 16948 17008 17000 17060
rect 18880 17051 18932 17060
rect 18880 17017 18914 17051
rect 18914 17017 18932 17051
rect 18880 17008 18932 17017
rect 11060 16940 11112 16992
rect 11428 16940 11480 16992
rect 13544 16940 13596 16992
rect 14280 16940 14332 16992
rect 19064 16940 19116 16992
rect 20996 16940 21048 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 11244 16779 11296 16788
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 12440 16736 12492 16788
rect 11060 16668 11112 16720
rect 11336 16600 11388 16652
rect 12716 16736 12768 16788
rect 14372 16779 14424 16788
rect 14372 16745 14381 16779
rect 14381 16745 14415 16779
rect 14415 16745 14424 16779
rect 14372 16736 14424 16745
rect 15016 16779 15068 16788
rect 15016 16745 15025 16779
rect 15025 16745 15059 16779
rect 15059 16745 15068 16779
rect 15016 16736 15068 16745
rect 11152 16532 11204 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 11888 16532 11940 16584
rect 14280 16600 14332 16652
rect 16304 16736 16356 16788
rect 18880 16779 18932 16788
rect 18880 16745 18889 16779
rect 18889 16745 18923 16779
rect 18923 16745 18932 16779
rect 18880 16736 18932 16745
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 22100 16736 22152 16788
rect 22376 16736 22428 16788
rect 23572 16736 23624 16788
rect 15384 16668 15436 16720
rect 17132 16711 17184 16720
rect 17132 16677 17166 16711
rect 17166 16677 17184 16711
rect 17132 16668 17184 16677
rect 18328 16668 18380 16720
rect 23204 16711 23256 16720
rect 23204 16677 23213 16711
rect 23213 16677 23247 16711
rect 23247 16677 23256 16711
rect 23204 16668 23256 16677
rect 23480 16668 23532 16720
rect 14832 16532 14884 16584
rect 14648 16464 14700 16516
rect 16948 16600 17000 16652
rect 20628 16600 20680 16652
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 21640 16600 21692 16652
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 23848 16575 23900 16584
rect 20904 16532 20956 16541
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 24216 16532 24268 16584
rect 24676 16736 24728 16788
rect 25136 16779 25188 16788
rect 25136 16745 25145 16779
rect 25145 16745 25179 16779
rect 25179 16745 25188 16779
rect 25136 16736 25188 16745
rect 24860 16600 24912 16652
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 20444 16396 20496 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 11060 16192 11112 16244
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 14648 16235 14700 16244
rect 14648 16201 14657 16235
rect 14657 16201 14691 16235
rect 14691 16201 14700 16235
rect 14648 16192 14700 16201
rect 15844 16192 15896 16244
rect 16028 16192 16080 16244
rect 11796 16124 11848 16176
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 16948 16192 17000 16244
rect 17132 16192 17184 16244
rect 20536 16192 20588 16244
rect 20720 16192 20772 16244
rect 20904 16124 20956 16176
rect 17040 16099 17092 16108
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 16304 15988 16356 16040
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 19064 16056 19116 16108
rect 20444 16056 20496 16108
rect 13636 15920 13688 15972
rect 16948 15988 17000 16040
rect 20076 15988 20128 16040
rect 23480 16192 23532 16244
rect 24216 16235 24268 16244
rect 24216 16201 24225 16235
rect 24225 16201 24259 16235
rect 24259 16201 24268 16235
rect 24216 16192 24268 16201
rect 24860 16192 24912 16244
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22376 16099 22428 16108
rect 22192 16056 22244 16065
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 24216 16056 24268 16108
rect 25044 16056 25096 16108
rect 24124 15988 24176 16040
rect 13728 15852 13780 15904
rect 14556 15852 14608 15904
rect 16396 15895 16448 15904
rect 16396 15861 16405 15895
rect 16405 15861 16439 15895
rect 16439 15861 16448 15895
rect 16396 15852 16448 15861
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 19156 15920 19208 15972
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 19524 15852 19576 15904
rect 23020 15852 23072 15904
rect 23848 15852 23900 15904
rect 24768 15895 24820 15904
rect 24768 15861 24777 15895
rect 24777 15861 24811 15895
rect 24811 15861 24820 15895
rect 24768 15852 24820 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 14556 15648 14608 15700
rect 14832 15648 14884 15700
rect 17040 15691 17092 15700
rect 17040 15657 17049 15691
rect 17049 15657 17083 15691
rect 17083 15657 17092 15691
rect 17040 15648 17092 15657
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 20076 15648 20128 15700
rect 20444 15648 20496 15700
rect 21364 15580 21416 15632
rect 15660 15512 15712 15564
rect 14832 15444 14884 15496
rect 16396 15512 16448 15564
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 17408 15555 17460 15564
rect 17408 15521 17442 15555
rect 17442 15521 17460 15555
rect 17408 15512 17460 15521
rect 24032 15512 24084 15564
rect 16212 15487 16264 15496
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 19432 15444 19484 15496
rect 20904 15444 20956 15496
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 15292 15308 15344 15360
rect 16488 15308 16540 15360
rect 18236 15308 18288 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 14832 15104 14884 15156
rect 16396 15104 16448 15156
rect 17132 15104 17184 15156
rect 16212 14968 16264 15020
rect 16580 14968 16632 15020
rect 21732 15104 21784 15156
rect 22192 15104 22244 15156
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 24032 15104 24084 15156
rect 20904 15036 20956 15088
rect 23388 15036 23440 15088
rect 12624 14900 12676 14952
rect 17408 14900 17460 14952
rect 21456 14943 21508 14952
rect 21456 14909 21465 14943
rect 21465 14909 21499 14943
rect 21499 14909 21508 14943
rect 21456 14900 21508 14909
rect 24584 14943 24636 14952
rect 18236 14832 18288 14884
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 14832 14764 14884 14816
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 19984 14764 20036 14816
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 23756 14764 23808 14816
rect 24768 14807 24820 14816
rect 24768 14773 24777 14807
rect 24777 14773 24811 14807
rect 24811 14773 24820 14807
rect 24768 14764 24820 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 15200 14560 15252 14612
rect 16028 14560 16080 14612
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 18052 14603 18104 14612
rect 18052 14569 18061 14603
rect 18061 14569 18095 14603
rect 18095 14569 18104 14603
rect 18052 14560 18104 14569
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 21456 14603 21508 14612
rect 21456 14569 21465 14603
rect 21465 14569 21499 14603
rect 21499 14569 21508 14603
rect 21456 14560 21508 14569
rect 24860 14560 24912 14612
rect 15292 14492 15344 14544
rect 16212 14492 16264 14544
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 13176 14424 13228 14476
rect 15476 14424 15528 14476
rect 16764 14424 16816 14476
rect 17132 14424 17184 14476
rect 20904 14467 20956 14476
rect 20904 14433 20913 14467
rect 20913 14433 20947 14467
rect 20947 14433 20956 14467
rect 20904 14424 20956 14433
rect 21916 14424 21968 14476
rect 18052 14356 18104 14408
rect 14280 14331 14332 14340
rect 14280 14297 14289 14331
rect 14289 14297 14323 14331
rect 14323 14297 14332 14331
rect 14280 14288 14332 14297
rect 19340 14288 19392 14340
rect 19984 14288 20036 14340
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 18236 14220 18288 14272
rect 18972 14220 19024 14272
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 22744 14220 22796 14272
rect 24032 14424 24084 14476
rect 24400 14424 24452 14476
rect 25596 14424 25648 14476
rect 23848 14399 23900 14408
rect 23848 14365 23857 14399
rect 23857 14365 23891 14399
rect 23891 14365 23900 14399
rect 23848 14356 23900 14365
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 13176 14016 13228 14068
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 14832 14016 14884 14068
rect 16212 14016 16264 14068
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 19432 14016 19484 14068
rect 19616 14016 19668 14068
rect 20812 14016 20864 14068
rect 21364 14016 21416 14068
rect 23848 14016 23900 14068
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 16764 13991 16816 14000
rect 16764 13957 16773 13991
rect 16773 13957 16807 13991
rect 16807 13957 16816 13991
rect 16764 13948 16816 13957
rect 20904 13948 20956 14000
rect 21916 13948 21968 14000
rect 23388 13991 23440 14000
rect 23388 13957 23397 13991
rect 23397 13957 23431 13991
rect 23431 13957 23440 13991
rect 23388 13948 23440 13957
rect 14188 13812 14240 13864
rect 14464 13812 14516 13864
rect 14832 13812 14884 13864
rect 15384 13812 15436 13864
rect 18236 13880 18288 13932
rect 19340 13880 19392 13932
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 18144 13812 18196 13864
rect 19616 13855 19668 13864
rect 19616 13821 19625 13855
rect 19625 13821 19659 13855
rect 19659 13821 19668 13855
rect 19616 13812 19668 13821
rect 23572 13744 23624 13796
rect 24032 13744 24084 13796
rect 16856 13676 16908 13728
rect 17592 13676 17644 13728
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 21640 13676 21692 13728
rect 23112 13676 23164 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 14740 13472 14792 13524
rect 17132 13472 17184 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 19340 13472 19392 13524
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 23848 13472 23900 13524
rect 24216 13472 24268 13524
rect 24768 13515 24820 13524
rect 24768 13481 24777 13515
rect 24777 13481 24811 13515
rect 24811 13481 24820 13515
rect 24768 13472 24820 13481
rect 16212 13404 16264 13456
rect 19432 13404 19484 13456
rect 19616 13447 19668 13456
rect 19616 13413 19625 13447
rect 19625 13413 19659 13447
rect 19659 13413 19668 13447
rect 19616 13404 19668 13413
rect 23112 13447 23164 13456
rect 23112 13413 23121 13447
rect 23121 13413 23155 13447
rect 23155 13413 23164 13447
rect 23112 13404 23164 13413
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 16304 13336 16356 13388
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 18788 13336 18840 13388
rect 19524 13336 19576 13388
rect 21088 13336 21140 13388
rect 24584 13379 24636 13388
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 16212 13311 16264 13320
rect 16212 13277 16221 13311
rect 16221 13277 16255 13311
rect 16255 13277 16264 13311
rect 16212 13268 16264 13277
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 18420 13268 18472 13320
rect 20996 13268 21048 13320
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 21640 13268 21692 13320
rect 16764 13200 16816 13252
rect 19248 13243 19300 13252
rect 19248 13209 19257 13243
rect 19257 13209 19291 13243
rect 19291 13209 19300 13243
rect 19248 13200 19300 13209
rect 19340 13200 19392 13252
rect 22744 13243 22796 13252
rect 22744 13209 22753 13243
rect 22753 13209 22787 13243
rect 22787 13209 22796 13243
rect 22744 13200 22796 13209
rect 16948 13175 17000 13184
rect 16948 13141 16957 13175
rect 16957 13141 16991 13175
rect 16991 13141 17000 13175
rect 16948 13132 17000 13141
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20628 13132 20680 13141
rect 21916 13175 21968 13184
rect 21916 13141 21925 13175
rect 21925 13141 21959 13175
rect 21959 13141 21968 13175
rect 21916 13132 21968 13141
rect 22100 13132 22152 13184
rect 23572 13132 23624 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 15476 12928 15528 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 16856 12928 16908 12980
rect 17684 12928 17736 12980
rect 20812 12928 20864 12980
rect 21364 12928 21416 12980
rect 21640 12928 21692 12980
rect 22284 12971 22336 12980
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 23112 12971 23164 12980
rect 23112 12937 23121 12971
rect 23121 12937 23155 12971
rect 23155 12937 23164 12971
rect 23112 12928 23164 12937
rect 24676 12928 24728 12980
rect 16304 12860 16356 12912
rect 19616 12860 19668 12912
rect 22560 12860 22612 12912
rect 23204 12860 23256 12912
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 21364 12792 21416 12844
rect 21916 12792 21968 12844
rect 16488 12724 16540 12776
rect 16948 12724 17000 12776
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 19340 12767 19392 12776
rect 19340 12733 19349 12767
rect 19349 12733 19383 12767
rect 19383 12733 19392 12767
rect 19340 12724 19392 12733
rect 20628 12724 20680 12776
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 24584 12767 24636 12776
rect 22100 12724 22152 12733
rect 24584 12733 24593 12767
rect 24593 12733 24627 12767
rect 24627 12733 24636 12767
rect 24584 12724 24636 12733
rect 12624 12656 12676 12708
rect 14372 12699 14424 12708
rect 14372 12665 14384 12699
rect 14384 12665 14424 12699
rect 14372 12656 14424 12665
rect 19248 12656 19300 12708
rect 20444 12656 20496 12708
rect 23020 12656 23072 12708
rect 12440 12588 12492 12640
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 17500 12588 17552 12640
rect 18052 12588 18104 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 19156 12588 19208 12640
rect 20536 12631 20588 12640
rect 20536 12597 20545 12631
rect 20545 12597 20579 12631
rect 20579 12597 20588 12631
rect 20536 12588 20588 12597
rect 21088 12588 21140 12640
rect 24768 12631 24820 12640
rect 24768 12597 24777 12631
rect 24777 12597 24811 12631
rect 24811 12597 24820 12631
rect 24768 12588 24820 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 13084 12384 13136 12436
rect 13544 12384 13596 12436
rect 16212 12384 16264 12436
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 19064 12384 19116 12436
rect 20536 12384 20588 12436
rect 23756 12427 23808 12436
rect 23756 12393 23765 12427
rect 23765 12393 23799 12427
rect 23799 12393 23808 12427
rect 23756 12384 23808 12393
rect 11612 12316 11664 12368
rect 13728 12316 13780 12368
rect 14280 12316 14332 12368
rect 14556 12316 14608 12368
rect 17132 12316 17184 12368
rect 19524 12316 19576 12368
rect 21364 12359 21416 12368
rect 21364 12325 21398 12359
rect 21398 12325 21416 12359
rect 21364 12316 21416 12325
rect 13176 12248 13228 12300
rect 15476 12248 15528 12300
rect 16304 12248 16356 12300
rect 19248 12248 19300 12300
rect 19984 12248 20036 12300
rect 20904 12248 20956 12300
rect 22744 12248 22796 12300
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13636 12180 13688 12232
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 20076 12180 20128 12232
rect 11704 12112 11756 12164
rect 14740 12112 14792 12164
rect 16856 12112 16908 12164
rect 23572 12112 23624 12164
rect 13176 12044 13228 12096
rect 14188 12044 14240 12096
rect 19248 12044 19300 12096
rect 19432 12044 19484 12096
rect 20444 12044 20496 12096
rect 22468 12087 22520 12096
rect 22468 12053 22477 12087
rect 22477 12053 22511 12087
rect 22511 12053 22520 12087
rect 22468 12044 22520 12053
rect 24216 12044 24268 12096
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 11612 11840 11664 11892
rect 12440 11840 12492 11892
rect 14280 11840 14332 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 16488 11840 16540 11892
rect 16580 11840 16632 11892
rect 20076 11883 20128 11892
rect 12624 11772 12676 11824
rect 16580 11704 16632 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 16948 11704 17000 11713
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 20904 11840 20956 11892
rect 21916 11883 21968 11892
rect 21916 11849 21925 11883
rect 21925 11849 21959 11883
rect 21959 11849 21968 11883
rect 21916 11840 21968 11849
rect 22744 11883 22796 11892
rect 22744 11849 22753 11883
rect 22753 11849 22787 11883
rect 22787 11849 22796 11883
rect 22744 11840 22796 11849
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 23940 11704 23992 11756
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 20536 11679 20588 11688
rect 20536 11645 20545 11679
rect 20545 11645 20579 11679
rect 20579 11645 20588 11679
rect 20536 11636 20588 11645
rect 14648 11568 14700 11620
rect 14924 11543 14976 11552
rect 14924 11509 14933 11543
rect 14933 11509 14967 11543
rect 14967 11509 14976 11543
rect 14924 11500 14976 11509
rect 16764 11500 16816 11552
rect 17592 11568 17644 11620
rect 18236 11568 18288 11620
rect 20260 11568 20312 11620
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 23664 11543 23716 11552
rect 23664 11509 23673 11543
rect 23673 11509 23707 11543
rect 23707 11509 23716 11543
rect 23664 11500 23716 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 12256 11296 12308 11348
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 14648 11339 14700 11348
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 16856 11296 16908 11348
rect 16948 11296 17000 11348
rect 19156 11296 19208 11348
rect 19432 11296 19484 11348
rect 19524 11296 19576 11348
rect 20628 11296 20680 11348
rect 20904 11296 20956 11348
rect 22008 11296 22060 11348
rect 11244 11160 11296 11212
rect 14004 11203 14056 11212
rect 14004 11169 14013 11203
rect 14013 11169 14047 11203
rect 14047 11169 14056 11203
rect 14004 11160 14056 11169
rect 15108 11160 15160 11212
rect 16488 11160 16540 11212
rect 16580 11160 16632 11212
rect 17132 11203 17184 11212
rect 17132 11169 17166 11203
rect 17166 11169 17184 11203
rect 17132 11160 17184 11169
rect 22468 11228 22520 11280
rect 25320 11228 25372 11280
rect 13728 11024 13780 11076
rect 14372 11092 14424 11144
rect 14924 11092 14976 11144
rect 16764 11092 16816 11144
rect 16304 11067 16356 11076
rect 16304 11033 16313 11067
rect 16313 11033 16347 11067
rect 16347 11033 16356 11067
rect 16304 11024 16356 11033
rect 18236 11067 18288 11076
rect 18236 11033 18245 11067
rect 18245 11033 18279 11067
rect 18279 11033 18288 11067
rect 18236 11024 18288 11033
rect 19984 11024 20036 11076
rect 1492 10956 1544 11008
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 12900 10956 12952 11008
rect 16764 10999 16816 11008
rect 16764 10965 16773 10999
rect 16773 10965 16807 10999
rect 16807 10965 16816 10999
rect 16764 10956 16816 10965
rect 20260 10956 20312 11008
rect 20720 10956 20772 11008
rect 22376 11160 22428 11212
rect 25596 11160 25648 11212
rect 21916 11092 21968 11144
rect 25412 11135 25464 11144
rect 25412 11101 25421 11135
rect 25421 11101 25455 11135
rect 25455 11101 25464 11135
rect 25412 11092 25464 11101
rect 24768 11067 24820 11076
rect 24768 11033 24777 11067
rect 24777 11033 24811 11067
rect 24811 11033 24820 11067
rect 24768 11024 24820 11033
rect 22100 10999 22152 11008
rect 22100 10965 22109 10999
rect 22109 10965 22143 10999
rect 22143 10965 22152 10999
rect 22100 10956 22152 10965
rect 23940 10956 23992 11008
rect 25412 10956 25464 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 11244 10795 11296 10804
rect 11244 10761 11253 10795
rect 11253 10761 11287 10795
rect 11287 10761 11296 10795
rect 11244 10752 11296 10761
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 13820 10752 13872 10804
rect 15292 10752 15344 10804
rect 16580 10752 16632 10804
rect 13452 10684 13504 10736
rect 17132 10752 17184 10804
rect 18880 10752 18932 10804
rect 20720 10752 20772 10804
rect 22376 10795 22428 10804
rect 22376 10761 22385 10795
rect 22385 10761 22419 10795
rect 22419 10761 22428 10795
rect 22376 10752 22428 10761
rect 22468 10752 22520 10804
rect 25412 10752 25464 10804
rect 23388 10727 23440 10736
rect 12532 10616 12584 10668
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 14464 10659 14516 10668
rect 13544 10616 13596 10625
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 14648 10659 14700 10668
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 16304 10616 16356 10668
rect 23388 10693 23397 10727
rect 23397 10693 23431 10727
rect 23431 10693 23440 10727
rect 23388 10684 23440 10693
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 1492 10548 1544 10600
rect 1676 10591 1728 10600
rect 1676 10557 1710 10591
rect 1710 10557 1728 10591
rect 1676 10548 1728 10557
rect 11336 10591 11388 10600
rect 11336 10557 11345 10591
rect 11345 10557 11379 10591
rect 11379 10557 11388 10591
rect 11336 10548 11388 10557
rect 12624 10548 12676 10600
rect 16672 10548 16724 10600
rect 19156 10591 19208 10600
rect 19156 10557 19190 10591
rect 19190 10557 19208 10591
rect 19156 10548 19208 10557
rect 23940 10591 23992 10600
rect 23940 10557 23974 10591
rect 23974 10557 23992 10591
rect 23940 10548 23992 10557
rect 11612 10480 11664 10532
rect 20720 10480 20772 10532
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 12900 10455 12952 10464
rect 2780 10412 2832 10421
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13544 10412 13596 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 16028 10412 16080 10464
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 21732 10455 21784 10464
rect 21732 10421 21741 10455
rect 21741 10421 21775 10455
rect 21775 10421 21784 10455
rect 21732 10412 21784 10421
rect 23480 10412 23532 10464
rect 24216 10412 24268 10464
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 14004 10208 14056 10260
rect 16304 10251 16356 10260
rect 16304 10217 16313 10251
rect 16313 10217 16347 10251
rect 16347 10217 16356 10251
rect 16304 10208 16356 10217
rect 16580 10208 16632 10260
rect 16764 10208 16816 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 21824 10208 21876 10260
rect 23020 10208 23072 10260
rect 11152 10140 11204 10192
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 11152 9868 11204 9877
rect 11336 9868 11388 9920
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 13728 10140 13780 10192
rect 13820 10072 13872 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15568 10004 15620 10056
rect 16304 10004 16356 10056
rect 17132 10004 17184 10056
rect 17408 10140 17460 10192
rect 23480 10140 23532 10192
rect 18788 10115 18840 10124
rect 18788 10081 18797 10115
rect 18797 10081 18831 10115
rect 18831 10081 18840 10115
rect 18788 10072 18840 10081
rect 19156 10072 19208 10124
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 18972 10047 19024 10056
rect 17408 10004 17460 10013
rect 18972 10013 18981 10047
rect 18981 10013 19015 10047
rect 19015 10013 19024 10047
rect 18972 10004 19024 10013
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 23388 10004 23440 10056
rect 13452 9936 13504 9988
rect 21732 9936 21784 9988
rect 11980 9868 12032 9920
rect 13636 9911 13688 9920
rect 13636 9877 13645 9911
rect 13645 9877 13679 9911
rect 13679 9877 13688 9911
rect 13636 9868 13688 9877
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 18328 9868 18380 9920
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 25320 9868 25372 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 14004 9707 14056 9716
rect 14004 9673 14013 9707
rect 14013 9673 14047 9707
rect 14047 9673 14056 9707
rect 14004 9664 14056 9673
rect 16304 9664 16356 9716
rect 16580 9664 16632 9716
rect 20720 9707 20772 9716
rect 11980 9596 12032 9648
rect 11796 9528 11848 9580
rect 16672 9596 16724 9648
rect 20720 9673 20729 9707
rect 20729 9673 20763 9707
rect 20763 9673 20772 9707
rect 20720 9664 20772 9673
rect 21364 9664 21416 9716
rect 21824 9664 21876 9716
rect 23388 9707 23440 9716
rect 23388 9673 23397 9707
rect 23397 9673 23431 9707
rect 23431 9673 23440 9707
rect 23388 9664 23440 9673
rect 9956 9460 10008 9512
rect 11980 9460 12032 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 13084 9460 13136 9512
rect 13728 9528 13780 9580
rect 14648 9528 14700 9580
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 21456 9596 21508 9648
rect 21640 9639 21692 9648
rect 21640 9605 21649 9639
rect 21649 9605 21683 9639
rect 21683 9605 21692 9639
rect 21640 9596 21692 9605
rect 17684 9528 17736 9580
rect 18236 9528 18288 9580
rect 18880 9528 18932 9580
rect 17040 9460 17092 9512
rect 20168 9460 20220 9512
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 24768 9460 24820 9512
rect 14832 9392 14884 9444
rect 15016 9435 15068 9444
rect 15016 9401 15050 9435
rect 15050 9401 15068 9435
rect 15016 9392 15068 9401
rect 17868 9435 17920 9444
rect 17868 9401 17877 9435
rect 17877 9401 17911 9435
rect 17911 9401 17920 9435
rect 17868 9392 17920 9401
rect 20812 9392 20864 9444
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 10876 9324 10928 9376
rect 11152 9324 11204 9376
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12808 9324 12860 9376
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 15568 9324 15620 9376
rect 16764 9324 16816 9376
rect 17132 9324 17184 9376
rect 18328 9324 18380 9376
rect 19156 9367 19208 9376
rect 19156 9333 19165 9367
rect 19165 9333 19199 9367
rect 19199 9333 19208 9367
rect 19156 9324 19208 9333
rect 21456 9324 21508 9376
rect 22284 9324 22336 9376
rect 23480 9392 23532 9444
rect 25504 9367 25556 9376
rect 25504 9333 25513 9367
rect 25513 9333 25547 9367
rect 25547 9333 25556 9367
rect 25504 9324 25556 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 12900 9120 12952 9172
rect 13728 9120 13780 9172
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 19432 9120 19484 9172
rect 20260 9120 20312 9172
rect 21548 9163 21600 9172
rect 21548 9129 21557 9163
rect 21557 9129 21591 9163
rect 21591 9129 21600 9163
rect 21548 9120 21600 9129
rect 22100 9120 22152 9172
rect 23664 9163 23716 9172
rect 23664 9129 23673 9163
rect 23673 9129 23707 9163
rect 23707 9129 23716 9163
rect 23664 9120 23716 9129
rect 24032 9120 24084 9172
rect 12072 9052 12124 9104
rect 12808 9052 12860 9104
rect 13452 9095 13504 9104
rect 13452 9061 13461 9095
rect 13461 9061 13495 9095
rect 13495 9061 13504 9095
rect 13452 9052 13504 9061
rect 14648 9052 14700 9104
rect 10876 8984 10928 9036
rect 9680 8916 9732 8968
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 12900 8984 12952 9036
rect 13176 8984 13228 9036
rect 14004 9027 14056 9036
rect 14004 8993 14013 9027
rect 14013 8993 14047 9027
rect 14047 8993 14056 9027
rect 14004 8984 14056 8993
rect 16212 9052 16264 9104
rect 17408 9052 17460 9104
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 18144 8984 18196 8993
rect 19340 8984 19392 9036
rect 21916 8984 21968 9036
rect 14372 8916 14424 8968
rect 17040 8916 17092 8968
rect 17776 8916 17828 8968
rect 22192 8916 22244 8968
rect 23296 8959 23348 8968
rect 16580 8848 16632 8900
rect 17224 8891 17276 8900
rect 17224 8857 17233 8891
rect 17233 8857 17267 8891
rect 17267 8857 17276 8891
rect 17224 8848 17276 8857
rect 20168 8848 20220 8900
rect 23296 8925 23305 8959
rect 23305 8925 23339 8959
rect 23339 8925 23348 8959
rect 24768 9052 24820 9104
rect 24860 8984 24912 9036
rect 24676 8959 24728 8968
rect 23296 8916 23348 8925
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24676 8916 24728 8925
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 13360 8780 13412 8832
rect 15476 8780 15528 8832
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 22376 8780 22428 8832
rect 23572 8780 23624 8832
rect 24768 8780 24820 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 14372 8619 14424 8628
rect 14372 8585 14381 8619
rect 14381 8585 14415 8619
rect 14415 8585 14424 8619
rect 14372 8576 14424 8585
rect 14648 8576 14700 8628
rect 17040 8619 17092 8628
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 18144 8576 18196 8628
rect 20720 8576 20772 8628
rect 22192 8576 22244 8628
rect 23296 8576 23348 8628
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 24768 8576 24820 8628
rect 21916 8551 21968 8560
rect 21916 8517 21925 8551
rect 21925 8517 21959 8551
rect 21959 8517 21968 8551
rect 21916 8508 21968 8517
rect 22284 8508 22336 8560
rect 14924 8483 14976 8492
rect 12532 8372 12584 8424
rect 14096 8372 14148 8424
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 17868 8440 17920 8492
rect 18788 8440 18840 8492
rect 18328 8372 18380 8424
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 20260 8415 20312 8424
rect 20260 8381 20294 8415
rect 20294 8381 20312 8415
rect 15844 8304 15896 8356
rect 17960 8304 18012 8356
rect 18696 8304 18748 8356
rect 19340 8304 19392 8356
rect 20260 8372 20312 8381
rect 22468 8415 22520 8424
rect 22468 8381 22477 8415
rect 22477 8381 22511 8415
rect 22511 8381 22520 8415
rect 22468 8372 22520 8381
rect 24032 8415 24084 8424
rect 24032 8381 24041 8415
rect 24041 8381 24075 8415
rect 24075 8381 24084 8415
rect 24032 8372 24084 8381
rect 24860 8372 24912 8424
rect 20076 8304 20128 8356
rect 20536 8304 20588 8356
rect 21732 8304 21784 8356
rect 24584 8304 24636 8356
rect 25504 8304 25556 8356
rect 16212 8236 16264 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 11980 8007 12032 8016
rect 11980 7973 11989 8007
rect 11989 7973 12023 8007
rect 12023 7973 12032 8007
rect 11980 7964 12032 7973
rect 12440 8007 12492 8016
rect 12440 7973 12449 8007
rect 12449 7973 12483 8007
rect 12483 7973 12492 8007
rect 13728 8032 13780 8084
rect 14188 8032 14240 8084
rect 14924 8075 14976 8084
rect 14924 8041 14933 8075
rect 14933 8041 14967 8075
rect 14967 8041 14976 8075
rect 14924 8032 14976 8041
rect 16488 8032 16540 8084
rect 17684 8032 17736 8084
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 21088 8075 21140 8084
rect 21088 8041 21097 8075
rect 21097 8041 21131 8075
rect 21131 8041 21140 8075
rect 21088 8032 21140 8041
rect 24584 8075 24636 8084
rect 24584 8041 24593 8075
rect 24593 8041 24627 8075
rect 24627 8041 24636 8075
rect 24584 8032 24636 8041
rect 24860 8032 24912 8084
rect 12440 7964 12492 7973
rect 14648 7964 14700 8016
rect 15844 8007 15896 8016
rect 15844 7973 15853 8007
rect 15853 7973 15887 8007
rect 15887 7973 15896 8007
rect 15844 7964 15896 7973
rect 16304 7964 16356 8016
rect 14004 7896 14056 7948
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12808 7828 12860 7880
rect 14832 7828 14884 7880
rect 17132 7828 17184 7880
rect 18512 7939 18564 7948
rect 18512 7905 18521 7939
rect 18521 7905 18555 7939
rect 18555 7905 18564 7939
rect 18512 7896 18564 7905
rect 20904 7896 20956 7948
rect 23388 7964 23440 8016
rect 22928 7939 22980 7948
rect 22928 7905 22962 7939
rect 22962 7905 22980 7939
rect 22928 7896 22980 7905
rect 17868 7828 17920 7880
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 19708 7871 19760 7880
rect 16212 7760 16264 7812
rect 16580 7803 16632 7812
rect 16580 7769 16589 7803
rect 16589 7769 16623 7803
rect 16623 7769 16632 7803
rect 16580 7760 16632 7769
rect 17776 7760 17828 7812
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 22100 7760 22152 7812
rect 22468 7803 22520 7812
rect 22468 7769 22477 7803
rect 22477 7769 22511 7803
rect 22511 7769 22520 7803
rect 22468 7760 22520 7769
rect 12624 7692 12676 7744
rect 19340 7692 19392 7744
rect 20628 7692 20680 7744
rect 22192 7735 22244 7744
rect 22192 7701 22201 7735
rect 22201 7701 22235 7735
rect 22235 7701 22244 7735
rect 22192 7692 22244 7701
rect 22652 7692 22704 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 12440 7488 12492 7540
rect 13360 7488 13412 7540
rect 13544 7488 13596 7540
rect 14832 7488 14884 7540
rect 16948 7488 17000 7540
rect 17500 7488 17552 7540
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 18512 7531 18564 7540
rect 18512 7497 18521 7531
rect 18521 7497 18555 7531
rect 18555 7497 18564 7531
rect 18512 7488 18564 7497
rect 18604 7488 18656 7540
rect 18788 7488 18840 7540
rect 12808 7420 12860 7472
rect 13912 7420 13964 7472
rect 14464 7420 14516 7472
rect 15200 7420 15252 7472
rect 20076 7488 20128 7540
rect 21456 7488 21508 7540
rect 22652 7488 22704 7540
rect 22744 7488 22796 7540
rect 23388 7488 23440 7540
rect 22376 7420 22428 7472
rect 12624 7352 12676 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15844 7352 15896 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 22192 7352 22244 7404
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 24124 7352 24176 7404
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 13636 7284 13688 7336
rect 13820 7284 13872 7336
rect 14280 7284 14332 7336
rect 12808 7259 12860 7268
rect 12808 7225 12817 7259
rect 12817 7225 12851 7259
rect 12851 7225 12860 7259
rect 12808 7216 12860 7225
rect 15660 7284 15712 7336
rect 22376 7327 22428 7336
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 19340 7216 19392 7268
rect 13360 7148 13412 7200
rect 13912 7148 13964 7200
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 16396 7191 16448 7200
rect 16396 7157 16405 7191
rect 16405 7157 16439 7191
rect 16439 7157 16448 7191
rect 16396 7148 16448 7157
rect 16488 7191 16540 7200
rect 16488 7157 16497 7191
rect 16497 7157 16531 7191
rect 16531 7157 16540 7191
rect 16488 7148 16540 7157
rect 17224 7148 17276 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 21548 7148 21600 7200
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 24676 7148 24728 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 12624 6944 12676 6996
rect 12900 6987 12952 6996
rect 12900 6953 12909 6987
rect 12909 6953 12943 6987
rect 12943 6953 12952 6987
rect 12900 6944 12952 6953
rect 14648 6987 14700 6996
rect 14648 6953 14657 6987
rect 14657 6953 14691 6987
rect 14691 6953 14700 6987
rect 14648 6944 14700 6953
rect 15568 6944 15620 6996
rect 16212 6944 16264 6996
rect 16304 6944 16356 6996
rect 18052 6944 18104 6996
rect 18972 6944 19024 6996
rect 12532 6876 12584 6928
rect 13636 6919 13688 6928
rect 13636 6885 13645 6919
rect 13645 6885 13679 6919
rect 13679 6885 13688 6919
rect 13636 6876 13688 6885
rect 16396 6876 16448 6928
rect 17684 6876 17736 6928
rect 20352 6876 20404 6928
rect 21640 6876 21692 6928
rect 22008 6876 22060 6928
rect 22100 6876 22152 6928
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 18880 6808 18932 6860
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 15936 6783 15988 6792
rect 13820 6740 13872 6749
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 22284 6851 22336 6860
rect 22284 6817 22293 6851
rect 22293 6817 22327 6851
rect 22327 6817 22336 6851
rect 22284 6808 22336 6817
rect 14188 6672 14240 6724
rect 18512 6715 18564 6724
rect 18512 6681 18521 6715
rect 18521 6681 18555 6715
rect 18555 6681 18564 6715
rect 18512 6672 18564 6681
rect 18604 6672 18656 6724
rect 21732 6740 21784 6792
rect 22100 6740 22152 6792
rect 22928 6944 22980 6996
rect 24124 6987 24176 6996
rect 24124 6953 24133 6987
rect 24133 6953 24167 6987
rect 24167 6953 24176 6987
rect 24124 6944 24176 6953
rect 23112 6876 23164 6928
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 25228 6851 25280 6860
rect 22744 6808 22796 6817
rect 25228 6817 25237 6851
rect 25237 6817 25271 6851
rect 25271 6817 25280 6851
rect 25228 6808 25280 6817
rect 20812 6672 20864 6724
rect 21916 6672 21968 6724
rect 12900 6604 12952 6656
rect 14556 6604 14608 6656
rect 15936 6604 15988 6656
rect 17132 6604 17184 6656
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 19708 6647 19760 6656
rect 19708 6613 19717 6647
rect 19717 6613 19751 6647
rect 19751 6613 19760 6647
rect 19708 6604 19760 6613
rect 20904 6604 20956 6656
rect 25412 6647 25464 6656
rect 25412 6613 25421 6647
rect 25421 6613 25455 6647
rect 25455 6613 25464 6647
rect 25412 6604 25464 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 14096 6400 14148 6452
rect 13544 6332 13596 6384
rect 11336 6128 11388 6180
rect 13820 6264 13872 6316
rect 15752 6400 15804 6452
rect 18880 6400 18932 6452
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 21732 6400 21784 6452
rect 22744 6443 22796 6452
rect 22744 6409 22753 6443
rect 22753 6409 22787 6443
rect 22787 6409 22796 6443
rect 22744 6400 22796 6409
rect 24032 6443 24084 6452
rect 24032 6409 24041 6443
rect 24041 6409 24075 6443
rect 24075 6409 24084 6443
rect 24032 6400 24084 6409
rect 25228 6443 25280 6452
rect 25228 6409 25237 6443
rect 25237 6409 25271 6443
rect 25271 6409 25280 6443
rect 25228 6400 25280 6409
rect 17592 6264 17644 6316
rect 19064 6264 19116 6316
rect 21640 6375 21692 6384
rect 21640 6341 21649 6375
rect 21649 6341 21683 6375
rect 21683 6341 21692 6375
rect 21640 6332 21692 6341
rect 24492 6332 24544 6384
rect 24676 6264 24728 6316
rect 16948 6196 17000 6248
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 19708 6196 19760 6248
rect 22284 6196 22336 6248
rect 13728 6128 13780 6180
rect 16396 6128 16448 6180
rect 25136 6128 25188 6180
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12532 6060 12584 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 15568 6060 15620 6112
rect 16212 6060 16264 6112
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 17684 6060 17736 6112
rect 17960 6060 18012 6112
rect 18144 6060 18196 6112
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 20996 6103 21048 6112
rect 20996 6069 21005 6103
rect 21005 6069 21039 6103
rect 21039 6069 21048 6103
rect 20996 6060 21048 6069
rect 22652 6060 22704 6112
rect 23572 6060 23624 6112
rect 24492 6060 24544 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 17408 5856 17460 5908
rect 18604 5856 18656 5908
rect 18972 5899 19024 5908
rect 18972 5865 18981 5899
rect 18981 5865 19015 5899
rect 19015 5865 19024 5899
rect 18972 5856 19024 5865
rect 19064 5856 19116 5908
rect 20996 5856 21048 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 22100 5856 22152 5908
rect 25136 5899 25188 5908
rect 25136 5865 25145 5899
rect 25145 5865 25179 5899
rect 25179 5865 25188 5899
rect 25136 5856 25188 5865
rect 12900 5788 12952 5840
rect 15660 5831 15712 5840
rect 15660 5797 15669 5831
rect 15669 5797 15703 5831
rect 15703 5797 15712 5831
rect 15660 5788 15712 5797
rect 17592 5788 17644 5840
rect 21272 5831 21324 5840
rect 21272 5797 21281 5831
rect 21281 5797 21315 5831
rect 21315 5797 21324 5831
rect 21272 5788 21324 5797
rect 12256 5720 12308 5772
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 16028 5720 16080 5772
rect 16396 5720 16448 5772
rect 16948 5720 17000 5772
rect 19524 5720 19576 5772
rect 20260 5720 20312 5772
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 22008 5720 22060 5772
rect 22560 5720 22612 5772
rect 23020 5720 23072 5772
rect 24860 5720 24912 5772
rect 20812 5584 20864 5636
rect 23296 5652 23348 5704
rect 22468 5584 22520 5636
rect 24676 5652 24728 5704
rect 12532 5516 12584 5568
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 17316 5516 17368 5568
rect 20352 5559 20404 5568
rect 20352 5525 20361 5559
rect 20361 5525 20395 5559
rect 20395 5525 20404 5559
rect 20352 5516 20404 5525
rect 20720 5516 20772 5568
rect 22928 5516 22980 5568
rect 23112 5559 23164 5568
rect 23112 5525 23121 5559
rect 23121 5525 23155 5559
rect 23155 5525 23164 5559
rect 23112 5516 23164 5525
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 24676 5559 24728 5568
rect 23480 5516 23532 5525
rect 24676 5525 24685 5559
rect 24685 5525 24719 5559
rect 24719 5525 24728 5559
rect 24676 5516 24728 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 15660 5312 15712 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 19984 5312 20036 5364
rect 20812 5312 20864 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 21824 5312 21876 5364
rect 23020 5355 23072 5364
rect 23020 5321 23029 5355
rect 23029 5321 23063 5355
rect 23063 5321 23072 5355
rect 23020 5312 23072 5321
rect 23112 5312 23164 5364
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 22744 5244 22796 5296
rect 24860 5312 24912 5364
rect 13636 5176 13688 5228
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 20352 5176 20404 5228
rect 20536 5219 20588 5228
rect 20536 5185 20545 5219
rect 20545 5185 20579 5219
rect 20579 5185 20588 5219
rect 20536 5176 20588 5185
rect 22468 5219 22520 5228
rect 22468 5185 22477 5219
rect 22477 5185 22511 5219
rect 22511 5185 22520 5219
rect 22468 5176 22520 5185
rect 23112 5176 23164 5228
rect 13176 5108 13228 5160
rect 14096 5108 14148 5160
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 19340 5108 19392 5160
rect 19984 5108 20036 5160
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23572 5108 23624 5160
rect 15108 5040 15160 5092
rect 19524 5040 19576 5092
rect 12164 5015 12216 5024
rect 12164 4981 12173 5015
rect 12173 4981 12207 5015
rect 12207 4981 12216 5015
rect 12164 4972 12216 4981
rect 12348 4972 12400 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 24676 5040 24728 5092
rect 24768 4972 24820 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 13176 4768 13228 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 15384 4768 15436 4820
rect 15936 4768 15988 4820
rect 16488 4768 16540 4820
rect 17316 4768 17368 4820
rect 17868 4768 17920 4820
rect 18328 4768 18380 4820
rect 18972 4768 19024 4820
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 21272 4768 21324 4820
rect 23480 4768 23532 4820
rect 12256 4700 12308 4752
rect 16396 4700 16448 4752
rect 17132 4743 17184 4752
rect 17132 4709 17141 4743
rect 17141 4709 17175 4743
rect 17175 4709 17184 4743
rect 17132 4700 17184 4709
rect 20352 4700 20404 4752
rect 20536 4700 20588 4752
rect 20996 4700 21048 4752
rect 12532 4675 12584 4684
rect 12532 4641 12566 4675
rect 12566 4641 12584 4675
rect 12532 4632 12584 4641
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 13176 4428 13228 4480
rect 13452 4428 13504 4480
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 14832 4428 14884 4480
rect 17592 4632 17644 4684
rect 19984 4632 20036 4684
rect 17408 4564 17460 4616
rect 19892 4607 19944 4616
rect 19892 4573 19901 4607
rect 19901 4573 19935 4607
rect 19935 4573 19944 4607
rect 19892 4564 19944 4573
rect 20812 4564 20864 4616
rect 20444 4496 20496 4548
rect 17132 4428 17184 4480
rect 17592 4428 17644 4480
rect 22284 4471 22336 4480
rect 22284 4437 22293 4471
rect 22293 4437 22327 4471
rect 22327 4437 22336 4471
rect 22284 4428 22336 4437
rect 22744 4428 22796 4480
rect 24768 4471 24820 4480
rect 24768 4437 24777 4471
rect 24777 4437 24811 4471
rect 24811 4437 24820 4471
rect 24768 4428 24820 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 12532 4224 12584 4276
rect 17408 4224 17460 4276
rect 14740 4156 14792 4208
rect 19892 4224 19944 4276
rect 20996 4267 21048 4276
rect 20996 4233 21005 4267
rect 21005 4233 21039 4267
rect 21039 4233 21048 4267
rect 20996 4224 21048 4233
rect 21456 4224 21508 4276
rect 22744 4224 22796 4276
rect 7748 4088 7800 4140
rect 8208 4088 8260 4140
rect 12532 4088 12584 4140
rect 12992 4088 13044 4140
rect 12348 4020 12400 4072
rect 13452 4020 13504 4072
rect 13636 4063 13688 4072
rect 13636 4029 13670 4063
rect 13670 4029 13688 4063
rect 13636 4020 13688 4029
rect 16396 4020 16448 4072
rect 16948 4088 17000 4140
rect 17776 4088 17828 4140
rect 18328 4088 18380 4140
rect 18880 4088 18932 4140
rect 24676 4224 24728 4276
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 12256 3884 12308 3936
rect 13452 3884 13504 3936
rect 14096 3884 14148 3936
rect 14832 3884 14884 3936
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 20812 4020 20864 4072
rect 18972 3952 19024 4004
rect 20076 3952 20128 4004
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 22744 3952 22796 4004
rect 23848 3952 23900 4004
rect 18328 3884 18380 3936
rect 22284 3927 22336 3936
rect 22284 3893 22293 3927
rect 22293 3893 22327 3927
rect 22327 3893 22336 3927
rect 22284 3884 22336 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 11704 3723 11756 3732
rect 11704 3689 11713 3723
rect 11713 3689 11747 3723
rect 11747 3689 11756 3723
rect 11704 3680 11756 3689
rect 13636 3680 13688 3732
rect 14188 3680 14240 3732
rect 14556 3680 14608 3732
rect 14832 3680 14884 3732
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 15108 3680 15160 3689
rect 19432 3680 19484 3732
rect 19984 3680 20036 3732
rect 20444 3680 20496 3732
rect 21364 3723 21416 3732
rect 21364 3689 21373 3723
rect 21373 3689 21407 3723
rect 21407 3689 21416 3723
rect 21364 3680 21416 3689
rect 22376 3680 22428 3732
rect 22560 3723 22612 3732
rect 22560 3689 22569 3723
rect 22569 3689 22603 3723
rect 22603 3689 22612 3723
rect 22560 3680 22612 3689
rect 23296 3723 23348 3732
rect 23296 3689 23305 3723
rect 23305 3689 23339 3723
rect 23339 3689 23348 3723
rect 23296 3680 23348 3689
rect 23756 3723 23808 3732
rect 23756 3689 23765 3723
rect 23765 3689 23799 3723
rect 23799 3689 23808 3723
rect 23756 3680 23808 3689
rect 24860 3723 24912 3732
rect 24860 3689 24869 3723
rect 24869 3689 24903 3723
rect 24903 3689 24912 3723
rect 24860 3680 24912 3689
rect 25228 3723 25280 3732
rect 25228 3689 25237 3723
rect 25237 3689 25271 3723
rect 25271 3689 25280 3723
rect 25228 3680 25280 3689
rect 25320 3723 25372 3732
rect 25320 3689 25329 3723
rect 25329 3689 25363 3723
rect 25363 3689 25372 3723
rect 25320 3680 25372 3689
rect 14096 3612 14148 3664
rect 16948 3612 17000 3664
rect 10784 3544 10836 3596
rect 12256 3544 12308 3596
rect 12716 3544 12768 3596
rect 15384 3587 15436 3596
rect 15384 3553 15393 3587
rect 15393 3553 15427 3587
rect 15427 3553 15436 3587
rect 15384 3544 15436 3553
rect 15660 3544 15712 3596
rect 20076 3655 20128 3664
rect 20076 3621 20085 3655
rect 20085 3621 20119 3655
rect 20119 3621 20128 3655
rect 20076 3612 20128 3621
rect 23204 3612 23256 3664
rect 19984 3544 20036 3596
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 13084 3476 13136 3528
rect 13912 3476 13964 3528
rect 14832 3476 14884 3528
rect 16396 3476 16448 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 18144 3408 18196 3460
rect 18880 3451 18932 3460
rect 18880 3417 18889 3451
rect 18889 3417 18923 3451
rect 18923 3417 18932 3451
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 25504 3519 25556 3528
rect 18880 3408 18932 3417
rect 23848 3408 23900 3460
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 24768 3408 24820 3460
rect 10692 3383 10744 3392
rect 10692 3349 10701 3383
rect 10701 3349 10735 3383
rect 10735 3349 10744 3383
rect 10692 3340 10744 3349
rect 13544 3340 13596 3392
rect 13728 3340 13780 3392
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 16672 3340 16724 3392
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 18972 3383 19024 3392
rect 18972 3349 18981 3383
rect 18981 3349 19015 3383
rect 19015 3349 19024 3383
rect 18972 3340 19024 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 12256 3179 12308 3188
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 12716 3136 12768 3188
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 13912 3136 13964 3188
rect 14096 3111 14148 3120
rect 11152 2932 11204 2984
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 16948 3136 17000 3188
rect 17316 3179 17368 3188
rect 17316 3145 17325 3179
rect 17325 3145 17359 3179
rect 17359 3145 17368 3179
rect 17316 3136 17368 3145
rect 20076 3136 20128 3188
rect 14096 3068 14148 3077
rect 16764 3068 16816 3120
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 14556 3043 14608 3052
rect 12440 3000 12492 3009
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 21272 3136 21324 3188
rect 23204 3136 23256 3188
rect 21088 3068 21140 3120
rect 21456 3068 21508 3120
rect 23756 3136 23808 3188
rect 25320 3136 25372 3188
rect 25504 3136 25556 3188
rect 13360 2932 13412 2984
rect 14832 2975 14884 2984
rect 14832 2941 14866 2975
rect 14866 2941 14884 2975
rect 14832 2932 14884 2941
rect 18328 2975 18380 2984
rect 16396 2864 16448 2916
rect 17592 2864 17644 2916
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 18420 2932 18472 2984
rect 21180 2975 21232 2984
rect 21180 2941 21189 2975
rect 21189 2941 21223 2975
rect 21223 2941 21232 2975
rect 21180 2932 21232 2941
rect 22560 2932 22612 2984
rect 25228 3000 25280 3052
rect 21088 2864 21140 2916
rect 21272 2907 21324 2916
rect 21272 2873 21281 2907
rect 21281 2873 21315 2907
rect 21315 2873 21324 2907
rect 21272 2864 21324 2873
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 13636 2839 13688 2848
rect 13636 2805 13645 2839
rect 13645 2805 13679 2839
rect 13679 2805 13688 2839
rect 13636 2796 13688 2805
rect 14372 2796 14424 2848
rect 15476 2796 15528 2848
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 16948 2796 17000 2805
rect 23204 2796 23256 2848
rect 24768 2839 24820 2848
rect 24768 2805 24777 2839
rect 24777 2805 24811 2839
rect 24811 2805 24820 2839
rect 24768 2796 24820 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 6000 2592 6052 2644
rect 8392 2592 8444 2644
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 14832 2592 14884 2644
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 16948 2592 17000 2644
rect 18144 2635 18196 2644
rect 12440 2567 12492 2576
rect 12440 2533 12449 2567
rect 12449 2533 12483 2567
rect 12483 2533 12492 2567
rect 12440 2524 12492 2533
rect 2964 2456 3016 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 8392 2456 8444 2508
rect 10692 2456 10744 2508
rect 11520 2456 11572 2508
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19984 2592 20036 2644
rect 21180 2592 21232 2644
rect 21364 2635 21416 2644
rect 21364 2601 21373 2635
rect 21373 2601 21407 2635
rect 21407 2601 21416 2635
rect 21364 2592 21416 2601
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 14372 2456 14424 2508
rect 15936 2456 15988 2508
rect 16120 2456 16172 2508
rect 16396 2431 16448 2440
rect 16396 2397 16405 2431
rect 16405 2397 16439 2431
rect 16439 2397 16448 2431
rect 16396 2388 16448 2397
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 4068 2320 4120 2372
rect 15384 2320 15436 2372
rect 8392 2252 8444 2304
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 18328 2363 18380 2372
rect 18328 2329 18337 2363
rect 18337 2329 18371 2363
rect 18371 2329 18380 2363
rect 18328 2320 18380 2329
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 20168 2456 20220 2508
rect 21732 2499 21784 2508
rect 21732 2465 21741 2499
rect 21741 2465 21775 2499
rect 21775 2465 21784 2499
rect 21732 2456 21784 2465
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 23940 2456 23992 2508
rect 18972 2320 19024 2372
rect 24676 2320 24728 2372
rect 26148 2320 26200 2372
rect 17224 2252 17276 2304
rect 18788 2252 18840 2304
rect 19340 2295 19392 2304
rect 19340 2261 19349 2295
rect 19349 2261 19383 2295
rect 19383 2261 19392 2295
rect 19340 2252 19392 2261
rect 20076 2295 20128 2304
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 21916 2295 21968 2304
rect 21916 2261 21925 2295
rect 21925 2261 21959 2295
rect 21959 2261 21968 2295
rect 21916 2252 21968 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 13912 552 13964 604
rect 14372 552 14424 604
rect 17132 552 17184 604
rect 17316 552 17368 604
rect 22928 552 22980 604
rect 23480 552 23532 604
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2318 27520 2374 28000
rect 2962 27520 3018 28000
rect 3698 27520 3754 28000
rect 4342 27520 4398 28000
rect 4986 27520 5042 28000
rect 5722 27520 5778 28000
rect 6366 27520 6422 28000
rect 7102 27520 7158 28000
rect 7746 27520 7802 28000
rect 8390 27520 8446 28000
rect 9126 27520 9182 28000
rect 9770 27520 9826 28000
rect 10506 27520 10562 28000
rect 11150 27520 11206 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13174 27520 13230 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15290 27520 15346 28000
rect 15934 27520 15990 28000
rect 16578 27520 16634 28000
rect 17314 27520 17370 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19338 27520 19394 28000
rect 20074 27520 20130 28000
rect 20718 27520 20774 28000
rect 21362 27520 21418 28000
rect 22098 27520 22154 28000
rect 22742 27520 22798 28000
rect 23294 27704 23350 27713
rect 23294 27639 23350 27648
rect 308 27418 336 27520
rect 308 27390 428 27418
rect 400 16289 428 27390
rect 952 22658 980 27520
rect 1596 24721 1624 27520
rect 1582 24712 1638 24721
rect 1582 24647 1638 24656
rect 1490 22672 1546 22681
rect 952 22630 1490 22658
rect 1490 22607 1546 22616
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 1582 20904 1638 20913
rect 1582 20839 1584 20848
rect 1636 20839 1638 20848
rect 1584 20810 1636 20816
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1582 20360 1638 20369
rect 1412 19718 1440 20334
rect 1582 20295 1638 20304
rect 1596 20262 1624 20295
rect 1964 20262 1992 20946
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 386 16280 442 16289
rect 386 16215 442 16224
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 294 3360 350 3369
rect 294 3295 350 3304
rect 308 480 336 3295
rect 952 480 980 3431
rect 1412 3346 1440 19654
rect 1674 13968 1730 13977
rect 1674 13903 1730 13912
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10606 1532 10950
rect 1688 10606 1716 13903
rect 1492 10600 1544 10606
rect 1490 10568 1492 10577
rect 1676 10600 1728 10606
rect 1544 10568 1546 10577
rect 1676 10542 1728 10548
rect 1490 10503 1546 10512
rect 1688 10266 1716 10542
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1964 3505 1992 20198
rect 2332 13161 2360 27520
rect 2976 24313 3004 27520
rect 2962 24304 3018 24313
rect 2962 24239 3018 24248
rect 3712 22409 3740 27520
rect 4356 24585 4384 27520
rect 4342 24576 4398 24585
rect 4342 24511 4398 24520
rect 5000 23633 5028 27520
rect 5736 25242 5764 27520
rect 5552 25214 5764 25242
rect 4986 23624 5042 23633
rect 4986 23559 5042 23568
rect 3698 22400 3754 22409
rect 3698 22335 3754 22344
rect 5552 22001 5580 25214
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5538 21992 5594 22001
rect 5538 21927 5594 21936
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6380 21457 6408 27520
rect 6366 21448 6422 21457
rect 6366 21383 6422 21392
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 7116 19281 7144 27520
rect 7760 19961 7788 27520
rect 8404 23526 8432 27520
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 9140 20777 9168 27520
rect 9784 24177 9812 27520
rect 10520 27418 10548 27520
rect 10520 27390 10732 27418
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10138 24576 10194 24585
rect 10138 24511 10194 24520
rect 10152 24342 10180 24511
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10140 24336 10192 24342
rect 10140 24278 10192 24284
rect 9770 24168 9826 24177
rect 9770 24103 9826 24112
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9126 20768 9182 20777
rect 9126 20703 9182 20712
rect 7746 19952 7802 19961
rect 7746 19887 7802 19896
rect 9600 19292 9628 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 23338 10732 27390
rect 10704 23310 10824 23338
rect 10796 23225 10824 23310
rect 10782 23216 10838 23225
rect 10782 23151 10838 23160
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10612 22642 10640 23054
rect 10888 22778 10916 23122
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10598 21992 10654 22001
rect 10598 21927 10654 21936
rect 10612 21690 10640 21927
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 11058 21448 11114 21457
rect 11058 21383 11114 21392
rect 11072 21350 11100 21383
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 20505 10824 21286
rect 11072 20806 11100 21286
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10782 20496 10838 20505
rect 10782 20431 10838 20440
rect 10968 20256 11020 20262
rect 10966 20224 10968 20233
rect 11020 20224 11022 20233
rect 10289 20156 10585 20176
rect 10966 20159 11022 20168
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 9876 19446 9904 19858
rect 10336 19514 10364 19858
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 9864 19440 9916 19446
rect 11164 19417 11192 27520
rect 11794 24304 11850 24313
rect 11794 24239 11850 24248
rect 11808 24206 11836 24239
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23662 11376 24006
rect 11426 23896 11482 23905
rect 11808 23866 11836 24142
rect 11426 23831 11428 23840
rect 11480 23831 11482 23840
rect 11796 23860 11848 23866
rect 11428 23802 11480 23808
rect 11796 23802 11848 23808
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11334 23488 11390 23497
rect 11334 23423 11390 23432
rect 11348 21978 11376 23423
rect 11900 23361 11928 27520
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 12084 23633 12112 24210
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12256 23656 12308 23662
rect 12070 23624 12126 23633
rect 12256 23598 12308 23604
rect 12070 23559 12126 23568
rect 12084 23526 12112 23559
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11886 23352 11942 23361
rect 11886 23287 11942 23296
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11348 21950 11560 21978
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11256 19922 11284 21286
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11440 20262 11468 20878
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11348 20058 11376 20198
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11440 19990 11468 20198
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 9864 19382 9916 19388
rect 11150 19408 11206 19417
rect 10968 19372 11020 19378
rect 11150 19343 11206 19352
rect 10968 19314 11020 19320
rect 9680 19304 9732 19310
rect 7102 19272 7158 19281
rect 9600 19264 9680 19292
rect 9680 19246 9732 19252
rect 10874 19272 10930 19281
rect 7102 19207 7158 19216
rect 10874 19207 10930 19216
rect 10888 19174 10916 19207
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 10336 18426 10364 18770
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18426 10640 18702
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10612 18136 10640 18362
rect 10704 18290 10732 19110
rect 10888 18630 10916 19110
rect 10980 18834 11008 19314
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10612 18108 10732 18136
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17746 10732 18108
rect 10888 17898 10916 18566
rect 11440 18290 11468 18566
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 10968 18080 11020 18086
rect 11152 18080 11204 18086
rect 11020 18028 11100 18034
rect 10968 18022 11100 18028
rect 11152 18022 11204 18028
rect 10980 18006 11100 18022
rect 10888 17870 11008 17898
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10876 17672 10928 17678
rect 10874 17640 10876 17649
rect 10928 17640 10930 17649
rect 10874 17575 10930 17584
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 8206 14376 8262 14385
rect 8206 14311 8262 14320
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 2318 13152 2374 13161
rect 2318 13087 2374 13096
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 4986 11112 5042 11121
rect 4986 11047 5042 11056
rect 2870 10568 2926 10577
rect 2870 10503 2926 10512
rect 4342 10568 4398 10577
rect 4342 10503 4398 10512
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 9625 2820 10406
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2884 9353 2912 10503
rect 2870 9344 2926 9353
rect 2870 9279 2926 9288
rect 2318 6352 2374 6361
rect 2318 6287 2374 6296
rect 1950 3496 2006 3505
rect 1950 3431 2006 3440
rect 1412 3318 1624 3346
rect 1596 480 1624 3318
rect 2332 480 2360 6287
rect 2884 4729 2912 9279
rect 3698 6760 3754 6769
rect 3698 6695 3754 6704
rect 2870 4720 2926 4729
rect 2870 4655 2926 4664
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2976 480 3004 2450
rect 3712 480 3740 6695
rect 4066 2408 4122 2417
rect 4066 2343 4068 2352
rect 4120 2343 4122 2352
rect 4068 2314 4120 2320
rect 4356 480 4384 10503
rect 5000 480 5028 11047
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6366 7440 6422 7449
rect 6366 7375 6422 7384
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5998 5536 6054 5545
rect 5622 5468 5918 5488
rect 5998 5471 6054 5480
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2650 6040 5471
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5552 1578 5580 2450
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5552 1550 5764 1578
rect 5736 480 5764 1550
rect 6380 480 6408 7375
rect 8220 4146 8248 14311
rect 10980 14113 11008 17870
rect 11072 17082 11100 18006
rect 11164 17649 11192 18022
rect 11440 17814 11468 18226
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11150 17640 11206 17649
rect 11150 17575 11206 17584
rect 11440 17202 11468 17750
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11072 17054 11192 17082
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16726 11100 16934
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16250 11100 16662
rect 11164 16590 11192 17054
rect 11256 16794 11284 17138
rect 11426 17096 11482 17105
rect 11336 17060 11388 17066
rect 11426 17031 11482 17040
rect 11336 17002 11388 17008
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11348 16658 11376 17002
rect 11440 16998 11468 17031
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11348 16114 11376 16594
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 10966 14104 11022 14113
rect 10966 14039 11022 14048
rect 11058 13696 11114 13705
rect 10289 13628 10585 13648
rect 11058 13631 11114 13640
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 8390 13288 8446 13297
rect 8390 13223 8446 13232
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 7116 480 7144 3975
rect 7760 480 7788 4082
rect 8404 2650 8432 13223
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9954 9616 10010 9625
rect 9954 9551 10010 9560
rect 9968 9518 9996 9551
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9680 9376 9732 9382
rect 9678 9344 9680 9353
rect 9732 9344 9734 9353
rect 9678 9279 9734 9288
rect 9126 9072 9182 9081
rect 9126 9007 9182 9016
rect 9034 6216 9090 6225
rect 9034 6151 9090 6160
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8404 2310 8432 2450
rect 9048 2417 9076 6151
rect 9034 2408 9090 2417
rect 9034 2343 9090 2352
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 480 8432 2246
rect 9140 480 9168 9007
rect 9692 8974 9720 9279
rect 9968 9178 9996 9454
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10888 9042 10916 9318
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 10888 8634 10916 8978
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10874 7712 10930 7721
rect 10874 7647 10930 7656
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 9770 5128 9826 5137
rect 9770 5063 9826 5072
rect 9784 480 9812 5063
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10782 4584 10838 4593
rect 10782 4519 10838 4528
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10796 3602 10824 4519
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2514 10732 3334
rect 10796 3194 10824 3538
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10888 3074 10916 7647
rect 10796 3046 10916 3074
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10520 1465 10548 2246
rect 10506 1456 10562 1465
rect 10506 1391 10562 1400
rect 10796 1034 10824 3046
rect 10520 1006 10824 1034
rect 10520 480 10548 1006
rect 11072 626 11100 13631
rect 11440 12424 11468 16934
rect 11164 12396 11468 12424
rect 11164 10690 11192 12396
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11256 10810 11284 11154
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11164 10662 11284 10690
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11164 9926 11192 10134
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9382 11192 9862
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8634 11192 8910
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11256 8537 11284 10662
rect 11348 10606 11376 10950
rect 11532 10810 11560 21950
rect 11992 21894 12020 22918
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11992 21554 12020 21830
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11992 21078 12020 21490
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11624 19378 11652 19654
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11624 11898 11652 12310
rect 11716 12170 11744 20742
rect 11992 20602 12020 21014
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11900 19922 11928 20198
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11808 17338 11836 17682
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11808 16182 11836 16526
rect 11900 16250 11928 16526
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 12084 13841 12112 23462
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12176 21486 12204 21830
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12070 13832 12126 13841
rect 12070 13767 12126 13776
rect 11886 12472 11942 12481
rect 11886 12407 11942 12416
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11624 10266 11652 10474
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11242 8528 11298 8537
rect 11348 8498 11376 9862
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9382 11836 9522
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11242 8463 11298 8472
rect 11336 8492 11388 8498
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 11164 3194 11192 6831
rect 11256 4049 11284 8463
rect 11336 8434 11388 8440
rect 11808 6361 11836 9318
rect 11794 6352 11850 6361
rect 11794 6287 11850 6296
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5234 11376 6122
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11702 4176 11758 4185
rect 11702 4111 11758 4120
rect 11242 4040 11298 4049
rect 11242 3975 11298 3984
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11164 2990 11192 3130
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11428 2848 11480 2854
rect 11426 2816 11428 2825
rect 11480 2816 11482 2825
rect 11426 2751 11482 2760
rect 11532 2514 11560 3878
rect 11716 3738 11744 4111
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1601 11652 2246
rect 11610 1592 11666 1601
rect 11610 1527 11666 1536
rect 11072 598 11192 626
rect 11164 480 11192 598
rect 11900 480 11928 12407
rect 12268 11354 12296 23598
rect 12360 22114 12388 24006
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 23254 12480 23598
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12452 22642 12480 23190
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12360 22098 12480 22114
rect 12360 22092 12492 22098
rect 12360 22086 12440 22092
rect 12440 22034 12492 22040
rect 12452 22003 12480 22034
rect 12544 21865 12572 27520
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12806 24168 12862 24177
rect 12728 23662 12756 24142
rect 12806 24103 12862 24112
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12530 21856 12586 21865
rect 12530 21791 12586 21800
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12544 20602 12572 21354
rect 12728 21350 12756 21422
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12438 20088 12494 20097
rect 12438 20023 12494 20032
rect 12532 20052 12584 20058
rect 12346 19952 12402 19961
rect 12346 19887 12402 19896
rect 12360 18408 12388 19887
rect 12452 19122 12480 20023
rect 12532 19994 12584 20000
rect 12544 19718 12572 19994
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19310 12572 19654
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12452 19094 12572 19122
rect 12360 18380 12480 18408
rect 12452 18154 12480 18380
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12452 16046 12480 16730
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12544 14770 12572 19094
rect 12636 14958 12664 21286
rect 12728 19174 12756 21286
rect 12820 21185 12848 24103
rect 12912 23497 12940 24686
rect 13188 24154 13216 27520
rect 13358 24848 13414 24857
rect 13358 24783 13414 24792
rect 13372 24614 13400 24783
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13004 24126 13216 24154
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 12898 23488 12954 23497
rect 12898 23423 12954 23432
rect 12806 21176 12862 21185
rect 12806 21111 12862 21120
rect 12898 20496 12954 20505
rect 12898 20431 12900 20440
rect 12952 20431 12954 20440
rect 12900 20402 12952 20408
rect 12806 19408 12862 19417
rect 12806 19343 12862 19352
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12820 18970 12848 19343
rect 12900 19168 12952 19174
rect 12898 19136 12900 19145
rect 12952 19136 12954 19145
rect 12898 19071 12954 19080
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12820 18222 12848 18906
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12808 18080 12860 18086
rect 12806 18048 12808 18057
rect 12860 18048 12862 18057
rect 12806 17983 12862 17992
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17134 12756 17478
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16794 12756 17070
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13004 16561 13032 24126
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13372 23322 13400 24006
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 12990 16552 13046 16561
rect 12990 16487 13046 16496
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12544 14742 12848 14770
rect 12714 13424 12770 13433
rect 12714 13359 12770 13368
rect 12728 12753 12756 13359
rect 12714 12744 12770 12753
rect 12624 12708 12676 12714
rect 12714 12679 12770 12688
rect 12624 12650 12676 12656
rect 12440 12640 12492 12646
rect 12346 12608 12402 12617
rect 12440 12582 12492 12588
rect 12346 12543 12402 12552
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12360 11121 12388 12543
rect 12452 12442 12480 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12452 11898 12480 12378
rect 12636 12238 12664 12650
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12636 11830 12664 12174
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12346 11112 12402 11121
rect 12346 11047 12402 11056
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9654 12020 9862
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11992 9518 12020 9590
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 12084 9110 12112 9998
rect 12360 9438 12480 9466
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12072 9104 12124 9110
rect 12176 9081 12204 9318
rect 12072 9046 12124 9052
rect 12162 9072 12218 9081
rect 12360 9058 12388 9438
rect 12452 9353 12480 9438
rect 12438 9344 12494 9353
rect 12438 9279 12494 9288
rect 12544 9178 12572 10610
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12360 9030 12480 9058
rect 12162 9007 12218 9016
rect 12452 8378 12480 9030
rect 12544 8430 12572 9114
rect 12360 8350 12480 8378
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 11980 8016 12032 8022
rect 11978 7984 11980 7993
rect 12032 7984 12034 7993
rect 11978 7919 12034 7928
rect 12360 7426 12388 8350
rect 12438 8120 12494 8129
rect 12438 8055 12494 8064
rect 12452 8022 12480 8055
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12452 7546 12480 7958
rect 12532 7880 12584 7886
rect 12530 7848 12532 7857
rect 12584 7848 12586 7857
rect 12530 7783 12586 7792
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12438 7440 12494 7449
rect 12360 7398 12438 7426
rect 12438 7375 12494 7384
rect 12544 6934 12572 7783
rect 12636 7750 12664 10542
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12636 7177 12664 7346
rect 12622 7168 12678 7177
rect 12622 7103 12678 7112
rect 12636 7002 12664 7103
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12256 6112 12308 6118
rect 12254 6080 12256 6089
rect 12532 6112 12584 6118
rect 12308 6080 12310 6089
rect 12532 6054 12584 6060
rect 12254 6015 12310 6024
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 5030 12204 5646
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12176 4570 12204 4966
rect 12268 4758 12296 5714
rect 12544 5574 12572 6054
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12256 4616 12308 4622
rect 12176 4564 12256 4570
rect 12176 4558 12308 4564
rect 12176 4542 12296 4558
rect 12268 3942 12296 4542
rect 12360 4078 12388 4966
rect 12544 4690 12572 5510
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12544 4282 12572 4626
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12438 3904 12494 3913
rect 12438 3839 12494 3848
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3505 12296 3538
rect 12254 3496 12310 3505
rect 12254 3431 12310 3440
rect 12268 3194 12296 3431
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12452 3058 12480 3839
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12440 2576 12492 2582
rect 12438 2544 12440 2553
rect 12492 2544 12494 2553
rect 12438 2479 12494 2488
rect 12544 480 12572 4082
rect 12728 3602 12756 12679
rect 12820 9518 12848 14742
rect 13096 14482 13124 22918
rect 13464 22506 13492 23462
rect 13544 23112 13596 23118
rect 13648 23089 13676 24142
rect 13740 23866 13768 24210
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13820 23112 13872 23118
rect 13544 23054 13596 23060
rect 13634 23080 13690 23089
rect 13452 22500 13504 22506
rect 13452 22442 13504 22448
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13372 21146 13400 22034
rect 13464 22030 13492 22442
rect 13556 22234 13584 23054
rect 13820 23054 13872 23060
rect 13634 23015 13690 23024
rect 13832 22778 13860 23054
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13556 22098 13584 22170
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13464 21690 13492 21966
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20466 13216 20742
rect 13266 20496 13322 20505
rect 13176 20460 13228 20466
rect 13266 20431 13322 20440
rect 13176 20402 13228 20408
rect 13188 20262 13216 20402
rect 13280 20330 13308 20431
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13188 19990 13216 20198
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13188 19378 13216 19926
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13556 19514 13584 19858
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13188 18970 13216 19314
rect 13358 19136 13414 19145
rect 13358 19071 13414 19080
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13266 18184 13322 18193
rect 13266 18119 13268 18128
rect 13320 18119 13322 18128
rect 13268 18090 13320 18096
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14482 13216 14758
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13096 14074 13124 14418
rect 13188 14074 13216 14418
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13280 13841 13308 14214
rect 12990 13832 13046 13841
rect 12990 13767 13046 13776
rect 13266 13832 13322 13841
rect 13266 13767 13322 13776
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10470 12940 10950
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 9110 12848 9318
rect 12912 9178 12940 10406
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12912 7834 12940 8978
rect 13004 8378 13032 13767
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13096 9518 13124 12378
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 12102 13216 12242
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11354 13216 12038
rect 13266 11656 13322 11665
rect 13266 11591 13322 11600
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13280 11234 13308 11591
rect 13188 11206 13308 11234
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13188 9042 13216 11206
rect 13372 10441 13400 19071
rect 13740 18970 13768 21286
rect 13832 21146 13860 22102
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13818 20768 13874 20777
rect 13818 20703 13874 20712
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13832 18902 13860 20703
rect 13924 18970 13952 27520
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14016 23526 14044 24142
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 14188 23112 14240 23118
rect 14186 23080 14188 23089
rect 14240 23080 14242 23089
rect 14186 23015 14242 23024
rect 14094 22128 14150 22137
rect 14094 22063 14150 22072
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14016 20058 14044 21490
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14108 19961 14136 22063
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14094 19952 14150 19961
rect 14094 19887 14150 19896
rect 14094 19816 14150 19825
rect 14094 19751 14150 19760
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13820 18760 13872 18766
rect 13740 18708 13820 18714
rect 13740 18702 13872 18708
rect 13740 18686 13860 18702
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13648 17320 13676 18226
rect 13740 17882 13768 18686
rect 13924 18426 13952 18906
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14016 18290 14044 18770
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13820 17332 13872 17338
rect 13648 17292 13820 17320
rect 13820 17274 13872 17280
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13450 16416 13506 16425
rect 13450 16351 13506 16360
rect 13464 10742 13492 16351
rect 13556 12442 13584 16934
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 14385 13676 15914
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15065 13768 15846
rect 13726 15056 13782 15065
rect 13726 14991 13782 15000
rect 13634 14376 13690 14385
rect 13634 14311 13690 14320
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 12889 13860 13670
rect 14016 13569 14044 18226
rect 14108 14634 14136 19751
rect 14200 19174 14228 20198
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14200 18766 14228 19110
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14200 17542 14228 18090
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14200 16114 14228 17478
rect 14292 17241 14320 24686
rect 14384 24682 14412 25298
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14384 21486 14412 24618
rect 14464 24608 14516 24614
rect 14462 24576 14464 24585
rect 14516 24576 14518 24585
rect 14462 24511 14518 24520
rect 14568 23905 14596 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24857 15332 27520
rect 15948 25498 15976 27520
rect 15936 25492 15988 25498
rect 15936 25434 15988 25440
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16408 24886 16436 25094
rect 16396 24880 16448 24886
rect 15290 24848 15346 24857
rect 16396 24822 16448 24828
rect 15290 24783 15346 24792
rect 15198 24712 15254 24721
rect 15198 24647 15200 24656
rect 15252 24647 15254 24656
rect 15200 24618 15252 24624
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15396 24410 15424 24550
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15764 24342 15792 24550
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15752 24336 15804 24342
rect 15752 24278 15804 24284
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14554 23896 14610 23905
rect 14956 23888 15252 23908
rect 14554 23831 14610 23840
rect 14462 23624 14518 23633
rect 14462 23559 14518 23568
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14384 20097 14412 20198
rect 14370 20088 14426 20097
rect 14370 20023 14426 20032
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14384 17542 14412 18158
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14278 17232 14334 17241
rect 14278 17167 14334 17176
rect 14292 16998 14320 17167
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14384 16697 14412 16730
rect 14370 16688 14426 16697
rect 14280 16652 14332 16658
rect 14370 16623 14426 16632
rect 14280 16594 14332 16600
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14292 15706 14320 16594
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14108 14606 14412 14634
rect 14186 14512 14242 14521
rect 14186 14447 14242 14456
rect 14200 14074 14228 14447
rect 14278 14376 14334 14385
rect 14278 14311 14280 14320
rect 14332 14311 14334 14320
rect 14280 14282 14332 14288
rect 14278 14104 14334 14113
rect 14188 14068 14240 14074
rect 14278 14039 14334 14048
rect 14188 14010 14240 14016
rect 14200 13870 14228 14010
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14002 13560 14058 13569
rect 14002 13495 14058 13504
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 13818 12880 13874 12889
rect 13818 12815 13874 12824
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13740 12186 13768 12310
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13556 10792 13584 11630
rect 13648 11354 13676 12174
rect 13740 12158 13860 12186
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13556 10764 13676 10792
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10577 13584 10610
rect 13542 10568 13598 10577
rect 13542 10503 13598 10512
rect 13544 10464 13596 10470
rect 13358 10432 13414 10441
rect 13544 10406 13596 10412
rect 13358 10367 13414 10376
rect 13372 9353 13400 10367
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13464 9110 13492 9930
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8412 13400 8774
rect 13280 8384 13400 8412
rect 13450 8392 13506 8401
rect 13004 8350 13124 8378
rect 12990 8256 13046 8265
rect 12990 8191 13046 8200
rect 13004 7993 13032 8191
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 12820 7478 12848 7822
rect 12912 7806 13032 7834
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12900 7336 12952 7342
rect 12806 7304 12862 7313
rect 12900 7278 12952 7284
rect 12806 7239 12808 7248
rect 12860 7239 12862 7248
rect 12808 7210 12860 7216
rect 12912 7002 12940 7278
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 5846 12940 6598
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12912 5234 12940 5782
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 13004 4146 13032 7806
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12728 3194 12756 3538
rect 13096 3534 13124 8350
rect 13280 8276 13308 8384
rect 13450 8327 13506 8336
rect 13280 8248 13400 8276
rect 13372 7546 13400 8248
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13372 7206 13400 7375
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13464 6769 13492 8327
rect 13556 7721 13584 10406
rect 13648 10010 13676 10764
rect 13740 10198 13768 11018
rect 13832 10810 13860 12158
rect 14200 12102 14228 13330
rect 14292 12374 14320 14039
rect 14384 13682 14412 14606
rect 14476 14074 14504 23559
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15304 22982 15332 23462
rect 15474 23352 15530 23361
rect 15474 23287 15530 23296
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14660 21690 14688 21966
rect 14648 21684 14700 21690
rect 14568 21644 14648 21672
rect 14568 17814 14596 21644
rect 14648 21626 14700 21632
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14660 18970 14688 19178
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14660 18426 14688 18906
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14556 17808 14608 17814
rect 14608 17756 14688 17762
rect 14556 17750 14688 17756
rect 14568 17734 14688 17750
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 15910 14596 17614
rect 14660 17338 14688 17734
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14660 16250 14688 16458
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15706 14596 15846
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14476 13870 14504 14010
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14384 13654 14504 13682
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14292 11898 14320 12174
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 13910 11520 13966 11529
rect 13910 11455 13966 11464
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13648 9982 13768 10010
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13542 7712 13598 7721
rect 13542 7647 13598 7656
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13450 6760 13506 6769
rect 13450 6695 13506 6704
rect 13556 6474 13584 7482
rect 13648 7342 13676 9862
rect 13740 9586 13768 9982
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13728 9376 13780 9382
rect 13832 9364 13860 10066
rect 13780 9336 13860 9364
rect 13728 9318 13780 9324
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13740 8090 13768 9114
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13832 7342 13860 9336
rect 13924 7478 13952 11455
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14016 10266 14044 11154
rect 14384 11150 14412 12650
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14476 10792 14504 13654
rect 14752 13530 14780 21422
rect 14844 21146 14872 22918
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 15292 22432 15344 22438
rect 15384 22432 15436 22438
rect 15292 22374 15344 22380
rect 15382 22400 15384 22409
rect 15436 22400 15438 22409
rect 14936 22166 14964 22374
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 15304 21894 15332 22374
rect 15382 22335 15438 22344
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21486 15332 21830
rect 15292 21480 15344 21486
rect 15290 21448 15292 21457
rect 15344 21448 15346 21457
rect 15290 21383 15346 21392
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14936 20890 14964 21286
rect 15304 21146 15332 21383
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15488 21049 15516 23287
rect 15474 21040 15530 21049
rect 15474 20975 15530 20984
rect 14844 20862 14964 20890
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14844 19802 14872 20862
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20618 15332 20878
rect 15382 20632 15438 20641
rect 15304 20590 15382 20618
rect 15304 20262 15332 20590
rect 15382 20567 15438 20576
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15488 19922 15516 20334
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 14844 19774 15332 19802
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14830 19408 14886 19417
rect 14830 19343 14886 19352
rect 14844 18737 14872 19343
rect 15304 18834 15332 19774
rect 15488 19446 15516 19858
rect 15580 19802 15608 24278
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 15764 23769 15792 24006
rect 16132 23866 16160 24142
rect 16316 23866 16344 24346
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 15750 23760 15806 23769
rect 15750 23695 15752 23704
rect 15804 23695 15806 23704
rect 15752 23666 15804 23672
rect 15764 23322 15792 23666
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15764 22642 15792 23258
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15856 22778 15884 23122
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15844 22024 15896 22030
rect 15896 21984 15976 22012
rect 15844 21966 15896 21972
rect 15948 21865 15976 21984
rect 15934 21856 15990 21865
rect 15934 21791 15990 21800
rect 15948 21690 15976 21791
rect 15936 21684 15988 21690
rect 15856 21644 15936 21672
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15672 20233 15700 20946
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15658 20224 15714 20233
rect 15658 20159 15714 20168
rect 15580 19774 15700 19802
rect 15566 19680 15622 19689
rect 15566 19615 15622 19624
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 14830 18728 14886 18737
rect 14830 18663 14886 18672
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 18154 14872 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 14844 17066 14872 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 15028 16794 15056 17070
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15396 16726 15424 17478
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14844 15706 14872 16526
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15106 16144 15162 16153
rect 15106 16079 15162 16088
rect 15120 16046 15148 16079
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14844 15162 14872 15438
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14844 14074 14872 14758
rect 15212 14618 15240 14758
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15304 14550 15332 15302
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14830 13968 14886 13977
rect 14830 13903 14886 13912
rect 14844 13870 14872 13903
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14384 10764 14504 10792
rect 14384 10470 14412 10764
rect 14462 10704 14518 10713
rect 14462 10639 14464 10648
rect 14516 10639 14518 10648
rect 14464 10610 14516 10616
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14186 10296 14242 10305
rect 14004 10260 14056 10266
rect 14186 10231 14242 10240
rect 14004 10202 14056 10208
rect 14200 10062 14228 10231
rect 14096 10056 14148 10062
rect 14094 10024 14096 10033
rect 14188 10056 14240 10062
rect 14148 10024 14150 10033
rect 14016 9982 14094 10010
rect 14016 9722 14044 9982
rect 14188 9998 14240 10004
rect 14094 9959 14150 9968
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14016 7993 14044 8978
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14384 8634 14412 8910
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14002 7984 14058 7993
rect 14002 7919 14004 7928
rect 14056 7919 14058 7928
rect 14004 7890 14056 7896
rect 14016 7859 14044 7890
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13648 6769 13676 6870
rect 13820 6792 13872 6798
rect 13634 6760 13690 6769
rect 13820 6734 13872 6740
rect 13634 6695 13690 6704
rect 13464 6446 13584 6474
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5166 13216 6054
rect 13358 5944 13414 5953
rect 13358 5879 13414 5888
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13188 4826 13216 5102
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 13188 480 13216 4422
rect 13372 3194 13400 5879
rect 13464 4486 13492 6446
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13556 5574 13584 6326
rect 13648 6089 13676 6695
rect 13832 6322 13860 6734
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13924 6202 13952 7142
rect 14108 6458 14136 8366
rect 14186 8256 14242 8265
rect 14186 8191 14242 8200
rect 14200 8090 14228 8191
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14568 7562 14596 12310
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 11354 14688 11562
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14660 10674 14688 11290
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14660 9110 14688 9522
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14660 8634 14688 9046
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14384 7534 14596 7562
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 13740 6186 13952 6202
rect 13728 6180 13952 6186
rect 13780 6174 13952 6180
rect 13728 6122 13780 6128
rect 13634 6080 13690 6089
rect 13634 6015 13690 6024
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13648 4826 13676 5170
rect 14108 5166 14136 6394
rect 14200 5914 14228 6666
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13648 4078 13676 4762
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13464 3942 13492 4014
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13648 3738 13676 4014
rect 14108 3942 14136 5102
rect 14096 3936 14148 3942
rect 14148 3896 14228 3924
rect 14096 3878 14148 3884
rect 14200 3738 14228 3896
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14096 3664 14148 3670
rect 14292 3641 14320 7278
rect 14096 3606 14148 3612
rect 14278 3632 14334 3641
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13372 2990 13400 3130
rect 13556 3097 13584 3334
rect 13542 3088 13598 3097
rect 13542 3023 13598 3032
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13634 2952 13690 2961
rect 13634 2887 13690 2896
rect 13648 2854 13676 2887
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13740 2666 13768 3334
rect 13924 3194 13952 3470
rect 13912 3188 13964 3194
rect 13648 2638 13768 2666
rect 13832 3148 13912 3176
rect 13832 2650 13860 3148
rect 13912 3130 13964 3136
rect 14108 3126 14136 3606
rect 14278 3567 14334 3576
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14384 2854 14412 7534
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13820 2644 13872 2650
rect 13648 2417 13676 2638
rect 13820 2586 13872 2592
rect 14384 2514 14412 2790
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 13634 2408 13690 2417
rect 14476 2394 14504 7414
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14568 6662 14596 7346
rect 14660 7002 14688 7958
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14752 4729 14780 12106
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14924 11552 14976 11558
rect 15396 11529 15424 13806
rect 15488 12986 15516 14418
rect 15580 13297 15608 19615
rect 15672 19514 15700 19774
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15764 18902 15792 20742
rect 15856 20505 15884 21644
rect 15936 21626 15988 21632
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16040 20942 16068 21490
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 20602 16068 20878
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15842 20496 15898 20505
rect 15842 20431 15898 20440
rect 16040 19990 16068 20538
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 16040 19514 16068 19926
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15752 18896 15804 18902
rect 16040 18850 16068 19314
rect 15752 18838 15804 18844
rect 15948 18822 16068 18850
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15750 18048 15806 18057
rect 15750 17983 15806 17992
rect 15764 17882 15792 17983
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 15672 17513 15700 17750
rect 15658 17504 15714 17513
rect 15658 17439 15714 17448
rect 15856 16590 15884 18362
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15672 15201 15700 15506
rect 15658 15192 15714 15201
rect 15658 15127 15714 15136
rect 15672 14822 15700 15127
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15566 13288 15622 13297
rect 15566 13223 15622 13232
rect 15476 12980 15528 12986
rect 15528 12940 15608 12968
rect 15476 12922 15528 12928
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12306 15516 12582
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15580 12238 15608 12940
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15580 11898 15608 12174
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 11778 15700 14758
rect 15948 14532 15976 18822
rect 16132 18766 16160 19382
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16040 18426 16068 18702
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 16040 17338 16068 17546
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16026 16552 16082 16561
rect 16026 16487 16082 16496
rect 16040 16250 16068 16487
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15488 11750 15700 11778
rect 15764 14504 15976 14532
rect 14924 11494 14976 11500
rect 15382 11520 15438 11529
rect 14936 11150 14964 11494
rect 15382 11455 15438 11464
rect 15108 11212 15160 11218
rect 15160 11172 15332 11200
rect 15108 11154 15160 11160
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10810 15332 11172
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 9450 14872 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14844 7886 14872 9386
rect 15028 9353 15056 9386
rect 15014 9344 15070 9353
rect 15014 9279 15070 9288
rect 15488 8838 15516 11750
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 9382 15608 9998
rect 15672 9897 15700 10066
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14936 8090 14964 8434
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7546 14872 7822
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15212 6905 15240 7414
rect 15580 7154 15608 9318
rect 15672 7342 15700 9823
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15580 7126 15700 7154
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15198 6896 15254 6905
rect 15198 6831 15254 6840
rect 15290 6760 15346 6769
rect 15290 6695 15346 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 5914 15332 6695
rect 15580 6118 15608 6938
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15672 5846 15700 7126
rect 15764 6866 15792 14504
rect 16040 13870 16068 14554
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15856 8022 15884 8298
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15856 7206 15884 7346
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15764 6458 15792 6802
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 5840 15712 5846
rect 15658 5808 15660 5817
rect 15712 5808 15714 5817
rect 15658 5743 15714 5752
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15672 5370 15700 5743
rect 15764 5409 15792 6394
rect 15750 5400 15806 5409
rect 15660 5364 15712 5370
rect 15750 5335 15806 5344
rect 15660 5306 15712 5312
rect 15856 5273 15884 7142
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15948 6662 15976 6734
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 5710 15976 6598
rect 16040 5778 16068 10406
rect 16132 7018 16160 17206
rect 16224 15722 16252 23598
rect 16408 23254 16436 24822
rect 16592 24585 16620 27520
rect 16948 25356 17000 25362
rect 16948 25298 17000 25304
rect 16960 24614 16988 25298
rect 17328 25226 17356 27520
rect 17972 25498 18000 27520
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17316 25220 17368 25226
rect 17316 25162 17368 25168
rect 17500 24676 17552 24682
rect 17500 24618 17552 24624
rect 16948 24608 17000 24614
rect 16578 24576 16634 24585
rect 16948 24550 17000 24556
rect 16578 24511 16634 24520
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16500 23338 16528 24142
rect 16684 23526 16712 24210
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16500 23322 16620 23338
rect 16500 23316 16632 23322
rect 16500 23310 16580 23316
rect 16580 23258 16632 23264
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16486 23216 16542 23225
rect 16408 22778 16436 23190
rect 16486 23151 16542 23160
rect 16500 22778 16528 23151
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16408 22658 16436 22714
rect 16316 22630 16436 22658
rect 16486 22672 16542 22681
rect 16316 22030 16344 22630
rect 16486 22607 16542 22616
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16316 21690 16344 21966
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16302 20496 16358 20505
rect 16302 20431 16358 20440
rect 16316 16794 16344 20431
rect 16408 17270 16436 22510
rect 16500 22012 16528 22607
rect 16684 22234 16712 23462
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16672 22228 16724 22234
rect 16672 22170 16724 22176
rect 16580 22024 16632 22030
rect 16500 21984 16580 22012
rect 16580 21966 16632 21972
rect 16672 20256 16724 20262
rect 16670 20224 16672 20233
rect 16724 20224 16726 20233
rect 16670 20159 16726 20168
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16684 18970 16712 19246
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16776 18850 16804 22510
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16868 21690 16896 21898
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16684 18822 16804 18850
rect 16592 18358 16620 18770
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16580 18216 16632 18222
rect 16500 18164 16580 18170
rect 16500 18158 16632 18164
rect 16500 18142 16620 18158
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16316 16046 16344 16730
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16224 15694 16344 15722
rect 16210 15600 16266 15609
rect 16210 15535 16266 15544
rect 16224 15502 16252 15535
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 15026 16252 15438
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16224 14550 16252 14962
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16224 14074 16252 14486
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16316 13546 16344 15694
rect 16408 15570 16436 15846
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16500 15450 16528 18142
rect 16408 15422 16528 15450
rect 16408 15162 16436 15422
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16500 15042 16528 15302
rect 16500 15026 16620 15042
rect 16500 15020 16632 15026
rect 16500 15014 16580 15020
rect 16580 14962 16632 14968
rect 16486 13832 16542 13841
rect 16486 13767 16542 13776
rect 16224 13518 16436 13546
rect 16224 13462 16252 13518
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16224 12442 16252 13262
rect 16316 13161 16344 13330
rect 16302 13152 16358 13161
rect 16302 13087 16358 13096
rect 16316 12918 16344 13087
rect 16408 12986 16436 13518
rect 16500 13433 16528 13767
rect 16486 13424 16542 13433
rect 16486 13359 16542 13368
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16316 12481 16344 12854
rect 16408 12617 16436 12922
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16394 12608 16450 12617
rect 16394 12543 16450 12552
rect 16302 12472 16358 12481
rect 16212 12436 16264 12442
rect 16302 12407 16358 12416
rect 16212 12378 16264 12384
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16316 11082 16344 12242
rect 16500 11898 16528 12718
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16592 11762 16620 11834
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16592 11218 16620 11698
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16316 10266 16344 10610
rect 16500 10282 16528 11154
rect 16592 10810 16620 11154
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16684 10713 16712 18822
rect 16868 18426 16896 19654
rect 16960 19174 16988 24550
rect 17038 23896 17094 23905
rect 17038 23831 17040 23840
rect 17092 23831 17094 23840
rect 17040 23802 17092 23808
rect 17038 23488 17094 23497
rect 17038 23423 17094 23432
rect 17052 22778 17080 23423
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17420 23118 17448 23258
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17420 22710 17448 23054
rect 17512 22778 17540 24618
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17408 22704 17460 22710
rect 17408 22646 17460 22652
rect 17512 22574 17540 22714
rect 17500 22568 17552 22574
rect 17314 22536 17370 22545
rect 17500 22510 17552 22516
rect 17314 22471 17370 22480
rect 17328 22098 17356 22471
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 21146 17172 21830
rect 17328 21350 17356 22034
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17420 21690 17448 21966
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17236 19281 17264 21286
rect 17222 19272 17278 19281
rect 17222 19207 17278 19216
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 17144 18358 17172 18702
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17144 17762 17172 18294
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17052 17746 17172 17762
rect 17040 17740 17172 17746
rect 17092 17734 17172 17740
rect 17040 17682 17092 17688
rect 17052 17338 17080 17682
rect 17040 17332 17092 17338
rect 16960 17292 17040 17320
rect 16960 17066 16988 17292
rect 17040 17274 17092 17280
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16960 16658 16988 17002
rect 17132 16720 17184 16726
rect 17052 16680 17132 16708
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16960 16250 16988 16594
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17052 16114 17080 16680
rect 17132 16662 17184 16668
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16960 15586 16988 15982
rect 17052 15706 17080 16050
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16960 15558 17080 15586
rect 17144 15570 17172 16186
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16776 14006 16804 14418
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16776 11694 16804 13194
rect 16868 12986 16896 13670
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16960 12782 16988 13126
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16868 11762 16896 12106
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16776 11150 16804 11494
rect 16868 11354 16896 11698
rect 16960 11354 16988 11698
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16670 10704 16726 10713
rect 16670 10639 16726 10648
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16500 10266 16620 10282
rect 16304 10260 16356 10266
rect 16500 10260 16632 10266
rect 16500 10254 16580 10260
rect 16304 10202 16356 10208
rect 16580 10202 16632 10208
rect 16316 10062 16344 10202
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16316 9722 16344 9998
rect 16592 9722 16620 10202
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16684 9654 16712 10542
rect 16776 10266 16804 10950
rect 17052 10713 17080 15558
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17144 15162 17172 15506
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17144 14482 17172 15098
rect 17236 14929 17264 18022
rect 17222 14920 17278 14929
rect 17222 14855 17278 14864
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17144 12481 17172 13466
rect 17130 12472 17186 12481
rect 17130 12407 17186 12416
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17144 11218 17172 12310
rect 17222 11792 17278 11801
rect 17222 11727 17278 11736
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17144 10810 17172 11154
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17038 10704 17094 10713
rect 17038 10639 17094 10648
rect 17236 10282 17264 11727
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16960 10254 17264 10282
rect 16856 9920 16908 9926
rect 16762 9888 16818 9897
rect 16856 9862 16908 9868
rect 16762 9823 16818 9832
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16776 9586 16804 9823
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16764 9376 16816 9382
rect 16670 9344 16726 9353
rect 16764 9318 16816 9324
rect 16670 9279 16726 9288
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16224 8294 16252 9046
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16592 8786 16620 8842
rect 16684 8838 16712 9279
rect 16500 8758 16620 8786
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 7818 16252 8230
rect 16500 8090 16528 8758
rect 16776 8650 16804 9318
rect 16684 8622 16804 8650
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16132 7002 16252 7018
rect 16316 7002 16344 7958
rect 16578 7848 16634 7857
rect 16578 7783 16580 7792
rect 16632 7783 16634 7792
rect 16580 7754 16632 7760
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16132 6996 16264 7002
rect 16132 6990 16212 6996
rect 16212 6938 16264 6944
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16408 6934 16436 7142
rect 16396 6928 16448 6934
rect 16394 6896 16396 6905
rect 16448 6896 16450 6905
rect 16394 6831 16450 6840
rect 16408 6805 16436 6831
rect 16396 6180 16448 6186
rect 16396 6122 16448 6128
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15106 5264 15162 5273
rect 15106 5199 15162 5208
rect 15842 5264 15898 5273
rect 15842 5199 15898 5208
rect 15120 5098 15148 5199
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4826 15424 4966
rect 15948 4826 15976 5646
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 14738 4720 14794 4729
rect 14738 4655 14794 4664
rect 15382 4720 15438 4729
rect 15382 4655 15438 4664
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14752 4214 14780 4422
rect 14740 4208 14792 4214
rect 14844 4185 14872 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14740 4150 14792 4156
rect 14830 4176 14886 4185
rect 14830 4111 14886 4120
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3738 14872 3878
rect 15106 3768 15162 3777
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14832 3732 14884 3738
rect 15106 3703 15108 3712
rect 14832 3674 14884 3680
rect 15160 3703 15162 3712
rect 15108 3674 15160 3680
rect 14568 3058 14596 3674
rect 14844 3534 14872 3674
rect 15396 3602 15424 4655
rect 15936 3936 15988 3942
rect 15934 3904 15936 3913
rect 16120 3936 16172 3942
rect 15988 3904 15990 3913
rect 16120 3878 16172 3884
rect 15934 3839 15990 3848
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15382 3496 15438 3505
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14844 2990 14872 3470
rect 15382 3431 15438 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14844 2650 14872 2926
rect 15290 2816 15346 2825
rect 15290 2751 15346 2760
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 13634 2343 13690 2352
rect 14384 2366 14504 2394
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13372 1737 13400 2246
rect 13358 1728 13414 1737
rect 13358 1663 13414 1672
rect 14384 610 14412 2366
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 1873 14504 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14462 1864 14518 1873
rect 14462 1799 14518 1808
rect 14554 1456 14610 1465
rect 14554 1391 14610 1400
rect 13912 604 13964 610
rect 13912 546 13964 552
rect 14372 604 14424 610
rect 14372 546 14424 552
rect 13924 480 13952 546
rect 14568 480 14596 1391
rect 15304 480 15332 2751
rect 15396 2378 15424 3431
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15580 3233 15608 3334
rect 15566 3224 15622 3233
rect 15566 3159 15622 3168
rect 15476 2848 15528 2854
rect 15474 2816 15476 2825
rect 15528 2816 15530 2825
rect 15474 2751 15530 2760
rect 15672 2650 15700 3538
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15934 2544 15990 2553
rect 16132 2514 16160 3878
rect 16224 2553 16252 6054
rect 16408 5914 16436 6122
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16302 5672 16358 5681
rect 16302 5607 16358 5616
rect 16316 4593 16344 5607
rect 16408 5030 16436 5714
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4865 16436 4966
rect 16394 4856 16450 4865
rect 16500 4826 16528 7142
rect 16684 5137 16712 8622
rect 16868 8265 16896 9862
rect 16854 8256 16910 8265
rect 16854 8191 16910 8200
rect 16960 8072 16988 10254
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17052 8974 17080 9454
rect 17144 9382 17172 9998
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8634 17080 8910
rect 17236 8906 17264 10066
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16868 8044 16988 8072
rect 16868 6225 16896 8044
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7546 16988 7890
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7698 17172 7822
rect 17144 7670 17264 7698
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17236 7206 17264 7670
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 16948 6248 17000 6254
rect 16854 6216 16910 6225
rect 16948 6190 17000 6196
rect 16854 6151 16910 6160
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16762 5400 16818 5409
rect 16762 5335 16818 5344
rect 16776 5166 16804 5335
rect 16868 5273 16896 6054
rect 16960 5778 16988 6190
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 16764 5160 16816 5166
rect 16670 5128 16726 5137
rect 16764 5102 16816 5108
rect 16670 5063 16726 5072
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16394 4791 16450 4800
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16302 4584 16358 4593
rect 16302 4519 16358 4528
rect 16408 4078 16436 4694
rect 16960 4321 16988 4966
rect 17144 4758 17172 6598
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16946 4312 17002 4321
rect 16946 4247 17002 4256
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16960 3670 16988 4082
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16408 2922 16436 3470
rect 16672 3392 16724 3398
rect 16500 3340 16672 3346
rect 16500 3334 16724 3340
rect 16500 3318 16712 3334
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16210 2544 16266 2553
rect 15934 2479 15936 2488
rect 15988 2479 15990 2488
rect 16120 2508 16172 2514
rect 15936 2450 15988 2456
rect 16210 2479 16266 2488
rect 16120 2450 16172 2456
rect 16500 2446 16528 3318
rect 16960 3194 16988 3606
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16764 3120 16816 3126
rect 16578 3088 16634 3097
rect 16578 3023 16634 3032
rect 16762 3088 16764 3097
rect 16816 3088 16818 3097
rect 16762 3023 16818 3032
rect 16396 2440 16448 2446
rect 16394 2408 16396 2417
rect 16488 2440 16540 2446
rect 16448 2408 16450 2417
rect 15384 2372 15436 2378
rect 16488 2382 16540 2388
rect 16394 2343 16450 2352
rect 15384 2314 15436 2320
rect 15934 1592 15990 1601
rect 15934 1527 15990 1536
rect 15948 480 15976 1527
rect 16592 480 16620 3023
rect 16960 2854 16988 3130
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16960 2650 16988 2790
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17144 610 17172 4422
rect 17236 3505 17264 7142
rect 17328 6848 17356 21286
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 17377 17448 17750
rect 17406 17368 17462 17377
rect 17406 17303 17408 17312
rect 17460 17303 17462 17312
rect 17408 17274 17460 17280
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17420 14958 17448 15506
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17420 14618 17448 14894
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17406 14240 17462 14249
rect 17406 14175 17462 14184
rect 17420 10198 17448 14175
rect 17604 13734 17632 25230
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24750 18184 25094
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17696 23322 17724 24074
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17788 23633 17816 24006
rect 17774 23624 17830 23633
rect 17774 23559 17830 23568
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 18064 22778 18092 24210
rect 18156 23322 18184 24550
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18340 23526 18368 24210
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18432 23594 18460 24142
rect 18510 23624 18566 23633
rect 18420 23588 18472 23594
rect 18510 23559 18566 23568
rect 18420 23530 18472 23536
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 18156 22574 18184 23258
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18156 21350 18184 21966
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 17682 21176 17738 21185
rect 17682 21111 17738 21120
rect 17696 19009 17724 21111
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17880 20602 17908 20878
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17880 20058 17908 20538
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17682 19000 17738 19009
rect 17682 18935 17738 18944
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17696 18426 17724 18770
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17788 16289 17816 19178
rect 17866 19000 17922 19009
rect 17866 18935 17922 18944
rect 17774 16280 17830 16289
rect 17774 16215 17830 16224
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17592 13728 17644 13734
rect 17788 13705 17816 13806
rect 17592 13670 17644 13676
rect 17774 13696 17830 13705
rect 17774 13631 17830 13640
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12646 17540 13330
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12986 17724 13262
rect 17684 12980 17736 12986
rect 17604 12940 17684 12968
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17498 12472 17554 12481
rect 17498 12407 17500 12416
rect 17552 12407 17554 12416
rect 17500 12378 17552 12384
rect 17604 11626 17632 12940
rect 17684 12922 17736 12928
rect 17880 12866 17908 18935
rect 17972 14521 18000 20742
rect 18064 20058 18092 21286
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18064 19310 18092 19994
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18050 17640 18106 17649
rect 18156 17626 18184 21286
rect 18340 19145 18368 23462
rect 18524 22642 18552 23559
rect 18708 23497 18736 27520
rect 18972 24948 19024 24954
rect 18972 24890 19024 24896
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18892 23730 18920 24006
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18694 23488 18750 23497
rect 18694 23423 18750 23432
rect 18892 23254 18920 23666
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18892 22778 18920 23190
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18524 22234 18552 22578
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21010 18644 21830
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18708 20330 18736 21898
rect 18892 21690 18920 22714
rect 18984 22234 19012 24890
rect 19352 23905 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20088 25498 20116 27520
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19444 24682 19472 25298
rect 20074 24848 20130 24857
rect 19524 24812 19576 24818
rect 20074 24783 20130 24792
rect 19524 24754 19576 24760
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19338 23896 19394 23905
rect 19338 23831 19394 23840
rect 19260 23594 19380 23610
rect 19248 23588 19380 23594
rect 19300 23582 19380 23588
rect 19248 23530 19300 23536
rect 19352 23322 19380 23582
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19536 23202 19564 24754
rect 20088 24614 20116 24783
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19352 23174 19564 23202
rect 19246 22672 19302 22681
rect 19246 22607 19302 22616
rect 19260 22409 19288 22607
rect 19246 22400 19302 22409
rect 19246 22335 19302 22344
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18892 20398 18920 21626
rect 19168 21457 19196 22170
rect 19260 22098 19288 22335
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19154 21448 19210 21457
rect 19154 21383 19210 21392
rect 19168 21078 19196 21383
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18616 19514 18644 19858
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18708 19417 18736 20266
rect 19260 20058 19288 20946
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 18694 19408 18750 19417
rect 18694 19343 18696 19352
rect 18748 19343 18750 19352
rect 18696 19314 18748 19320
rect 18696 19168 18748 19174
rect 18326 19136 18382 19145
rect 18696 19110 18748 19116
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 18326 19071 18382 19080
rect 18106 17598 18184 17626
rect 18050 17575 18106 17584
rect 18064 14618 18092 17575
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18340 16726 18368 17478
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18248 15609 18276 16390
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18234 15600 18290 15609
rect 18234 15535 18290 15544
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18248 14890 18276 15302
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17958 14512 18014 14521
rect 18064 14498 18092 14554
rect 18064 14470 18184 14498
rect 17958 14447 18014 14456
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18064 14074 18092 14350
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18156 13870 18184 14470
rect 18248 14278 18276 14826
rect 18616 14521 18644 15846
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13938 18276 14214
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18248 13530 18276 13874
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 17696 12838 17908 12866
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9110 17448 9998
rect 17696 9738 17724 12838
rect 18432 12646 18460 13262
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18064 12442 18092 12582
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18248 11082 18276 11562
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18432 10305 18460 12582
rect 18418 10296 18474 10305
rect 18418 10231 18474 10240
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17604 9710 17724 9738
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17408 6860 17460 6866
rect 17328 6820 17408 6848
rect 17328 5953 17356 6820
rect 17408 6802 17460 6808
rect 17314 5944 17370 5953
rect 17314 5879 17370 5888
rect 17408 5908 17460 5914
rect 17328 5574 17356 5879
rect 17408 5850 17460 5856
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 17328 3194 17356 4762
rect 17420 4622 17448 5850
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 4282 17448 4558
rect 17512 4457 17540 7482
rect 17604 6916 17632 9710
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 17696 8090 17724 9522
rect 17866 9480 17922 9489
rect 17866 9415 17868 9424
rect 17920 9415 17922 9424
rect 17868 9386 17920 9392
rect 18248 9178 18276 9522
rect 18340 9382 18368 9862
rect 18510 9616 18566 9625
rect 18510 9551 18566 9560
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18340 9058 18368 9318
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18248 9030 18368 9058
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17788 7818 17816 8910
rect 18156 8634 18184 8978
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 7886 17908 8434
rect 18156 8401 18184 8570
rect 17958 8392 18014 8401
rect 17958 8327 17960 8336
rect 18012 8327 18014 8336
rect 18142 8392 18198 8401
rect 18142 8327 18198 8336
rect 17960 8298 18012 8304
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 8129 18092 8230
rect 18050 8120 18106 8129
rect 18050 8055 18106 8064
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18156 7993 18184 8026
rect 18142 7984 18198 7993
rect 18142 7919 18198 7928
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7546 17816 7754
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 7002 18092 7142
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17684 6928 17736 6934
rect 17604 6888 17684 6916
rect 17684 6870 17736 6876
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17604 6322 17632 6734
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17604 5846 17632 6258
rect 17696 6118 17724 6870
rect 18144 6656 18196 6662
rect 18248 6644 18276 9030
rect 18524 8430 18552 9551
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18196 6616 18276 6644
rect 18144 6598 18196 6604
rect 18156 6118 18184 6598
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17604 4690 17632 5782
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17592 4480 17644 4486
rect 17498 4448 17554 4457
rect 17592 4422 17644 4428
rect 17498 4383 17554 4392
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17604 2922 17632 4422
rect 17696 4185 17724 6054
rect 17776 5024 17828 5030
rect 17774 4992 17776 5001
rect 17828 4992 17830 5001
rect 17774 4927 17830 4936
rect 17972 4842 18000 6054
rect 17880 4826 18000 4842
rect 18340 4826 18368 8366
rect 18708 8362 18736 19110
rect 19168 18970 19196 19110
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19260 18834 19288 19790
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19246 18184 19302 18193
rect 19064 18148 19116 18154
rect 19246 18119 19302 18128
rect 19064 18090 19116 18096
rect 19076 17542 19104 18090
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18880 17060 18932 17066
rect 18880 17002 18932 17008
rect 18892 16794 18920 17002
rect 19076 16998 19104 17478
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 19076 16114 19104 16934
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19062 16008 19118 16017
rect 19062 15943 19118 15952
rect 19156 15972 19208 15978
rect 19076 15910 19104 15943
rect 19156 15914 19208 15920
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19168 15706 19196 15914
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 18972 14272 19024 14278
rect 19260 14249 19288 18119
rect 19352 17105 19380 23174
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 21486 19656 21830
rect 19616 21480 19668 21486
rect 19536 21440 19616 21468
rect 19536 20602 19564 21440
rect 19616 21422 19668 21428
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 20596 19576 20602
rect 19444 20556 19524 20584
rect 19444 19854 19472 20556
rect 19524 20538 19576 20544
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19444 19009 19472 19110
rect 19430 19000 19486 19009
rect 19536 18970 19564 19926
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20088 19310 20116 19858
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19996 18970 20024 19110
rect 19430 18935 19486 18944
rect 19524 18964 19576 18970
rect 19444 18902 19472 18935
rect 19524 18906 19576 18912
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 20088 18902 20116 19110
rect 19432 18896 19484 18902
rect 20076 18896 20128 18902
rect 19432 18838 19484 18844
rect 19798 18864 19854 18873
rect 20076 18838 20128 18844
rect 19798 18799 19800 18808
rect 19852 18799 19854 18808
rect 19800 18770 19852 18776
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18329 20024 18566
rect 19982 18320 20038 18329
rect 19982 18255 20038 18264
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20074 17912 20130 17921
rect 20074 17847 20076 17856
rect 20128 17847 20130 17856
rect 20076 17818 20128 17824
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19812 17649 19840 17682
rect 19798 17640 19854 17649
rect 19798 17575 19854 17584
rect 19338 17096 19394 17105
rect 19338 17031 19394 17040
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 14618 19472 15438
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 18972 14214 19024 14220
rect 19246 14240 19302 14249
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18800 12782 18828 13330
rect 18788 12776 18840 12782
rect 18786 12744 18788 12753
rect 18840 12744 18842 12753
rect 18786 12679 18842 12688
rect 18984 11937 19012 14214
rect 19246 14175 19302 14184
rect 19352 13938 19380 14282
rect 19444 14074 19472 14554
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19352 13530 19380 13874
rect 19430 13560 19486 13569
rect 19340 13524 19392 13530
rect 19430 13495 19486 13504
rect 19340 13466 19392 13472
rect 19444 13462 19472 13495
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19536 13394 19564 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20088 15706 20116 15982
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14346 20024 14758
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19628 13870 19656 14010
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19062 12744 19118 12753
rect 19260 12714 19288 13194
rect 19352 12782 19380 13194
rect 19628 12918 19656 13398
rect 20180 13025 20208 24618
rect 20732 24426 20760 27520
rect 21376 24857 21404 27520
rect 21914 27160 21970 27169
rect 21914 27095 21970 27104
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21362 24848 21418 24857
rect 21362 24783 21418 24792
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 20640 24410 20760 24426
rect 20628 24404 20760 24410
rect 20680 24398 20760 24404
rect 21454 24440 21510 24449
rect 21454 24375 21456 24384
rect 20628 24346 20680 24352
rect 21508 24375 21510 24384
rect 21456 24346 21508 24352
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20626 23760 20682 23769
rect 20626 23695 20682 23704
rect 20640 23526 20668 23695
rect 21100 23526 21128 24210
rect 21362 23624 21418 23633
rect 21362 23559 21418 23568
rect 21376 23526 21404 23559
rect 20628 23520 20680 23526
rect 20812 23520 20864 23526
rect 20680 23480 20760 23508
rect 20628 23462 20680 23468
rect 20732 23118 20760 23480
rect 20812 23462 20864 23468
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 21364 23520 21416 23526
rect 21560 23474 21588 24686
rect 21652 23662 21680 25094
rect 21732 24880 21784 24886
rect 21732 24822 21784 24828
rect 21744 23730 21772 24822
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21364 23462 21416 23468
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20272 22234 20300 22442
rect 20350 22400 20406 22409
rect 20350 22335 20406 22344
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20272 21690 20300 22170
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20272 20942 20300 21626
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20272 20602 20300 20878
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20364 19825 20392 22335
rect 20732 22234 20760 23054
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20456 20482 20484 20742
rect 20456 20466 20760 20482
rect 20456 20460 20772 20466
rect 20456 20454 20720 20460
rect 20350 19816 20406 19825
rect 20350 19751 20406 19760
rect 20456 19417 20484 20454
rect 20720 20402 20772 20408
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19990 20576 20198
rect 20536 19984 20588 19990
rect 20824 19938 20852 23462
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20902 23080 20958 23089
rect 20902 23015 20904 23024
rect 20956 23015 20958 23024
rect 20904 22986 20956 22992
rect 21008 22930 21036 23122
rect 20916 22902 21036 22930
rect 20916 22574 20944 22902
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20916 20262 20944 22510
rect 21100 20641 21128 23462
rect 21468 23446 21588 23474
rect 21362 22536 21418 22545
rect 21362 22471 21418 22480
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21086 20632 21142 20641
rect 21086 20567 21142 20576
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 20058 20944 20198
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20916 19961 20944 19994
rect 20536 19926 20588 19932
rect 20640 19922 20852 19938
rect 20628 19916 20852 19922
rect 20680 19910 20852 19916
rect 20628 19858 20680 19864
rect 20442 19408 20498 19417
rect 20442 19343 20498 19352
rect 20350 18864 20406 18873
rect 20350 18799 20406 18808
rect 20364 17882 20392 18799
rect 20456 18426 20484 19343
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20720 18148 20772 18154
rect 20548 18108 20720 18136
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20258 17776 20314 17785
rect 20258 17711 20314 17720
rect 20272 16674 20300 17711
rect 20350 17640 20406 17649
rect 20350 17575 20406 17584
rect 20364 16794 20392 17575
rect 20442 17504 20498 17513
rect 20442 17439 20498 17448
rect 20456 17338 20484 17439
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20272 16646 20392 16674
rect 20166 13016 20222 13025
rect 20166 12951 20222 12960
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19340 12776 19392 12782
rect 19392 12736 19472 12764
rect 19340 12718 19392 12724
rect 19062 12679 19118 12688
rect 19248 12708 19300 12714
rect 19076 12442 19104 12679
rect 19248 12650 19300 12656
rect 19156 12640 19208 12646
rect 19444 12594 19472 12736
rect 19156 12582 19208 12588
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18970 11928 19026 11937
rect 18970 11863 19026 11872
rect 19168 11506 19196 12582
rect 19260 12566 19472 12594
rect 19260 12306 19288 12566
rect 19536 12458 19564 12786
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19444 12430 19564 12458
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19444 12102 19472 12430
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19076 11478 19196 11506
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18800 9489 18828 10066
rect 18892 10044 18920 10746
rect 18972 10056 19024 10062
rect 18892 10016 18972 10044
rect 18892 9586 18920 10016
rect 18972 9998 19024 10004
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18786 9480 18842 9489
rect 18842 9438 18920 9466
rect 18786 9415 18842 9424
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8498 18828 8774
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18524 7857 18552 7890
rect 18604 7880 18656 7886
rect 18510 7848 18566 7857
rect 18604 7822 18656 7828
rect 18510 7783 18566 7792
rect 18524 7546 18552 7783
rect 18616 7546 18644 7822
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18510 6896 18566 6905
rect 18510 6831 18566 6840
rect 18418 6760 18474 6769
rect 18524 6730 18552 6831
rect 18418 6695 18474 6704
rect 18512 6724 18564 6730
rect 18432 6254 18460 6695
rect 18512 6666 18564 6672
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 17868 4820 18000 4826
rect 17920 4814 18000 4820
rect 18328 4820 18380 4826
rect 17868 4762 17920 4768
rect 18328 4762 18380 4768
rect 17682 4176 17738 4185
rect 18340 4146 18368 4762
rect 18432 4185 18460 4966
rect 18418 4176 18474 4185
rect 17682 4111 17738 4120
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 18328 4140 18380 4146
rect 18418 4111 18474 4120
rect 18328 4082 18380 4088
rect 17788 3942 17816 4082
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 17788 3641 17816 3878
rect 18142 3768 18198 3777
rect 18142 3703 18198 3712
rect 17774 3632 17830 3641
rect 17774 3567 17830 3576
rect 18156 3466 18184 3703
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 17958 2952 18014 2961
rect 17592 2916 17644 2922
rect 17958 2887 18014 2896
rect 17592 2858 17644 2864
rect 17224 2304 17276 2310
rect 17222 2272 17224 2281
rect 17276 2272 17278 2281
rect 17222 2207 17278 2216
rect 17132 604 17184 610
rect 17132 546 17184 552
rect 17316 604 17368 610
rect 17316 546 17368 552
rect 17328 480 17356 546
rect 17972 480 18000 2887
rect 18156 2650 18184 3402
rect 18340 2990 18368 3878
rect 18420 3392 18472 3398
rect 18524 3369 18552 6054
rect 18616 5914 18644 6666
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18800 4729 18828 7482
rect 18892 6866 18920 9438
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18892 6458 18920 6802
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18984 5914 19012 6938
rect 19076 6497 19104 11478
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19168 10606 19196 11290
rect 19260 11257 19288 12038
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11354 19472 11494
rect 19536 11354 19564 12310
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19246 11248 19302 11257
rect 19246 11183 19302 11192
rect 19522 11112 19578 11121
rect 19996 11082 20024 12242
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 12073 20116 12174
rect 20074 12064 20130 12073
rect 20074 11999 20130 12008
rect 20088 11898 20116 11999
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 19522 11047 19578 11056
rect 19984 11076 20036 11082
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19430 10296 19486 10305
rect 19430 10231 19486 10240
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19168 9382 19196 10066
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19168 6769 19196 9318
rect 19444 9178 19472 10231
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8362 19380 8978
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 8242 19380 8298
rect 19260 8214 19380 8242
rect 19154 6760 19210 6769
rect 19154 6695 19210 6704
rect 19062 6488 19118 6497
rect 19062 6423 19118 6432
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19076 5914 19104 6258
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18984 4826 19012 5170
rect 19260 4826 19288 8214
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7274 19380 7686
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 7177 19380 7210
rect 19338 7168 19394 7177
rect 19338 7103 19394 7112
rect 19444 6458 19472 7346
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19536 5930 19564 11047
rect 19984 11018 20036 11024
rect 20272 11014 20300 11562
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20272 10470 20300 10950
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 20272 9602 20300 10406
rect 20180 9574 20300 9602
rect 20180 9518 20208 9574
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19982 7848 20038 7857
rect 19720 7313 19748 7822
rect 19982 7783 20038 7792
rect 19706 7304 19762 7313
rect 19706 7239 19762 7248
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19720 6254 19748 6598
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19352 5902 19564 5930
rect 19352 5273 19380 5902
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19536 5370 19564 5714
rect 19996 5370 20024 7783
rect 20088 7546 20116 8298
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19338 5264 19394 5273
rect 19338 5199 19394 5208
rect 19352 5166 19380 5199
rect 19996 5166 20024 5306
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19524 5092 19576 5098
rect 19524 5034 19576 5040
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 18786 4720 18842 4729
rect 18786 4655 18842 4664
rect 18694 4312 18750 4321
rect 18694 4247 18750 4256
rect 18420 3334 18472 3340
rect 18510 3360 18566 3369
rect 18432 2990 18460 3334
rect 18510 3295 18566 3304
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18326 2408 18382 2417
rect 18326 2343 18328 2352
rect 18380 2343 18382 2352
rect 18328 2314 18380 2320
rect 18708 480 18736 4247
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18892 3466 18920 4082
rect 18984 4010 19012 4762
rect 19536 4457 19564 5034
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4690 20024 4966
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19892 4616 19944 4622
rect 19892 4558 19944 4564
rect 19904 4457 19932 4558
rect 19522 4448 19578 4457
rect 19444 4406 19522 4434
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 19444 3738 19472 4406
rect 19522 4383 19578 4392
rect 19890 4448 19946 4457
rect 19890 4383 19946 4392
rect 19904 4282 19932 4383
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3738 20024 4626
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 20088 3670 20116 3946
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19432 3528 19484 3534
rect 19338 3496 19394 3505
rect 18880 3460 18932 3466
rect 19394 3476 19432 3482
rect 19394 3470 19484 3476
rect 19394 3454 19472 3470
rect 19338 3431 19394 3440
rect 18880 3402 18932 3408
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18800 2310 18828 2382
rect 18984 2378 19012 3334
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 19352 2310 19380 3431
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2650 20024 3538
rect 20088 3194 20116 3606
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20180 2514 20208 8842
rect 20272 8430 20300 9114
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20364 6934 20392 16646
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 16114 20484 16390
rect 20548 16250 20576 18108
rect 20720 18090 20772 18096
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20732 17241 20760 17682
rect 20718 17232 20774 17241
rect 20718 17167 20720 17176
rect 20772 17167 20774 17176
rect 20720 17138 20772 17144
rect 20824 17134 20852 19910
rect 20902 19952 20958 19961
rect 20902 19887 20958 19896
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20916 19446 20944 19790
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20916 17270 20944 19382
rect 21008 19378 21036 19858
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21008 18698 21036 19314
rect 21192 18850 21220 21966
rect 21284 21350 21312 22034
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21284 19514 21312 21286
rect 21376 20913 21404 22471
rect 21362 20904 21418 20913
rect 21362 20839 21418 20848
rect 21362 19816 21418 19825
rect 21362 19751 21418 19760
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21192 18822 21312 18850
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 21192 18222 21220 18702
rect 21180 18216 21232 18222
rect 21178 18184 21180 18193
rect 21232 18184 21234 18193
rect 21178 18119 21234 18128
rect 20994 17776 21050 17785
rect 20994 17711 21050 17720
rect 21008 17338 21036 17711
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20640 16266 20668 16594
rect 20916 16590 20944 17206
rect 21008 16998 21036 17274
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20640 16250 20760 16266
rect 20536 16244 20588 16250
rect 20640 16244 20772 16250
rect 20640 16238 20720 16244
rect 20536 16186 20588 16192
rect 20720 16186 20772 16192
rect 20916 16182 20944 16526
rect 21284 16425 21312 18822
rect 21270 16416 21326 16425
rect 21270 16351 21326 16360
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 15706 20484 16050
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20916 15502 20944 16118
rect 21376 15722 21404 19751
rect 21468 18766 21496 23446
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21652 22234 21680 23258
rect 21744 22982 21772 23666
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21836 22658 21864 24550
rect 21928 24410 21956 27095
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22020 24886 22048 25298
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 21928 23594 21956 24346
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22778 21956 22918
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 21836 22630 21956 22658
rect 21732 22500 21784 22506
rect 21732 22442 21784 22448
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21652 20398 21680 22170
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21546 19272 21602 19281
rect 21546 19207 21602 19216
rect 21560 18902 21588 19207
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18970 21680 19110
rect 21640 18964 21692 18970
rect 21640 18906 21692 18912
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 16017 21496 18022
rect 21560 17882 21588 18838
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21652 17202 21680 17614
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21652 16658 21680 17138
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21454 16008 21510 16017
rect 21454 15943 21510 15952
rect 21376 15694 21588 15722
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 15094 20944 15438
rect 20904 15088 20956 15094
rect 20824 15048 20904 15076
rect 20824 14074 20852 15048
rect 20904 15030 20956 15036
rect 21376 14822 21404 15574
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20824 13138 20852 14010
rect 20916 14006 20944 14418
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20904 14000 20956 14006
rect 20902 13968 20904 13977
rect 20956 13968 20958 13977
rect 20902 13903 20958 13912
rect 20916 13877 20944 13903
rect 21100 13841 21128 14214
rect 21376 14074 21404 14758
rect 21468 14618 21496 14894
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13326 21036 13670
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20640 12782 20668 13126
rect 20824 13110 20944 13138
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20456 12102 20484 12650
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 12442 20576 12582
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11665 20484 12038
rect 20536 11688 20588 11694
rect 20442 11656 20498 11665
rect 20536 11630 20588 11636
rect 20442 11591 20498 11600
rect 20548 8362 20576 11630
rect 20640 11354 20668 12718
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20626 11248 20682 11257
rect 20626 11183 20682 11192
rect 20640 8616 20668 11183
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10810 20760 10950
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20732 9722 20760 10474
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20824 9450 20852 12922
rect 20916 12306 20944 13110
rect 21100 12646 21128 13330
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12986 21404 13262
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21560 12866 21588 15694
rect 21744 15162 21772 22442
rect 21928 22030 21956 22630
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21836 20942 21864 21286
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 20262 21864 20878
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21836 19446 21864 20198
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21928 18193 21956 21830
rect 21914 18184 21970 18193
rect 21914 18119 21970 18128
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17338 21864 18022
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21914 14512 21970 14521
rect 21914 14447 21916 14456
rect 21968 14447 21970 14456
rect 21916 14418 21968 14424
rect 21928 14006 21956 14418
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21652 13326 21680 13670
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 12986 21680 13262
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21364 12844 21416 12850
rect 21560 12838 21680 12866
rect 21928 12850 21956 13126
rect 21364 12786 21416 12792
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20916 11898 20944 12242
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20916 11354 20944 11834
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 21100 9518 21128 12582
rect 21376 12374 21404 12786
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21546 11112 21602 11121
rect 21546 11047 21602 11056
rect 21270 10568 21326 10577
rect 21270 10503 21326 10512
rect 21284 10266 21312 10503
rect 21362 10296 21418 10305
rect 21272 10260 21324 10266
rect 21362 10231 21418 10240
rect 21272 10202 21324 10208
rect 21376 10062 21404 10231
rect 21364 10056 21416 10062
rect 21362 10024 21364 10033
rect 21456 10056 21508 10062
rect 21416 10024 21418 10033
rect 21456 9998 21508 10004
rect 21362 9959 21418 9968
rect 21376 9722 21404 9959
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21468 9654 21496 9998
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20824 9353 20852 9386
rect 20810 9344 20866 9353
rect 20810 9279 20866 9288
rect 21100 9217 21128 9454
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21086 9208 21142 9217
rect 21086 9143 21142 9152
rect 21086 8936 21142 8945
rect 21086 8871 21142 8880
rect 20720 8628 20772 8634
rect 20640 8588 20720 8616
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20640 7750 20668 8588
rect 20720 8570 20772 8576
rect 20994 8392 21050 8401
rect 20994 8327 21050 8336
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20352 6928 20404 6934
rect 20272 6888 20352 6916
rect 20272 5778 20300 6888
rect 20352 6870 20404 6876
rect 20824 6730 20852 7142
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20718 5672 20774 5681
rect 20824 5642 20852 6666
rect 20916 6662 20944 7890
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20718 5607 20774 5616
rect 20812 5636 20864 5642
rect 20732 5574 20760 5607
rect 20812 5578 20864 5584
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20364 5234 20392 5510
rect 20824 5370 20852 5578
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4758 20392 4966
rect 20548 4758 20576 5170
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20456 3738 20484 4490
rect 20824 4078 20852 4558
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20916 3777 20944 6598
rect 21008 6202 21036 8327
rect 21100 8090 21128 8871
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21468 7546 21496 9318
rect 21560 9178 21588 11047
rect 21652 9654 21680 12838
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21928 11898 21956 12786
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21928 11150 21956 11834
rect 22020 11354 22048 24822
rect 22112 24682 22140 27520
rect 22756 25498 22784 27520
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22558 24848 22614 24857
rect 22558 24783 22614 24792
rect 22374 24712 22430 24721
rect 22100 24676 22152 24682
rect 22374 24647 22430 24656
rect 22100 24618 22152 24624
rect 22388 24614 22416 24647
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22572 24410 22600 24783
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 22388 23526 22416 24210
rect 22928 23588 22980 23594
rect 22928 23530 22980 23536
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22388 22409 22416 23462
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22374 22400 22430 22409
rect 22374 22335 22430 22344
rect 22100 22092 22152 22098
rect 22100 22034 22152 22040
rect 22112 21690 22140 22034
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22112 21146 22140 21626
rect 22388 21486 22416 21966
rect 22480 21554 22508 22918
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22940 21078 22968 23530
rect 23124 23526 23152 24210
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23018 23216 23074 23225
rect 23018 23151 23074 23160
rect 23032 23118 23060 23151
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 23032 22778 23060 23054
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23124 22506 23152 23462
rect 23308 22642 23336 27639
rect 23478 27520 23534 28000
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25502 27520 25558 28000
rect 26146 27520 26202 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 23386 26616 23442 26625
rect 23386 26551 23442 26560
rect 23400 23322 23428 26551
rect 23492 24449 23520 27520
rect 23570 25392 23626 25401
rect 23570 25327 23626 25336
rect 23584 24954 23612 25327
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 24136 24721 24164 27520
rect 24674 25936 24730 25945
rect 24674 25871 24730 25880
rect 24688 25158 24716 25871
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24857 24808 27520
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 25318 24848 25374 24857
rect 25318 24783 25374 24792
rect 24122 24712 24178 24721
rect 24122 24647 24178 24656
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23754 24576 23810 24585
rect 23478 24440 23534 24449
rect 23478 24375 23534 24384
rect 23570 24168 23626 24177
rect 23570 24103 23626 24112
rect 23478 23624 23534 23633
rect 23478 23559 23534 23568
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23400 22778 23428 23258
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 23296 22432 23348 22438
rect 23294 22400 23296 22409
rect 23348 22400 23350 22409
rect 23294 22335 23350 22344
rect 23400 22234 23428 22578
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23400 22098 23428 22170
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21350 23152 21966
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 22928 21072 22980 21078
rect 22928 21014 22980 21020
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22112 20602 22140 20946
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22112 20058 22140 20538
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22112 19514 22140 19994
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22928 19440 22980 19446
rect 22650 19408 22706 19417
rect 22928 19382 22980 19388
rect 22650 19343 22706 19352
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22112 17134 22140 18226
rect 22204 18154 22232 18566
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22112 16794 22140 17070
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22204 16114 22232 17546
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 17338 22324 17478
rect 22480 17338 22508 17750
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22388 16114 22416 16730
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22204 15162 22232 16050
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 12782 22140 13126
rect 22100 12776 22152 12782
rect 22098 12744 22100 12753
rect 22152 12744 22154 12753
rect 22098 12679 22154 12688
rect 22204 12345 22232 14214
rect 22572 13161 22600 18770
rect 22664 15162 22692 19343
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22756 18766 22784 19110
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22756 18426 22784 18702
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22756 13258 22784 14214
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22558 13152 22614 13161
rect 22558 13087 22614 13096
rect 22282 13016 22338 13025
rect 22282 12951 22284 12960
rect 22336 12951 22338 12960
rect 22284 12922 22336 12928
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22190 12336 22246 12345
rect 22190 12271 22246 12280
rect 22468 12096 22520 12102
rect 22466 12064 22468 12073
rect 22520 12064 22522 12073
rect 22466 11999 22522 12008
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22480 11286 22508 11999
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21928 10674 21956 11086
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21744 9994 21772 10406
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21836 9722 21864 10202
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 22112 9178 22140 10950
rect 22388 10810 22416 11154
rect 22480 10810 22508 11222
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22296 9058 22324 9318
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 22204 9030 22324 9058
rect 21928 8566 21956 8978
rect 22204 8974 22232 9030
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22204 8634 22232 8910
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 21916 8560 21968 8566
rect 21914 8528 21916 8537
rect 22284 8560 22336 8566
rect 21968 8528 21970 8537
rect 22284 8502 22336 8508
rect 21914 8463 21970 8472
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21744 7886 21772 8298
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21270 7440 21326 7449
rect 21270 7375 21326 7384
rect 21008 6174 21128 6202
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 21008 5914 21036 6054
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 21008 4282 21036 4694
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20994 4040 21050 4049
rect 20994 3975 21050 3984
rect 20902 3768 20958 3777
rect 20444 3732 20496 3738
rect 20902 3703 20958 3712
rect 20444 3674 20496 3680
rect 21008 3641 21036 3975
rect 20994 3632 21050 3641
rect 20994 3567 21050 3576
rect 20718 3224 20774 3233
rect 20718 3159 20774 3168
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 19352 1601 19380 2246
rect 19430 1728 19486 1737
rect 19430 1663 19486 1672
rect 19338 1592 19394 1601
rect 19338 1527 19394 1536
rect 19444 1170 19472 1663
rect 19352 1142 19472 1170
rect 19352 480 19380 1142
rect 20088 480 20116 2246
rect 20732 480 20760 3159
rect 21100 3126 21128 6174
rect 21284 5846 21312 7375
rect 21560 7206 21588 7822
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22112 7698 22140 7754
rect 21836 7670 22140 7698
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21362 6488 21418 6497
rect 21362 6423 21418 6432
rect 21376 5914 21404 6423
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21178 4992 21234 5001
rect 21178 4927 21234 4936
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 21100 2922 21128 3062
rect 21192 2990 21220 4927
rect 21284 4826 21312 5782
rect 21376 5370 21404 5850
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21362 4176 21418 4185
rect 21362 4111 21418 4120
rect 21376 3738 21404 4111
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21284 3194 21312 3538
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 21192 2650 21220 2926
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21284 921 21312 2858
rect 21376 2650 21404 3674
rect 21468 3534 21496 4218
rect 21560 4185 21588 7142
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21652 6390 21680 6870
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21744 6458 21772 6734
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21640 6384 21692 6390
rect 21638 6352 21640 6361
rect 21692 6352 21694 6361
rect 21638 6287 21694 6296
rect 21836 5370 21864 7670
rect 22204 7410 22232 7686
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22204 7290 22232 7346
rect 21928 7262 22232 7290
rect 21928 6730 21956 7262
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22020 6934 22048 7142
rect 22008 6928 22060 6934
rect 22100 6928 22152 6934
rect 22008 6870 22060 6876
rect 22098 6896 22100 6905
rect 22152 6896 22154 6905
rect 22296 6866 22324 8502
rect 22388 7478 22416 8774
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22480 7818 22508 8366
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22388 7342 22416 7414
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22098 6831 22154 6840
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 22112 5914 22140 6734
rect 22296 6254 22324 6802
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22572 5778 22600 12854
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22756 11937 22784 12242
rect 22742 11928 22798 11937
rect 22742 11863 22744 11872
rect 22796 11863 22798 11872
rect 22744 11834 22796 11840
rect 22756 11803 22784 11834
rect 22940 9704 22968 19382
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 15910 23060 18770
rect 23202 18728 23258 18737
rect 23202 18663 23258 18672
rect 23216 18426 23244 18663
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23204 18148 23256 18154
rect 23204 18090 23256 18096
rect 23216 17814 23244 18090
rect 23308 17814 23336 21830
rect 23400 21146 23428 22034
rect 23492 21865 23520 23559
rect 23584 22681 23612 24103
rect 23676 23322 23704 24550
rect 23754 24511 23810 24520
rect 23768 24410 23796 24511
rect 24766 24440 24822 24449
rect 23756 24404 23808 24410
rect 24766 24375 24768 24384
rect 23756 24346 23808 24352
rect 24820 24375 24822 24384
rect 24768 24346 24820 24352
rect 24216 24268 24268 24274
rect 24216 24210 24268 24216
rect 24228 23730 24256 24210
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24766 23896 24822 23905
rect 24766 23831 24768 23840
rect 24820 23831 24822 23840
rect 24768 23802 24820 23808
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 23570 22672 23626 22681
rect 23952 22642 23980 23054
rect 23570 22607 23626 22616
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 24044 22574 24072 23258
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 23676 22166 23704 22374
rect 23664 22160 23716 22166
rect 23664 22102 23716 22108
rect 23478 21856 23534 21865
rect 23478 21791 23534 21800
rect 23768 21706 23796 22374
rect 24136 22098 24164 23462
rect 24228 22438 24256 23666
rect 24766 23488 24822 23497
rect 24766 23423 24822 23432
rect 24780 23322 24808 23423
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22438 24716 23122
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 24216 21888 24268 21894
rect 24596 21876 24624 22034
rect 24688 22012 24716 22374
rect 24688 21984 24900 22012
rect 24596 21848 24716 21876
rect 24216 21830 24268 21836
rect 23492 21678 23796 21706
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23492 18834 23520 21678
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23662 21312 23718 21321
rect 23662 21247 23718 21256
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23584 20602 23612 21014
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23400 17762 23428 18702
rect 23584 18154 23612 20538
rect 23676 20074 23704 21247
rect 23768 21146 23796 21490
rect 24228 21486 24256 21830
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23754 21040 23810 21049
rect 23754 20975 23810 20984
rect 23768 20942 23796 20975
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23676 20046 23796 20074
rect 23662 19952 23718 19961
rect 23662 19887 23718 19896
rect 23676 18970 23704 19887
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23676 18222 23704 18906
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23572 18148 23624 18154
rect 23572 18090 23624 18096
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23676 17882 23704 18022
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23400 17734 23520 17762
rect 23296 17672 23348 17678
rect 23202 17640 23258 17649
rect 23296 17614 23348 17620
rect 23202 17575 23204 17584
rect 23256 17575 23258 17584
rect 23204 17546 23256 17552
rect 23202 17368 23258 17377
rect 23308 17354 23336 17614
rect 23258 17338 23336 17354
rect 23258 17332 23348 17338
rect 23258 17326 23296 17332
rect 23202 17303 23258 17312
rect 23216 16726 23244 17303
rect 23296 17274 23348 17280
rect 23308 17243 23336 17274
rect 23492 16726 23520 17734
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23584 16794 23612 17682
rect 23768 16946 23796 20046
rect 23860 19922 23888 21286
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23860 19242 23888 19858
rect 23952 19446 23980 20198
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23860 18766 23888 19178
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18873 23980 19110
rect 23938 18864 23994 18873
rect 23938 18799 23994 18808
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 18426 23888 18702
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 24044 17785 24072 20538
rect 24136 20398 24164 20742
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 20058 24164 20198
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24136 19310 24164 19994
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24228 19242 24256 20742
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24308 19440 24360 19446
rect 24308 19382 24360 19388
rect 24216 19236 24268 19242
rect 24216 19178 24268 19184
rect 24320 18970 24348 19382
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24596 18902 24624 19314
rect 24216 18896 24268 18902
rect 24216 18838 24268 18844
rect 24584 18896 24636 18902
rect 24584 18838 24636 18844
rect 24228 17882 24256 18838
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18408 24716 21848
rect 24766 21856 24822 21865
rect 24766 21791 24822 21800
rect 24780 20369 24808 21791
rect 24766 20360 24822 20369
rect 24872 20330 24900 21984
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 24950 20768 25006 20777
rect 24950 20703 25006 20712
rect 24766 20295 24822 20304
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24964 19530 24992 20703
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 25056 19990 25084 20402
rect 25148 20262 25176 20810
rect 25332 20602 25360 24783
rect 25516 24585 25544 27520
rect 25502 24576 25558 24585
rect 25502 24511 25558 24520
rect 26160 23497 26188 27520
rect 26896 24449 26924 27520
rect 26882 24440 26938 24449
rect 26882 24375 26938 24384
rect 27540 23905 27568 27520
rect 27526 23896 27582 23905
rect 27526 23831 27582 23840
rect 26146 23488 26202 23497
rect 26146 23423 26202 23432
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25424 22778 25452 23015
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25516 20942 25544 21286
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25516 20602 25544 20878
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25044 19984 25096 19990
rect 25044 19926 25096 19932
rect 24872 19514 24992 19530
rect 25056 19514 25084 19926
rect 24860 19508 24992 19514
rect 24912 19502 24992 19508
rect 25044 19508 25096 19514
rect 24860 19450 24912 19456
rect 25044 19450 25096 19456
rect 25148 19394 25176 20198
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25056 19366 25176 19394
rect 25332 19378 25360 19654
rect 25320 19372 25372 19378
rect 24766 19000 24822 19009
rect 24766 18935 24822 18944
rect 24596 18380 24716 18408
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24030 17776 24086 17785
rect 24030 17711 24086 17720
rect 24596 17610 24624 18380
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 23940 17604 23992 17610
rect 23940 17546 23992 17552
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 23676 16918 23796 16946
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23480 16720 23532 16726
rect 23480 16662 23532 16668
rect 23202 16416 23258 16425
rect 23202 16351 23258 16360
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 23032 12714 23060 15846
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 23124 13462 23152 13670
rect 23216 13530 23244 16351
rect 23492 16250 23520 16662
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23400 14006 23428 15030
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23572 13796 23624 13802
rect 23572 13738 23624 13744
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23112 13456 23164 13462
rect 23112 13398 23164 13404
rect 23124 12986 23152 13398
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23216 12918 23244 13466
rect 23584 13190 23612 13738
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 23020 12708 23072 12714
rect 23020 12650 23072 12656
rect 23584 12170 23612 13126
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 10266 23060 11494
rect 23388 10736 23440 10742
rect 23202 10704 23258 10713
rect 23388 10678 23440 10684
rect 23202 10639 23258 10648
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22848 9676 22968 9704
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7546 22692 7686
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22664 7410 22692 7482
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22756 6866 22784 7482
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22756 6458 22784 6802
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21730 5264 21786 5273
rect 21730 5199 21786 5208
rect 21546 4176 21602 4185
rect 21546 4111 21602 4120
rect 21546 4040 21602 4049
rect 21546 3975 21602 3984
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21468 3126 21496 3470
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21560 2961 21588 3975
rect 21546 2952 21602 2961
rect 21546 2887 21602 2896
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21744 2514 21772 5199
rect 22020 2666 22048 5714
rect 22558 5672 22614 5681
rect 22468 5636 22520 5642
rect 22558 5607 22614 5616
rect 22468 5578 22520 5584
rect 22480 5234 22508 5578
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22284 4480 22336 4486
rect 22282 4448 22284 4457
rect 22336 4448 22338 4457
rect 22282 4383 22338 4392
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22112 3641 22140 4014
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22098 3632 22154 3641
rect 22098 3567 22154 3576
rect 22296 3505 22324 3878
rect 22388 3738 22416 5102
rect 22572 3738 22600 5607
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22282 3496 22338 3505
rect 22282 3431 22338 3440
rect 22572 2990 22600 3674
rect 22664 3074 22692 6054
rect 22756 5302 22784 6394
rect 22848 5545 22876 9676
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 22940 7002 22968 7890
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 22928 5568 22980 5574
rect 22834 5536 22890 5545
rect 22928 5510 22980 5516
rect 22834 5471 22890 5480
rect 22744 5296 22796 5302
rect 22744 5238 22796 5244
rect 22756 4486 22784 5238
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22756 4282 22784 4422
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22756 4010 22784 4218
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 22664 3046 22876 3074
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22848 2666 22876 3046
rect 22020 2638 22140 2666
rect 21732 2508 21784 2514
rect 21732 2450 21784 2456
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 21362 1864 21418 1873
rect 21362 1799 21418 1808
rect 21270 912 21326 921
rect 21270 847 21326 856
rect 21376 480 21404 1799
rect 21928 1465 21956 2246
rect 21914 1456 21970 1465
rect 21914 1391 21970 1400
rect 22112 480 22140 2638
rect 22756 2638 22876 2666
rect 22756 480 22784 2638
rect 22834 2544 22890 2553
rect 22834 2479 22836 2488
rect 22888 2479 22890 2488
rect 22836 2450 22888 2456
rect 22940 610 22968 5510
rect 23032 5370 23060 5714
rect 23124 5574 23152 6870
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23124 5370 23152 5510
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23124 5234 23152 5306
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 23216 3670 23244 10639
rect 23400 10062 23428 10678
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23492 10198 23520 10406
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23400 9722 23428 9998
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23308 8634 23336 8910
rect 23400 8650 23428 9658
rect 23492 9450 23520 10134
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 23584 8838 23612 12106
rect 23676 11801 23704 16918
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23860 15910 23888 16526
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23952 15201 23980 17546
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17134 24716 18226
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24688 16794 24716 17070
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24030 16688 24086 16697
rect 24030 16623 24086 16632
rect 24044 15570 24072 16623
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24122 16280 24178 16289
rect 24228 16250 24256 16526
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24122 16215 24178 16224
rect 24216 16244 24268 16250
rect 24136 16046 24164 16215
rect 24216 16186 24268 16192
rect 24780 16130 24808 18935
rect 24858 18184 24914 18193
rect 24858 18119 24914 18128
rect 24872 16658 24900 18119
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 17241 24992 17478
rect 24950 17232 25006 17241
rect 24950 17167 25006 17176
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24872 16250 24900 16594
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24688 16102 24808 16130
rect 25056 16114 25084 19366
rect 25320 19314 25372 19320
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18426 25268 18566
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25226 18320 25282 18329
rect 25226 18255 25282 18264
rect 25240 18222 25268 18255
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25424 17785 25452 18022
rect 25516 17921 25544 19246
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18465 25728 19110
rect 25686 18456 25742 18465
rect 25686 18391 25742 18400
rect 25502 17912 25558 17921
rect 25502 17847 25558 17856
rect 25410 17776 25466 17785
rect 25410 17711 25466 17720
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25608 17338 25636 17682
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25148 16697 25176 16730
rect 25134 16688 25190 16697
rect 25134 16623 25190 16632
rect 25044 16108 25096 16114
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 23938 15192 23994 15201
rect 24044 15162 24072 15506
rect 23938 15127 23994 15136
rect 24032 15156 24084 15162
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23768 12442 23796 14758
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23860 14074 23888 14350
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23662 11792 23718 11801
rect 23662 11727 23718 11736
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23676 9178 23704 11494
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23400 8634 23520 8650
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23400 8628 23532 8634
rect 23400 8622 23480 8628
rect 23400 8022 23428 8622
rect 23480 8570 23532 8576
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 23400 7546 23428 7958
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23308 3738 23336 5646
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23492 4826 23520 5510
rect 23584 5166 23612 6054
rect 23572 5160 23624 5166
rect 23572 5102 23624 5108
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23570 4584 23626 4593
rect 23570 4519 23626 4528
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 23216 3194 23244 3606
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23204 2848 23256 2854
rect 23202 2816 23204 2825
rect 23256 2816 23258 2825
rect 23202 2751 23258 2760
rect 23584 2009 23612 4519
rect 23860 4162 23888 13466
rect 23952 11762 23980 15127
rect 24032 15098 24084 15104
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24044 13802 24072 14418
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23952 10606 23980 10950
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23938 9208 23994 9217
rect 24044 9178 24072 13738
rect 24228 13530 24256 16050
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24582 15056 24638 15065
rect 24582 14991 24638 15000
rect 24596 14958 24624 14991
rect 24584 14952 24636 14958
rect 24398 14920 24454 14929
rect 24584 14894 24636 14900
rect 24398 14855 24454 14864
rect 24412 14482 24440 14855
rect 24688 14634 24716 16102
rect 25044 16050 25096 16056
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24780 15910 24808 15943
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24766 15464 24822 15473
rect 24766 15399 24768 15408
rect 24820 15399 24822 15408
rect 24768 15370 24820 15376
rect 24766 14920 24822 14929
rect 24766 14855 24822 14864
rect 24780 14822 24808 14855
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24688 14618 24900 14634
rect 24688 14612 24912 14618
rect 24688 14606 24860 14612
rect 24860 14554 24912 14560
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 25608 14074 25636 14418
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 24674 13832 24730 13841
rect 24674 13767 24730 13776
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24582 13424 24638 13433
rect 24688 13410 24716 13767
rect 24766 13696 24822 13705
rect 24766 13631 24822 13640
rect 24780 13530 24808 13631
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24688 13382 24808 13410
rect 24582 13359 24584 13368
rect 24636 13359 24638 13368
rect 24584 13330 24636 13336
rect 24596 13172 24624 13330
rect 24596 13144 24716 13172
rect 24780 13161 24808 13382
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12986 24716 13144
rect 24766 13152 24822 13161
rect 24766 13087 24822 13096
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24582 12880 24638 12889
rect 24582 12815 24638 12824
rect 24596 12782 24624 12815
rect 24584 12776 24636 12782
rect 24584 12718 24636 12724
rect 24768 12640 24820 12646
rect 24766 12608 24768 12617
rect 24820 12608 24822 12617
rect 24766 12543 24822 12552
rect 24582 12336 24638 12345
rect 24582 12271 24584 12280
rect 24636 12271 24638 12280
rect 24584 12242 24636 12248
rect 24596 12186 24624 12242
rect 24596 12158 24716 12186
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11762 24256 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12158
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11937 24808 12038
rect 24766 11928 24822 11937
rect 24676 11892 24728 11898
rect 24766 11863 24822 11872
rect 24676 11834 24728 11840
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24228 10470 24256 11698
rect 24674 11384 24730 11393
rect 24674 11319 24730 11328
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24688 10305 24716 11319
rect 25320 11280 25372 11286
rect 25320 11222 25372 11228
rect 24766 11112 24822 11121
rect 24766 11047 24768 11056
rect 24820 11047 24822 11056
rect 24768 11018 24820 11024
rect 24766 10840 24822 10849
rect 24766 10775 24822 10784
rect 24674 10296 24730 10305
rect 24674 10231 24730 10240
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24780 9704 24808 10775
rect 25332 9926 25360 11222
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25424 11014 25452 11086
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10810 25452 10950
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25608 10470 25636 11154
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 24688 9676 24808 9704
rect 24688 9489 24716 9676
rect 24872 9602 24900 9862
rect 24780 9574 24900 9602
rect 24780 9518 24808 9574
rect 24768 9512 24820 9518
rect 24674 9480 24730 9489
rect 24768 9454 24820 9460
rect 24674 9415 24730 9424
rect 24122 9344 24178 9353
rect 24122 9279 24178 9288
rect 23938 9143 23994 9152
rect 24032 9172 24084 9178
rect 23952 7313 23980 9143
rect 24032 9114 24084 9120
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23938 7304 23994 7313
rect 23938 7239 23994 7248
rect 24044 6458 24072 8366
rect 24136 7698 24164 9279
rect 24780 9110 24808 9454
rect 24768 9104 24820 9110
rect 24214 9072 24270 9081
rect 24768 9046 24820 9052
rect 24214 9007 24270 9016
rect 24860 9036 24912 9042
rect 24228 7857 24256 9007
rect 24860 8978 24912 8984
rect 24676 8968 24728 8974
rect 24674 8936 24676 8945
rect 24768 8968 24820 8974
rect 24728 8936 24730 8945
rect 24768 8910 24820 8916
rect 24674 8871 24730 8880
rect 24780 8838 24808 8910
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24780 8634 24808 8774
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24584 8356 24636 8362
rect 24584 8298 24636 8304
rect 24596 8090 24624 8298
rect 24780 8242 24808 8570
rect 24872 8537 24900 8978
rect 24858 8528 24914 8537
rect 24858 8463 24914 8472
rect 24872 8430 24900 8463
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24780 8214 24900 8242
rect 24872 8090 24900 8214
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24214 7848 24270 7857
rect 24214 7783 24270 7792
rect 24674 7848 24730 7857
rect 24674 7783 24730 7792
rect 24136 7670 24256 7698
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24136 7002 24164 7346
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24122 6352 24178 6361
rect 24122 6287 24178 6296
rect 23860 4134 23980 4162
rect 23754 4040 23810 4049
rect 23754 3975 23810 3984
rect 23848 4004 23900 4010
rect 23768 3738 23796 3975
rect 23848 3946 23900 3952
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23662 3360 23718 3369
rect 23662 3295 23718 3304
rect 23676 2689 23704 3295
rect 23768 3194 23796 3674
rect 23860 3466 23888 3946
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23662 2680 23718 2689
rect 23860 2650 23888 3402
rect 23952 3233 23980 4134
rect 24136 3913 24164 6287
rect 24122 3904 24178 3913
rect 24122 3839 24178 3848
rect 24122 3496 24178 3505
rect 24122 3431 24178 3440
rect 23938 3224 23994 3233
rect 23938 3159 23994 3168
rect 23662 2615 23718 2624
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23952 2514 23980 3159
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23570 2000 23626 2009
rect 23570 1935 23626 1944
rect 22928 604 22980 610
rect 22928 546 22980 552
rect 23480 604 23532 610
rect 23480 546 23532 552
rect 23492 480 23520 546
rect 24136 480 24164 3431
rect 24228 3097 24256 7670
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7206 24716 7783
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 25226 6896 25282 6905
rect 25226 6831 25228 6840
rect 25280 6831 25282 6840
rect 25228 6802 25280 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 25240 6458 25268 6802
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 24492 6384 24544 6390
rect 25332 6361 25360 9862
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25516 8362 25544 9318
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25608 7857 25636 10406
rect 25594 7848 25650 7857
rect 25594 7783 25650 7792
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 24492 6326 24544 6332
rect 25318 6352 25374 6361
rect 24504 6118 24532 6326
rect 24676 6316 24728 6322
rect 25318 6287 25374 6296
rect 24676 6258 24728 6264
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24688 5710 24716 6258
rect 25136 6180 25188 6186
rect 25136 6122 25188 6128
rect 25148 5914 25176 6122
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24688 5574 24716 5646
rect 24676 5568 24728 5574
rect 24676 5510 24728 5516
rect 24766 5536 24822 5545
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5098 24716 5510
rect 24766 5471 24822 5480
rect 24676 5092 24728 5098
rect 24676 5034 24728 5040
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 5034
rect 24780 5030 24808 5471
rect 24872 5370 24900 5714
rect 25424 5681 25452 6598
rect 25410 5672 25466 5681
rect 25410 5607 25466 5616
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24780 3466 24808 4422
rect 24872 3738 24900 5306
rect 25226 4448 25282 4457
rect 25226 4383 25282 4392
rect 25240 3777 25268 4383
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25226 3768 25282 3777
rect 24860 3732 24912 3738
rect 25332 3738 25360 3975
rect 25226 3703 25228 3712
rect 24860 3674 24912 3680
rect 25280 3703 25282 3712
rect 25320 3732 25372 3738
rect 25228 3674 25280 3680
rect 25320 3674 25372 3680
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24214 3088 24270 3097
rect 25240 3058 25268 3674
rect 25332 3194 25360 3674
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25516 3194 25544 3470
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 24214 3023 24270 3032
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 24766 2952 24822 2961
rect 24766 2887 24822 2896
rect 24780 2854 24808 2887
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 24676 2372 24728 2378
rect 24676 2314 24728 2320
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1170 24716 2314
rect 24688 1142 24808 1170
rect 24780 480 24808 1142
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2318 0 2374 480
rect 2962 0 3018 480
rect 3698 0 3754 480
rect 4342 0 4398 480
rect 4986 0 5042 480
rect 5722 0 5778 480
rect 6366 0 6422 480
rect 7102 0 7158 480
rect 7746 0 7802 480
rect 8390 0 8446 480
rect 9126 0 9182 480
rect 9770 0 9826 480
rect 10506 0 10562 480
rect 11150 0 11206 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15290 0 15346 480
rect 15934 0 15990 480
rect 16578 0 16634 480
rect 17314 0 17370 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19338 0 19394 480
rect 20074 0 20130 480
rect 20718 0 20774 480
rect 21362 0 21418 480
rect 22098 0 22154 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25332 377 25360 3130
rect 27526 2952 27582 2961
rect 27526 2887 27582 2896
rect 25502 2816 25558 2825
rect 25502 2751 25558 2760
rect 25516 480 25544 2751
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 26160 480 26188 2314
rect 26790 1456 26846 1465
rect 26846 1414 26924 1442
rect 26790 1391 26846 1400
rect 26896 480 26924 1414
rect 27540 480 27568 2887
rect 25318 368 25374 377
rect 25318 303 25374 312
rect 25502 0 25558 480
rect 26146 0 26202 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 23294 27648 23350 27704
rect 1582 24656 1638 24712
rect 1490 22616 1546 22672
rect 1582 20868 1638 20904
rect 1582 20848 1584 20868
rect 1584 20848 1636 20868
rect 1636 20848 1638 20868
rect 1582 20304 1638 20360
rect 386 16224 442 16280
rect 938 3440 994 3496
rect 294 3304 350 3360
rect 1674 13912 1730 13968
rect 1490 10548 1492 10568
rect 1492 10548 1544 10568
rect 1544 10548 1546 10568
rect 1490 10512 1546 10548
rect 2962 24248 3018 24304
rect 4342 24520 4398 24576
rect 4986 23568 5042 23624
rect 3698 22344 3754 22400
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5538 21936 5594 21992
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6366 21392 6422 21448
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10138 24520 10194 24576
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9770 24112 9826 24168
rect 9126 20712 9182 20768
rect 7746 19896 7802 19952
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10782 23160 10838 23216
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10598 21936 10654 21992
rect 11058 21392 11114 21448
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10782 20440 10838 20496
rect 10966 20204 10968 20224
rect 10968 20204 11020 20224
rect 11020 20204 11022 20224
rect 10966 20168 11022 20204
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 11794 24248 11850 24304
rect 11426 23860 11482 23896
rect 11426 23840 11428 23860
rect 11428 23840 11480 23860
rect 11480 23840 11482 23860
rect 11334 23432 11390 23488
rect 12070 23568 12126 23624
rect 11886 23296 11942 23352
rect 11150 19352 11206 19408
rect 7102 19216 7158 19272
rect 10874 19216 10930 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10874 17620 10876 17640
rect 10876 17620 10928 17640
rect 10928 17620 10930 17640
rect 10874 17584 10930 17620
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 8206 14320 8262 14376
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 2318 13096 2374 13152
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 4986 11056 5042 11112
rect 2870 10512 2926 10568
rect 4342 10512 4398 10568
rect 2778 9560 2834 9616
rect 2870 9288 2926 9344
rect 2318 6296 2374 6352
rect 1950 3440 2006 3496
rect 3698 6704 3754 6760
rect 2870 4664 2926 4720
rect 4066 2372 4122 2408
rect 4066 2352 4068 2372
rect 4068 2352 4120 2372
rect 4120 2352 4122 2372
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6366 7384 6422 7440
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5998 5480 6054 5536
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 11150 17584 11206 17640
rect 11426 17040 11482 17096
rect 10966 14048 11022 14104
rect 11058 13640 11114 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 8390 13232 8446 13288
rect 7102 3984 7158 4040
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9954 9560 10010 9616
rect 9678 9324 9680 9344
rect 9680 9324 9732 9344
rect 9732 9324 9734 9344
rect 9678 9288 9734 9324
rect 9126 9016 9182 9072
rect 9034 6160 9090 6216
rect 9034 2352 9090 2408
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10874 7656 10930 7712
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 9770 5072 9826 5128
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10782 4528 10838 4584
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10506 1400 10562 1456
rect 12070 13776 12126 13832
rect 11886 12416 11942 12472
rect 11242 8472 11298 8528
rect 11150 6840 11206 6896
rect 11794 6296 11850 6352
rect 11702 4120 11758 4176
rect 11242 3984 11298 4040
rect 11426 2796 11428 2816
rect 11428 2796 11480 2816
rect 11480 2796 11482 2816
rect 11426 2760 11482 2796
rect 11610 1536 11666 1592
rect 12806 24112 12862 24168
rect 12530 21800 12586 21856
rect 12438 20032 12494 20088
rect 12346 19896 12402 19952
rect 13358 24792 13414 24848
rect 12898 23432 12954 23488
rect 12806 21120 12862 21176
rect 12898 20460 12954 20496
rect 12898 20440 12900 20460
rect 12900 20440 12952 20460
rect 12952 20440 12954 20460
rect 12806 19352 12862 19408
rect 12898 19116 12900 19136
rect 12900 19116 12952 19136
rect 12952 19116 12954 19136
rect 12898 19080 12954 19116
rect 12806 18028 12808 18048
rect 12808 18028 12860 18048
rect 12860 18028 12862 18048
rect 12806 17992 12862 18028
rect 12990 16496 13046 16552
rect 12714 13368 12770 13424
rect 12714 12688 12770 12744
rect 12346 12552 12402 12608
rect 12346 11056 12402 11112
rect 12162 9016 12218 9072
rect 12438 9288 12494 9344
rect 11978 7964 11980 7984
rect 11980 7964 12032 7984
rect 12032 7964 12034 7984
rect 11978 7928 12034 7964
rect 12438 8064 12494 8120
rect 12530 7828 12532 7848
rect 12532 7828 12584 7848
rect 12584 7828 12586 7848
rect 12530 7792 12586 7828
rect 12438 7384 12494 7440
rect 12622 7112 12678 7168
rect 12254 6060 12256 6080
rect 12256 6060 12308 6080
rect 12308 6060 12310 6080
rect 12254 6024 12310 6060
rect 12438 3848 12494 3904
rect 12254 3440 12310 3496
rect 12438 2524 12440 2544
rect 12440 2524 12492 2544
rect 12492 2524 12494 2544
rect 12438 2488 12494 2524
rect 13634 23024 13690 23080
rect 13266 20440 13322 20496
rect 13358 19080 13414 19136
rect 13266 18148 13322 18184
rect 13266 18128 13268 18148
rect 13268 18128 13320 18148
rect 13320 18128 13322 18148
rect 12990 13776 13046 13832
rect 13266 13776 13322 13832
rect 13266 11600 13322 11656
rect 13818 20712 13874 20768
rect 14186 23060 14188 23080
rect 14188 23060 14240 23080
rect 14240 23060 14242 23080
rect 14186 23024 14242 23060
rect 14094 22072 14150 22128
rect 14094 19896 14150 19952
rect 14094 19760 14150 19816
rect 13450 16360 13506 16416
rect 13726 15000 13782 15056
rect 13634 14320 13690 14376
rect 14462 24556 14464 24576
rect 14464 24556 14516 24576
rect 14516 24556 14518 24576
rect 14462 24520 14518 24556
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15290 24792 15346 24848
rect 15198 24676 15254 24712
rect 15198 24656 15200 24676
rect 15200 24656 15252 24676
rect 15252 24656 15254 24676
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14554 23840 14610 23896
rect 14462 23568 14518 23624
rect 14370 20032 14426 20088
rect 14278 17176 14334 17232
rect 14370 16632 14426 16688
rect 14186 14456 14242 14512
rect 14278 14340 14334 14376
rect 14278 14320 14280 14340
rect 14280 14320 14332 14340
rect 14332 14320 14334 14340
rect 14278 14048 14334 14104
rect 14002 13504 14058 13560
rect 13818 12824 13874 12880
rect 13542 10512 13598 10568
rect 13358 10376 13414 10432
rect 13358 9288 13414 9344
rect 12990 8200 13046 8256
rect 12990 7928 13046 7984
rect 12806 7268 12862 7304
rect 12806 7248 12808 7268
rect 12808 7248 12860 7268
rect 12860 7248 12862 7268
rect 13450 8336 13506 8392
rect 13358 7384 13414 7440
rect 15474 23296 15530 23352
rect 13910 11464 13966 11520
rect 13542 7656 13598 7712
rect 13450 6704 13506 6760
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15382 22380 15384 22400
rect 15384 22380 15436 22400
rect 15436 22380 15438 22400
rect 15382 22344 15438 22380
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15290 21428 15292 21448
rect 15292 21428 15344 21448
rect 15344 21428 15346 21448
rect 15290 21392 15346 21428
rect 15474 20984 15530 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15382 20576 15438 20632
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14830 19352 14886 19408
rect 15750 23724 15806 23760
rect 15750 23704 15752 23724
rect 15752 23704 15804 23724
rect 15804 23704 15806 23724
rect 15934 21800 15990 21856
rect 15658 20168 15714 20224
rect 15566 19624 15622 19680
rect 14830 18672 14886 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15106 16088 15162 16144
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14830 13912 14886 13968
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14462 10668 14518 10704
rect 14462 10648 14464 10668
rect 14464 10648 14516 10668
rect 14516 10648 14518 10668
rect 14186 10240 14242 10296
rect 14094 10004 14096 10024
rect 14096 10004 14148 10024
rect 14148 10004 14150 10024
rect 14094 9968 14150 10004
rect 14002 7948 14058 7984
rect 14002 7928 14004 7948
rect 14004 7928 14056 7948
rect 14056 7928 14058 7948
rect 13634 6704 13690 6760
rect 13358 5888 13414 5944
rect 14186 8200 14242 8256
rect 13634 6024 13690 6080
rect 13542 3032 13598 3088
rect 13634 2896 13690 2952
rect 14278 3576 14334 3632
rect 13634 2352 13690 2408
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15842 20440 15898 20496
rect 15750 17992 15806 18048
rect 15658 17448 15714 17504
rect 15658 15136 15714 15192
rect 15566 13232 15622 13288
rect 16026 16496 16082 16552
rect 15382 11464 15438 11520
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15014 9288 15070 9344
rect 15658 9832 15714 9888
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15198 6840 15254 6896
rect 15290 6704 15346 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15658 5788 15660 5808
rect 15660 5788 15712 5808
rect 15712 5788 15714 5808
rect 15658 5752 15714 5788
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15750 5344 15806 5400
rect 16578 24520 16634 24576
rect 16486 23160 16542 23216
rect 16486 22616 16542 22672
rect 16302 20440 16358 20496
rect 16670 20204 16672 20224
rect 16672 20204 16724 20224
rect 16724 20204 16726 20224
rect 16670 20168 16726 20204
rect 16210 15544 16266 15600
rect 16486 13776 16542 13832
rect 16302 13096 16358 13152
rect 16486 13368 16542 13424
rect 16394 12552 16450 12608
rect 16302 12416 16358 12472
rect 17038 23860 17094 23896
rect 17038 23840 17040 23860
rect 17040 23840 17092 23860
rect 17092 23840 17094 23860
rect 17038 23432 17094 23488
rect 17314 22480 17370 22536
rect 17222 19216 17278 19272
rect 16670 10648 16726 10704
rect 17222 14864 17278 14920
rect 17130 12416 17186 12472
rect 17222 11736 17278 11792
rect 17038 10648 17094 10704
rect 16762 9832 16818 9888
rect 16670 9288 16726 9344
rect 16578 7812 16634 7848
rect 16578 7792 16580 7812
rect 16580 7792 16632 7812
rect 16632 7792 16634 7812
rect 16394 6876 16396 6896
rect 16396 6876 16448 6896
rect 16448 6876 16450 6896
rect 16394 6840 16450 6876
rect 15106 5208 15162 5264
rect 15842 5208 15898 5264
rect 14738 4664 14794 4720
rect 15382 4664 15438 4720
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14830 4120 14886 4176
rect 15106 3732 15162 3768
rect 15106 3712 15108 3732
rect 15108 3712 15160 3732
rect 15160 3712 15162 3732
rect 15934 3884 15936 3904
rect 15936 3884 15988 3904
rect 15988 3884 15990 3904
rect 15934 3848 15990 3884
rect 15382 3440 15438 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15290 2760 15346 2816
rect 13358 1672 13414 1728
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14462 1808 14518 1864
rect 14554 1400 14610 1456
rect 15566 3168 15622 3224
rect 15474 2796 15476 2816
rect 15476 2796 15528 2816
rect 15528 2796 15530 2816
rect 15474 2760 15530 2796
rect 15934 2508 15990 2544
rect 16302 5616 16358 5672
rect 16394 4800 16450 4856
rect 16854 8200 16910 8256
rect 16854 6160 16910 6216
rect 16762 5344 16818 5400
rect 16854 5208 16910 5264
rect 16670 5072 16726 5128
rect 16302 4528 16358 4584
rect 16946 4256 17002 4312
rect 15934 2488 15936 2508
rect 15936 2488 15988 2508
rect 15988 2488 15990 2508
rect 16210 2488 16266 2544
rect 16578 3032 16634 3088
rect 16762 3068 16764 3088
rect 16764 3068 16816 3088
rect 16816 3068 16818 3088
rect 16762 3032 16818 3068
rect 16394 2388 16396 2408
rect 16396 2388 16448 2408
rect 16448 2388 16450 2408
rect 16394 2352 16450 2388
rect 15934 1536 15990 1592
rect 17406 17332 17462 17368
rect 17406 17312 17408 17332
rect 17408 17312 17460 17332
rect 17460 17312 17462 17332
rect 17406 14184 17462 14240
rect 17774 23568 17830 23624
rect 18510 23568 18566 23624
rect 17682 21120 17738 21176
rect 17682 18944 17738 19000
rect 17866 18944 17922 19000
rect 17774 16224 17830 16280
rect 17774 13640 17830 13696
rect 17498 12436 17554 12472
rect 17498 12416 17500 12436
rect 17500 12416 17552 12436
rect 17552 12416 17554 12436
rect 18050 17584 18106 17640
rect 18694 23432 18750 23488
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20074 24792 20130 24848
rect 19338 23840 19394 23896
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19246 22616 19302 22672
rect 19246 22344 19302 22400
rect 19154 21392 19210 21448
rect 18694 19372 18750 19408
rect 18694 19352 18696 19372
rect 18696 19352 18748 19372
rect 18748 19352 18750 19372
rect 18326 19080 18382 19136
rect 18234 15544 18290 15600
rect 17958 14456 18014 14512
rect 18602 14456 18658 14512
rect 18418 10240 18474 10296
rect 17314 5888 17370 5944
rect 17222 3440 17278 3496
rect 17866 9444 17922 9480
rect 17866 9424 17868 9444
rect 17868 9424 17920 9444
rect 17920 9424 17922 9444
rect 18510 9560 18566 9616
rect 17958 8356 18014 8392
rect 17958 8336 17960 8356
rect 17960 8336 18012 8356
rect 18012 8336 18014 8356
rect 18142 8336 18198 8392
rect 18050 8064 18106 8120
rect 18142 7928 18198 7984
rect 17498 4392 17554 4448
rect 17774 4972 17776 4992
rect 17776 4972 17828 4992
rect 17828 4972 17830 4992
rect 17774 4936 17830 4972
rect 19246 18128 19302 18184
rect 19062 15952 19118 16008
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19430 18944 19486 19000
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19798 18828 19854 18864
rect 19798 18808 19800 18828
rect 19800 18808 19852 18828
rect 19852 18808 19854 18828
rect 19982 18264 20038 18320
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20074 17876 20130 17912
rect 20074 17856 20076 17876
rect 20076 17856 20128 17876
rect 20128 17856 20130 17876
rect 19798 17584 19854 17640
rect 19338 17040 19394 17096
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 18786 12724 18788 12744
rect 18788 12724 18840 12744
rect 18840 12724 18842 12744
rect 18786 12688 18842 12724
rect 19246 14184 19302 14240
rect 19430 13504 19486 13560
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19062 12688 19118 12744
rect 21914 27104 21970 27160
rect 21362 24792 21418 24848
rect 21454 24404 21510 24440
rect 21454 24384 21456 24404
rect 21456 24384 21508 24404
rect 21508 24384 21510 24404
rect 20626 23704 20682 23760
rect 21362 23568 21418 23624
rect 20350 22344 20406 22400
rect 20350 19760 20406 19816
rect 20902 23044 20958 23080
rect 20902 23024 20904 23044
rect 20904 23024 20956 23044
rect 20956 23024 20958 23044
rect 21362 22480 21418 22536
rect 21086 20576 21142 20632
rect 20442 19352 20498 19408
rect 20350 18808 20406 18864
rect 20258 17720 20314 17776
rect 20350 17584 20406 17640
rect 20442 17448 20498 17504
rect 20166 12960 20222 13016
rect 18970 11872 19026 11928
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18786 9424 18842 9480
rect 18510 7792 18566 7848
rect 18510 6840 18566 6896
rect 18418 6704 18474 6760
rect 17682 4120 17738 4176
rect 18418 4120 18474 4176
rect 18142 3712 18198 3768
rect 17774 3576 17830 3632
rect 17958 2896 18014 2952
rect 17222 2252 17224 2272
rect 17224 2252 17276 2272
rect 17276 2252 17278 2272
rect 17222 2216 17278 2252
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19246 11192 19302 11248
rect 19522 11056 19578 11112
rect 20074 12008 20130 12064
rect 19430 10240 19486 10296
rect 19154 6704 19210 6760
rect 19062 6432 19118 6488
rect 19338 7112 19394 7168
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19982 7792 20038 7848
rect 19706 7248 19762 7304
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19338 5208 19394 5264
rect 18786 4664 18842 4720
rect 18694 4256 18750 4312
rect 18510 3304 18566 3360
rect 18326 2372 18382 2408
rect 18326 2352 18328 2372
rect 18328 2352 18380 2372
rect 18380 2352 18382 2372
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19522 4392 19578 4448
rect 19890 4392 19946 4448
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19338 3440 19394 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20718 17196 20774 17232
rect 20718 17176 20720 17196
rect 20720 17176 20772 17196
rect 20772 17176 20774 17196
rect 20902 19896 20958 19952
rect 21362 20848 21418 20904
rect 21362 19760 21418 19816
rect 21178 18164 21180 18184
rect 21180 18164 21232 18184
rect 21232 18164 21234 18184
rect 21178 18128 21234 18164
rect 20994 17720 21050 17776
rect 21270 16360 21326 16416
rect 21546 19216 21602 19272
rect 21454 15952 21510 16008
rect 20902 13948 20904 13968
rect 20904 13948 20956 13968
rect 20956 13948 20958 13968
rect 20902 13912 20958 13948
rect 21086 13776 21142 13832
rect 20442 11600 20498 11656
rect 20626 11192 20682 11248
rect 21914 18128 21970 18184
rect 21914 14476 21970 14512
rect 21914 14456 21916 14476
rect 21916 14456 21968 14476
rect 21968 14456 21970 14476
rect 21546 11056 21602 11112
rect 21270 10512 21326 10568
rect 21362 10240 21418 10296
rect 21362 10004 21364 10024
rect 21364 10004 21416 10024
rect 21416 10004 21418 10024
rect 21362 9968 21418 10004
rect 20810 9288 20866 9344
rect 21086 9152 21142 9208
rect 21086 8880 21142 8936
rect 20994 8336 21050 8392
rect 20718 5616 20774 5672
rect 22558 24792 22614 24848
rect 22374 24656 22430 24712
rect 22374 22344 22430 22400
rect 23018 23160 23074 23216
rect 23386 26560 23442 26616
rect 23570 25336 23626 25392
rect 24674 25880 24730 25936
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24792 24822 24848
rect 25318 24792 25374 24848
rect 24122 24656 24178 24712
rect 23478 24384 23534 24440
rect 23570 24112 23626 24168
rect 23478 23568 23534 23624
rect 23294 22380 23296 22400
rect 23296 22380 23348 22400
rect 23348 22380 23350 22400
rect 23294 22344 23350 22380
rect 22650 19352 22706 19408
rect 22098 12724 22100 12744
rect 22100 12724 22152 12744
rect 22152 12724 22154 12744
rect 22098 12688 22154 12724
rect 22558 13096 22614 13152
rect 22282 12980 22338 13016
rect 22282 12960 22284 12980
rect 22284 12960 22336 12980
rect 22336 12960 22338 12980
rect 22190 12280 22246 12336
rect 22466 12044 22468 12064
rect 22468 12044 22520 12064
rect 22520 12044 22522 12064
rect 22466 12008 22522 12044
rect 21914 8508 21916 8528
rect 21916 8508 21968 8528
rect 21968 8508 21970 8528
rect 21914 8472 21970 8508
rect 21270 7384 21326 7440
rect 20994 3984 21050 4040
rect 20902 3712 20958 3768
rect 20994 3576 21050 3632
rect 20718 3168 20774 3224
rect 19430 1672 19486 1728
rect 19338 1536 19394 1592
rect 21362 6432 21418 6488
rect 21178 4936 21234 4992
rect 21362 4120 21418 4176
rect 21638 6332 21640 6352
rect 21640 6332 21692 6352
rect 21692 6332 21694 6352
rect 21638 6296 21694 6332
rect 22098 6876 22100 6896
rect 22100 6876 22152 6896
rect 22152 6876 22154 6896
rect 22098 6840 22154 6876
rect 22742 11892 22798 11928
rect 22742 11872 22744 11892
rect 22744 11872 22796 11892
rect 22796 11872 22798 11892
rect 23202 18672 23258 18728
rect 23754 24520 23810 24576
rect 24766 24404 24822 24440
rect 24766 24384 24768 24404
rect 24768 24384 24820 24404
rect 24820 24384 24822 24404
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23860 24822 23896
rect 24766 23840 24768 23860
rect 24768 23840 24820 23860
rect 24820 23840 24822 23860
rect 23570 22616 23626 22672
rect 23478 21800 23534 21856
rect 24766 23432 24822 23488
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23662 21256 23718 21312
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 23754 20984 23810 21040
rect 23662 19896 23718 19952
rect 23202 17604 23258 17640
rect 23202 17584 23204 17604
rect 23204 17584 23256 17604
rect 23256 17584 23258 17604
rect 23202 17312 23258 17368
rect 23938 18808 23994 18864
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 21800 24822 21856
rect 24766 20304 24822 20360
rect 24950 20712 25006 20768
rect 25502 24520 25558 24576
rect 26882 24384 26938 24440
rect 27526 23840 27582 23896
rect 26146 23432 26202 23488
rect 25410 23024 25466 23080
rect 24766 18944 24822 19000
rect 24030 17720 24086 17776
rect 23202 16360 23258 16416
rect 23202 10648 23258 10704
rect 21730 5208 21786 5264
rect 21546 4120 21602 4176
rect 21546 3984 21602 4040
rect 21546 2896 21602 2952
rect 22558 5616 22614 5672
rect 22282 4428 22284 4448
rect 22284 4428 22336 4448
rect 22336 4428 22338 4448
rect 22282 4392 22338 4428
rect 22098 3576 22154 3632
rect 22282 3440 22338 3496
rect 22834 5480 22890 5536
rect 21362 1808 21418 1864
rect 21270 856 21326 912
rect 21914 1400 21970 1456
rect 22834 2508 22890 2544
rect 22834 2488 22836 2508
rect 22836 2488 22888 2508
rect 22888 2488 22890 2508
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24030 16632 24086 16688
rect 24122 16224 24178 16280
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24858 18128 24914 18184
rect 24950 17176 25006 17232
rect 25226 18264 25282 18320
rect 25686 18400 25742 18456
rect 25502 17856 25558 17912
rect 25410 17720 25466 17776
rect 25134 16632 25190 16688
rect 23938 15136 23994 15192
rect 23662 11736 23718 11792
rect 23570 4528 23626 4584
rect 23202 2796 23204 2816
rect 23204 2796 23256 2816
rect 23256 2796 23258 2816
rect 23202 2760 23258 2796
rect 23938 9152 23994 9208
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24582 15000 24638 15056
rect 24398 14864 24454 14920
rect 24766 15952 24822 16008
rect 24766 15428 24822 15464
rect 24766 15408 24768 15428
rect 24768 15408 24820 15428
rect 24820 15408 24822 15428
rect 24766 14864 24822 14920
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24674 13776 24730 13832
rect 24582 13388 24638 13424
rect 24582 13368 24584 13388
rect 24584 13368 24636 13388
rect 24636 13368 24638 13388
rect 24766 13640 24822 13696
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24766 13096 24822 13152
rect 24582 12824 24638 12880
rect 24766 12588 24768 12608
rect 24768 12588 24820 12608
rect 24820 12588 24822 12608
rect 24766 12552 24822 12588
rect 24582 12300 24638 12336
rect 24582 12280 24584 12300
rect 24584 12280 24636 12300
rect 24636 12280 24638 12300
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11872 24822 11928
rect 24674 11328 24730 11384
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24766 11076 24822 11112
rect 24766 11056 24768 11076
rect 24768 11056 24820 11076
rect 24820 11056 24822 11076
rect 24766 10784 24822 10840
rect 24674 10240 24730 10296
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9424 24730 9480
rect 24122 9288 24178 9344
rect 23938 7248 23994 7304
rect 24214 9016 24270 9072
rect 24674 8916 24676 8936
rect 24676 8916 24728 8936
rect 24728 8916 24730 8936
rect 24674 8880 24730 8916
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24858 8472 24914 8528
rect 24214 7792 24270 7848
rect 24674 7792 24730 7848
rect 24122 6296 24178 6352
rect 23754 3984 23810 4040
rect 23662 3304 23718 3360
rect 23662 2624 23718 2680
rect 24122 3848 24178 3904
rect 24122 3440 24178 3496
rect 23938 3168 23994 3224
rect 23570 1944 23626 2000
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 25226 6860 25282 6896
rect 25226 6840 25228 6860
rect 25228 6840 25280 6860
rect 25280 6840 25282 6860
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25594 7792 25650 7848
rect 25318 6296 25374 6352
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24766 5480 24822 5536
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25410 5616 25466 5672
rect 25226 4392 25282 4448
rect 25318 3984 25374 4040
rect 25226 3732 25282 3768
rect 25226 3712 25228 3732
rect 25228 3712 25280 3732
rect 25280 3712 25282 3732
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24214 3032 24270 3088
rect 24766 2896 24822 2952
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27526 2896 27582 2952
rect 25502 2760 25558 2816
rect 26790 1400 26846 1456
rect 25318 312 25374 368
<< metal3 >>
rect 23289 27706 23355 27709
rect 27520 27706 28000 27736
rect 23289 27704 28000 27706
rect 23289 27648 23294 27704
rect 23350 27648 28000 27704
rect 23289 27646 28000 27648
rect 23289 27643 23355 27646
rect 27520 27616 28000 27646
rect 21909 27162 21975 27165
rect 27520 27162 28000 27192
rect 21909 27160 28000 27162
rect 21909 27104 21914 27160
rect 21970 27104 28000 27160
rect 21909 27102 28000 27104
rect 21909 27099 21975 27102
rect 27520 27072 28000 27102
rect 23381 26618 23447 26621
rect 27520 26618 28000 26648
rect 23381 26616 28000 26618
rect 23381 26560 23386 26616
rect 23442 26560 28000 26616
rect 23381 26558 28000 26560
rect 23381 26555 23447 26558
rect 27520 26528 28000 26558
rect 24669 25938 24735 25941
rect 27520 25938 28000 25968
rect 24669 25936 28000 25938
rect 24669 25880 24674 25936
rect 24730 25880 28000 25936
rect 24669 25878 28000 25880
rect 24669 25875 24735 25878
rect 27520 25848 28000 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 23565 25394 23631 25397
rect 27520 25394 28000 25424
rect 23565 25392 28000 25394
rect 23565 25336 23570 25392
rect 23626 25336 28000 25392
rect 23565 25334 28000 25336
rect 23565 25331 23631 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 13353 24850 13419 24853
rect 15285 24850 15351 24853
rect 13353 24848 15351 24850
rect 13353 24792 13358 24848
rect 13414 24792 15290 24848
rect 15346 24792 15351 24848
rect 13353 24790 15351 24792
rect 13353 24787 13419 24790
rect 15285 24787 15351 24790
rect 20069 24850 20135 24853
rect 21357 24850 21423 24853
rect 20069 24848 21423 24850
rect 20069 24792 20074 24848
rect 20130 24792 21362 24848
rect 21418 24792 21423 24848
rect 20069 24790 21423 24792
rect 20069 24787 20135 24790
rect 21357 24787 21423 24790
rect 22553 24850 22619 24853
rect 24761 24850 24827 24853
rect 22553 24848 24827 24850
rect 22553 24792 22558 24848
rect 22614 24792 24766 24848
rect 24822 24792 24827 24848
rect 22553 24790 24827 24792
rect 22553 24787 22619 24790
rect 24761 24787 24827 24790
rect 25313 24850 25379 24853
rect 27520 24850 28000 24880
rect 25313 24848 28000 24850
rect 25313 24792 25318 24848
rect 25374 24792 28000 24848
rect 25313 24790 28000 24792
rect 25313 24787 25379 24790
rect 27520 24760 28000 24790
rect 1577 24714 1643 24717
rect 15193 24714 15259 24717
rect 1577 24712 15259 24714
rect 1577 24656 1582 24712
rect 1638 24656 15198 24712
rect 15254 24656 15259 24712
rect 1577 24654 15259 24656
rect 1577 24651 1643 24654
rect 15193 24651 15259 24654
rect 22369 24714 22435 24717
rect 24117 24714 24183 24717
rect 22369 24712 24183 24714
rect 22369 24656 22374 24712
rect 22430 24656 24122 24712
rect 24178 24656 24183 24712
rect 22369 24654 24183 24656
rect 22369 24651 22435 24654
rect 24117 24651 24183 24654
rect 4337 24578 4403 24581
rect 10133 24578 10199 24581
rect 4337 24576 10199 24578
rect 4337 24520 4342 24576
rect 4398 24520 10138 24576
rect 10194 24520 10199 24576
rect 4337 24518 10199 24520
rect 4337 24515 4403 24518
rect 10133 24515 10199 24518
rect 14457 24578 14523 24581
rect 16573 24578 16639 24581
rect 14457 24576 16639 24578
rect 14457 24520 14462 24576
rect 14518 24520 16578 24576
rect 16634 24520 16639 24576
rect 14457 24518 16639 24520
rect 14457 24515 14523 24518
rect 16573 24515 16639 24518
rect 23749 24578 23815 24581
rect 25497 24578 25563 24581
rect 23749 24576 25563 24578
rect 23749 24520 23754 24576
rect 23810 24520 25502 24576
rect 25558 24520 25563 24576
rect 23749 24518 25563 24520
rect 23749 24515 23815 24518
rect 25497 24515 25563 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 21449 24442 21515 24445
rect 23473 24442 23539 24445
rect 21449 24440 23539 24442
rect 21449 24384 21454 24440
rect 21510 24384 23478 24440
rect 23534 24384 23539 24440
rect 21449 24382 23539 24384
rect 21449 24379 21515 24382
rect 23473 24379 23539 24382
rect 24761 24442 24827 24445
rect 26877 24442 26943 24445
rect 24761 24440 26943 24442
rect 24761 24384 24766 24440
rect 24822 24384 26882 24440
rect 26938 24384 26943 24440
rect 24761 24382 26943 24384
rect 24761 24379 24827 24382
rect 26877 24379 26943 24382
rect 2957 24306 3023 24309
rect 11789 24306 11855 24309
rect 2957 24304 11855 24306
rect 2957 24248 2962 24304
rect 3018 24248 11794 24304
rect 11850 24248 11855 24304
rect 2957 24246 11855 24248
rect 2957 24243 3023 24246
rect 11789 24243 11855 24246
rect 9765 24170 9831 24173
rect 12801 24170 12867 24173
rect 9765 24168 12867 24170
rect 9765 24112 9770 24168
rect 9826 24112 12806 24168
rect 12862 24112 12867 24168
rect 9765 24110 12867 24112
rect 9765 24107 9831 24110
rect 12801 24107 12867 24110
rect 23565 24170 23631 24173
rect 27520 24170 28000 24200
rect 23565 24168 28000 24170
rect 23565 24112 23570 24168
rect 23626 24112 28000 24168
rect 23565 24110 28000 24112
rect 23565 24107 23631 24110
rect 27520 24080 28000 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 11421 23898 11487 23901
rect 14549 23898 14615 23901
rect 11421 23896 14615 23898
rect 11421 23840 11426 23896
rect 11482 23840 14554 23896
rect 14610 23840 14615 23896
rect 11421 23838 14615 23840
rect 11421 23835 11487 23838
rect 14549 23835 14615 23838
rect 17033 23898 17099 23901
rect 19333 23898 19399 23901
rect 17033 23896 19399 23898
rect 17033 23840 17038 23896
rect 17094 23840 19338 23896
rect 19394 23840 19399 23896
rect 17033 23838 19399 23840
rect 17033 23835 17099 23838
rect 19333 23835 19399 23838
rect 24761 23898 24827 23901
rect 27521 23898 27587 23901
rect 24761 23896 27587 23898
rect 24761 23840 24766 23896
rect 24822 23840 27526 23896
rect 27582 23840 27587 23896
rect 24761 23838 27587 23840
rect 24761 23835 24827 23838
rect 27521 23835 27587 23838
rect 15745 23762 15811 23765
rect 20621 23762 20687 23765
rect 15745 23760 20687 23762
rect 15745 23704 15750 23760
rect 15806 23704 20626 23760
rect 20682 23704 20687 23760
rect 15745 23702 20687 23704
rect 15745 23699 15811 23702
rect 20621 23699 20687 23702
rect 4981 23626 5047 23629
rect 12065 23626 12131 23629
rect 4981 23624 12131 23626
rect 4981 23568 4986 23624
rect 5042 23568 12070 23624
rect 12126 23568 12131 23624
rect 4981 23566 12131 23568
rect 4981 23563 5047 23566
rect 12065 23563 12131 23566
rect 14457 23626 14523 23629
rect 17769 23626 17835 23629
rect 14457 23624 17835 23626
rect 14457 23568 14462 23624
rect 14518 23568 17774 23624
rect 17830 23568 17835 23624
rect 14457 23566 17835 23568
rect 14457 23563 14523 23566
rect 17769 23563 17835 23566
rect 18505 23626 18571 23629
rect 21357 23626 21423 23629
rect 18505 23624 21423 23626
rect 18505 23568 18510 23624
rect 18566 23568 21362 23624
rect 21418 23568 21423 23624
rect 18505 23566 21423 23568
rect 18505 23563 18571 23566
rect 21357 23563 21423 23566
rect 23473 23626 23539 23629
rect 27520 23626 28000 23656
rect 23473 23624 28000 23626
rect 23473 23568 23478 23624
rect 23534 23568 28000 23624
rect 23473 23566 28000 23568
rect 23473 23563 23539 23566
rect 27520 23536 28000 23566
rect 11329 23490 11395 23493
rect 12893 23490 12959 23493
rect 11329 23488 12959 23490
rect 11329 23432 11334 23488
rect 11390 23432 12898 23488
rect 12954 23432 12959 23488
rect 11329 23430 12959 23432
rect 11329 23427 11395 23430
rect 12893 23427 12959 23430
rect 17033 23490 17099 23493
rect 18689 23490 18755 23493
rect 17033 23488 18755 23490
rect 17033 23432 17038 23488
rect 17094 23432 18694 23488
rect 18750 23432 18755 23488
rect 17033 23430 18755 23432
rect 17033 23427 17099 23430
rect 18689 23427 18755 23430
rect 24761 23490 24827 23493
rect 26141 23490 26207 23493
rect 24761 23488 26207 23490
rect 24761 23432 24766 23488
rect 24822 23432 26146 23488
rect 26202 23432 26207 23488
rect 24761 23430 26207 23432
rect 24761 23427 24827 23430
rect 26141 23427 26207 23430
rect 10277 23424 10597 23425
rect 0 23354 480 23384
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 11881 23354 11947 23357
rect 15469 23354 15535 23357
rect 0 23294 1226 23354
rect 0 23264 480 23294
rect 1166 22130 1226 23294
rect 11881 23352 15535 23354
rect 11881 23296 11886 23352
rect 11942 23296 15474 23352
rect 15530 23296 15535 23352
rect 11881 23294 15535 23296
rect 11881 23291 11947 23294
rect 15469 23291 15535 23294
rect 10777 23218 10843 23221
rect 16481 23218 16547 23221
rect 23013 23218 23079 23221
rect 10777 23216 23079 23218
rect 10777 23160 10782 23216
rect 10838 23160 16486 23216
rect 16542 23160 23018 23216
rect 23074 23160 23079 23216
rect 10777 23158 23079 23160
rect 10777 23155 10843 23158
rect 16481 23155 16547 23158
rect 23013 23155 23079 23158
rect 13629 23082 13695 23085
rect 14181 23082 14247 23085
rect 20897 23082 20963 23085
rect 13629 23080 20963 23082
rect 13629 23024 13634 23080
rect 13690 23024 14186 23080
rect 14242 23024 20902 23080
rect 20958 23024 20963 23080
rect 13629 23022 20963 23024
rect 13629 23019 13695 23022
rect 14181 23019 14247 23022
rect 20897 23019 20963 23022
rect 25405 23082 25471 23085
rect 27520 23082 28000 23112
rect 25405 23080 28000 23082
rect 25405 23024 25410 23080
rect 25466 23024 28000 23080
rect 25405 23022 28000 23024
rect 25405 23019 25471 23022
rect 27520 22992 28000 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1485 22674 1551 22677
rect 16481 22674 16547 22677
rect 1485 22672 16547 22674
rect 1485 22616 1490 22672
rect 1546 22616 16486 22672
rect 16542 22616 16547 22672
rect 1485 22614 16547 22616
rect 1485 22611 1551 22614
rect 16481 22611 16547 22614
rect 19241 22674 19307 22677
rect 23565 22674 23631 22677
rect 19241 22672 23631 22674
rect 19241 22616 19246 22672
rect 19302 22616 23570 22672
rect 23626 22616 23631 22672
rect 19241 22614 23631 22616
rect 19241 22611 19307 22614
rect 23565 22611 23631 22614
rect 17309 22538 17375 22541
rect 9998 22536 17375 22538
rect 9998 22480 17314 22536
rect 17370 22480 17375 22536
rect 9998 22478 17375 22480
rect 3693 22402 3759 22405
rect 9998 22402 10058 22478
rect 17309 22475 17375 22478
rect 21357 22538 21423 22541
rect 27520 22538 28000 22568
rect 21357 22536 28000 22538
rect 21357 22480 21362 22536
rect 21418 22480 28000 22536
rect 21357 22478 28000 22480
rect 21357 22475 21423 22478
rect 27520 22448 28000 22478
rect 3693 22400 10058 22402
rect 3693 22344 3698 22400
rect 3754 22344 10058 22400
rect 3693 22342 10058 22344
rect 15377 22402 15443 22405
rect 19241 22402 19307 22405
rect 15377 22400 19307 22402
rect 15377 22344 15382 22400
rect 15438 22344 19246 22400
rect 19302 22344 19307 22400
rect 15377 22342 19307 22344
rect 3693 22339 3759 22342
rect 15377 22339 15443 22342
rect 19241 22339 19307 22342
rect 20345 22402 20411 22405
rect 22369 22402 22435 22405
rect 23289 22402 23355 22405
rect 20345 22400 23355 22402
rect 20345 22344 20350 22400
rect 20406 22344 22374 22400
rect 22430 22344 23294 22400
rect 23350 22344 23355 22400
rect 20345 22342 23355 22344
rect 20345 22339 20411 22342
rect 22369 22339 22435 22342
rect 23289 22339 23355 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 14089 22130 14155 22133
rect 1166 22128 14155 22130
rect 1166 22072 14094 22128
rect 14150 22072 14155 22128
rect 1166 22070 14155 22072
rect 14089 22067 14155 22070
rect 5533 21994 5599 21997
rect 10593 21994 10659 21997
rect 5533 21992 10659 21994
rect 5533 21936 5538 21992
rect 5594 21936 10598 21992
rect 10654 21936 10659 21992
rect 5533 21934 10659 21936
rect 5533 21931 5599 21934
rect 10593 21931 10659 21934
rect 12525 21858 12591 21861
rect 14774 21858 14780 21860
rect 12525 21856 14780 21858
rect 12525 21800 12530 21856
rect 12586 21800 14780 21856
rect 12525 21798 14780 21800
rect 12525 21795 12591 21798
rect 14774 21796 14780 21798
rect 14844 21796 14850 21860
rect 15929 21858 15995 21861
rect 23473 21858 23539 21861
rect 15929 21856 23539 21858
rect 15929 21800 15934 21856
rect 15990 21800 23478 21856
rect 23534 21800 23539 21856
rect 15929 21798 23539 21800
rect 15929 21795 15995 21798
rect 23473 21795 23539 21798
rect 24761 21858 24827 21861
rect 27520 21858 28000 21888
rect 24761 21856 28000 21858
rect 24761 21800 24766 21856
rect 24822 21800 28000 21856
rect 24761 21798 28000 21800
rect 24761 21795 24827 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21798
rect 24277 21727 24597 21728
rect 6361 21450 6427 21453
rect 11053 21450 11119 21453
rect 6361 21448 11119 21450
rect 6361 21392 6366 21448
rect 6422 21392 11058 21448
rect 11114 21392 11119 21448
rect 6361 21390 11119 21392
rect 6361 21387 6427 21390
rect 11053 21387 11119 21390
rect 15285 21450 15351 21453
rect 19149 21450 19215 21453
rect 15285 21448 19215 21450
rect 15285 21392 15290 21448
rect 15346 21392 19154 21448
rect 19210 21392 19215 21448
rect 15285 21390 19215 21392
rect 15285 21387 15351 21390
rect 19149 21387 19215 21390
rect 23657 21314 23723 21317
rect 27520 21314 28000 21344
rect 23657 21312 28000 21314
rect 23657 21256 23662 21312
rect 23718 21256 28000 21312
rect 23657 21254 28000 21256
rect 23657 21251 23723 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 12801 21178 12867 21181
rect 17677 21178 17743 21181
rect 12801 21176 17743 21178
rect 12801 21120 12806 21176
rect 12862 21120 17682 21176
rect 17738 21120 17743 21176
rect 12801 21118 17743 21120
rect 12801 21115 12867 21118
rect 17677 21115 17743 21118
rect 15469 21042 15535 21045
rect 23749 21042 23815 21045
rect 15469 21040 23815 21042
rect 15469 20984 15474 21040
rect 15530 20984 23754 21040
rect 23810 20984 23815 21040
rect 15469 20982 23815 20984
rect 15469 20979 15535 20982
rect 23749 20979 23815 20982
rect 1577 20906 1643 20909
rect 21357 20906 21423 20909
rect 1577 20904 21423 20906
rect 1577 20848 1582 20904
rect 1638 20848 21362 20904
rect 21418 20848 21423 20904
rect 1577 20846 21423 20848
rect 1577 20843 1643 20846
rect 21357 20843 21423 20846
rect 9121 20770 9187 20773
rect 13813 20770 13879 20773
rect 9121 20768 13879 20770
rect 9121 20712 9126 20768
rect 9182 20712 13818 20768
rect 13874 20712 13879 20768
rect 9121 20710 13879 20712
rect 9121 20707 9187 20710
rect 13813 20707 13879 20710
rect 24945 20770 25011 20773
rect 27520 20770 28000 20800
rect 24945 20768 28000 20770
rect 24945 20712 24950 20768
rect 25006 20712 28000 20768
rect 24945 20710 28000 20712
rect 24945 20707 25011 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 15377 20634 15443 20637
rect 21081 20634 21147 20637
rect 15377 20632 21147 20634
rect 15377 20576 15382 20632
rect 15438 20576 21086 20632
rect 21142 20576 21147 20632
rect 15377 20574 21147 20576
rect 15377 20571 15443 20574
rect 21081 20571 21147 20574
rect 10777 20498 10843 20501
rect 12893 20498 12959 20501
rect 10777 20496 12959 20498
rect 10777 20440 10782 20496
rect 10838 20440 12898 20496
rect 12954 20440 12959 20496
rect 10777 20438 12959 20440
rect 10777 20435 10843 20438
rect 12893 20435 12959 20438
rect 13261 20498 13327 20501
rect 15837 20498 15903 20501
rect 16297 20498 16363 20501
rect 13261 20496 16363 20498
rect 13261 20440 13266 20496
rect 13322 20440 15842 20496
rect 15898 20440 16302 20496
rect 16358 20440 16363 20496
rect 13261 20438 16363 20440
rect 13261 20435 13327 20438
rect 15837 20435 15903 20438
rect 16297 20435 16363 20438
rect 1577 20362 1643 20365
rect 24761 20362 24827 20365
rect 1577 20360 24827 20362
rect 1577 20304 1582 20360
rect 1638 20304 24766 20360
rect 24822 20304 24827 20360
rect 1577 20302 24827 20304
rect 1577 20299 1643 20302
rect 24761 20299 24827 20302
rect 10961 20226 11027 20229
rect 15653 20226 15719 20229
rect 16665 20226 16731 20229
rect 10961 20224 16731 20226
rect 10961 20168 10966 20224
rect 11022 20168 15658 20224
rect 15714 20168 16670 20224
rect 16726 20168 16731 20224
rect 10961 20166 16731 20168
rect 10961 20163 11027 20166
rect 15653 20163 15719 20166
rect 16665 20163 16731 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 12433 20090 12499 20093
rect 14365 20090 14431 20093
rect 27520 20090 28000 20120
rect 12433 20088 14431 20090
rect 12433 20032 12438 20088
rect 12494 20032 14370 20088
rect 14426 20032 14431 20088
rect 12433 20030 14431 20032
rect 12433 20027 12499 20030
rect 14365 20027 14431 20030
rect 23982 20030 28000 20090
rect 7741 19954 7807 19957
rect 12341 19954 12407 19957
rect 7741 19952 12407 19954
rect 7741 19896 7746 19952
rect 7802 19896 12346 19952
rect 12402 19896 12407 19952
rect 7741 19894 12407 19896
rect 7741 19891 7807 19894
rect 12341 19891 12407 19894
rect 14089 19954 14155 19957
rect 20897 19954 20963 19957
rect 23657 19954 23723 19957
rect 14089 19952 20546 19954
rect 14089 19896 14094 19952
rect 14150 19896 20546 19952
rect 14089 19894 20546 19896
rect 14089 19891 14155 19894
rect 14089 19818 14155 19821
rect 20345 19818 20411 19821
rect 14089 19816 20411 19818
rect 14089 19760 14094 19816
rect 14150 19760 20350 19816
rect 20406 19760 20411 19816
rect 14089 19758 20411 19760
rect 20486 19818 20546 19894
rect 20897 19952 23723 19954
rect 20897 19896 20902 19952
rect 20958 19896 23662 19952
rect 23718 19896 23723 19952
rect 20897 19894 23723 19896
rect 20897 19891 20963 19894
rect 23657 19891 23723 19894
rect 21357 19818 21423 19821
rect 20486 19816 21423 19818
rect 20486 19760 21362 19816
rect 21418 19760 21423 19816
rect 20486 19758 21423 19760
rect 14089 19755 14155 19758
rect 20345 19755 20411 19758
rect 21357 19755 21423 19758
rect 15561 19682 15627 19685
rect 23982 19682 24042 20030
rect 27520 20000 28000 20030
rect 15561 19680 24042 19682
rect 15561 19624 15566 19680
rect 15622 19624 24042 19680
rect 15561 19622 24042 19624
rect 15561 19619 15627 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19546 28000 19576
rect 24718 19486 28000 19546
rect 11145 19410 11211 19413
rect 12801 19410 12867 19413
rect 14825 19412 14891 19413
rect 11145 19408 12867 19410
rect 11145 19352 11150 19408
rect 11206 19352 12806 19408
rect 12862 19352 12867 19408
rect 11145 19350 12867 19352
rect 11145 19347 11211 19350
rect 12801 19347 12867 19350
rect 14774 19348 14780 19412
rect 14844 19410 14891 19412
rect 18689 19410 18755 19413
rect 20437 19410 20503 19413
rect 14844 19408 14936 19410
rect 14886 19352 14936 19408
rect 14844 19350 14936 19352
rect 18689 19408 20503 19410
rect 18689 19352 18694 19408
rect 18750 19352 20442 19408
rect 20498 19352 20503 19408
rect 18689 19350 20503 19352
rect 14844 19348 14891 19350
rect 14825 19347 14891 19348
rect 18689 19347 18755 19350
rect 20437 19347 20503 19350
rect 22645 19410 22711 19413
rect 24718 19410 24778 19486
rect 27520 19456 28000 19486
rect 22645 19408 24778 19410
rect 22645 19352 22650 19408
rect 22706 19352 24778 19408
rect 22645 19350 24778 19352
rect 22645 19347 22711 19350
rect 7097 19274 7163 19277
rect 10869 19274 10935 19277
rect 7097 19272 10935 19274
rect 7097 19216 7102 19272
rect 7158 19216 10874 19272
rect 10930 19216 10935 19272
rect 7097 19214 10935 19216
rect 7097 19211 7163 19214
rect 10869 19211 10935 19214
rect 17217 19274 17283 19277
rect 21541 19274 21607 19277
rect 17217 19272 21607 19274
rect 17217 19216 17222 19272
rect 17278 19216 21546 19272
rect 21602 19216 21607 19272
rect 17217 19214 21607 19216
rect 17217 19211 17283 19214
rect 21541 19211 21607 19214
rect 12893 19138 12959 19141
rect 13353 19138 13419 19141
rect 18321 19138 18387 19141
rect 12893 19136 18387 19138
rect 12893 19080 12898 19136
rect 12954 19080 13358 19136
rect 13414 19080 18326 19136
rect 18382 19080 18387 19136
rect 12893 19078 18387 19080
rect 12893 19075 12959 19078
rect 13353 19075 13419 19078
rect 18321 19075 18387 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 17677 19002 17743 19005
rect 17861 19002 17927 19005
rect 19425 19002 19491 19005
rect 17677 19000 19491 19002
rect 17677 18944 17682 19000
rect 17738 18944 17866 19000
rect 17922 18944 19430 19000
rect 19486 18944 19491 19000
rect 17677 18942 19491 18944
rect 17677 18939 17743 18942
rect 17861 18939 17927 18942
rect 19425 18939 19491 18942
rect 24761 19002 24827 19005
rect 27520 19002 28000 19032
rect 24761 19000 28000 19002
rect 24761 18944 24766 19000
rect 24822 18944 28000 19000
rect 24761 18942 28000 18944
rect 24761 18939 24827 18942
rect 27520 18912 28000 18942
rect 19793 18866 19859 18869
rect 20345 18866 20411 18869
rect 23933 18866 23999 18869
rect 19793 18864 23999 18866
rect 19793 18808 19798 18864
rect 19854 18808 20350 18864
rect 20406 18808 23938 18864
rect 23994 18808 23999 18864
rect 19793 18806 23999 18808
rect 19793 18803 19859 18806
rect 20345 18803 20411 18806
rect 23933 18803 23999 18806
rect 14825 18730 14891 18733
rect 19374 18730 19380 18732
rect 14825 18728 19380 18730
rect 14825 18672 14830 18728
rect 14886 18672 19380 18728
rect 14825 18670 19380 18672
rect 14825 18667 14891 18670
rect 19374 18668 19380 18670
rect 19444 18730 19450 18732
rect 23197 18730 23263 18733
rect 19444 18728 23263 18730
rect 19444 18672 23202 18728
rect 23258 18672 23263 18728
rect 19444 18670 23263 18672
rect 19444 18668 19450 18670
rect 23197 18667 23263 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 25681 18458 25747 18461
rect 27520 18458 28000 18488
rect 25681 18456 28000 18458
rect 25681 18400 25686 18456
rect 25742 18400 28000 18456
rect 25681 18398 28000 18400
rect 25681 18395 25747 18398
rect 27520 18368 28000 18398
rect 19977 18322 20043 18325
rect 25221 18322 25287 18325
rect 19977 18320 25287 18322
rect 19977 18264 19982 18320
rect 20038 18264 25226 18320
rect 25282 18264 25287 18320
rect 19977 18262 25287 18264
rect 19977 18259 20043 18262
rect 25221 18259 25287 18262
rect 13261 18186 13327 18189
rect 19241 18186 19307 18189
rect 21173 18186 21239 18189
rect 13261 18184 15946 18186
rect 13261 18128 13266 18184
rect 13322 18128 15946 18184
rect 13261 18126 15946 18128
rect 13261 18123 13327 18126
rect 12801 18050 12867 18053
rect 15745 18050 15811 18053
rect 12801 18048 15811 18050
rect 12801 17992 12806 18048
rect 12862 17992 15750 18048
rect 15806 17992 15811 18048
rect 12801 17990 15811 17992
rect 12801 17987 12867 17990
rect 15745 17987 15811 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 15886 17778 15946 18126
rect 19241 18184 21239 18186
rect 19241 18128 19246 18184
rect 19302 18128 21178 18184
rect 21234 18128 21239 18184
rect 19241 18126 21239 18128
rect 19241 18123 19307 18126
rect 21173 18123 21239 18126
rect 21909 18186 21975 18189
rect 24853 18186 24919 18189
rect 21909 18184 24919 18186
rect 21909 18128 21914 18184
rect 21970 18128 24858 18184
rect 24914 18128 24919 18184
rect 21909 18126 24919 18128
rect 21909 18123 21975 18126
rect 24853 18123 24919 18126
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 20069 17914 20135 17917
rect 25497 17914 25563 17917
rect 20069 17912 25563 17914
rect 20069 17856 20074 17912
rect 20130 17856 25502 17912
rect 25558 17856 25563 17912
rect 20069 17854 25563 17856
rect 20069 17851 20135 17854
rect 25497 17851 25563 17854
rect 20253 17778 20319 17781
rect 15886 17776 20319 17778
rect 15886 17720 20258 17776
rect 20314 17720 20319 17776
rect 15886 17718 20319 17720
rect 20253 17715 20319 17718
rect 20989 17778 21055 17781
rect 24025 17778 24091 17781
rect 20989 17776 24091 17778
rect 20989 17720 20994 17776
rect 21050 17720 24030 17776
rect 24086 17720 24091 17776
rect 20989 17718 24091 17720
rect 20989 17715 21055 17718
rect 24025 17715 24091 17718
rect 25405 17778 25471 17781
rect 27520 17778 28000 17808
rect 25405 17776 28000 17778
rect 25405 17720 25410 17776
rect 25466 17720 28000 17776
rect 25405 17718 28000 17720
rect 25405 17715 25471 17718
rect 27520 17688 28000 17718
rect 10869 17642 10935 17645
rect 11145 17642 11211 17645
rect 18045 17642 18111 17645
rect 10869 17640 18111 17642
rect 10869 17584 10874 17640
rect 10930 17584 11150 17640
rect 11206 17584 18050 17640
rect 18106 17584 18111 17640
rect 10869 17582 18111 17584
rect 10869 17579 10935 17582
rect 11145 17579 11211 17582
rect 18045 17579 18111 17582
rect 19793 17642 19859 17645
rect 20345 17642 20411 17645
rect 23197 17642 23263 17645
rect 19793 17640 23263 17642
rect 19793 17584 19798 17640
rect 19854 17584 20350 17640
rect 20406 17584 23202 17640
rect 23258 17584 23263 17640
rect 19793 17582 23263 17584
rect 19793 17579 19859 17582
rect 20345 17579 20411 17582
rect 23197 17579 23263 17582
rect 15653 17506 15719 17509
rect 20437 17506 20503 17509
rect 15653 17504 20503 17506
rect 15653 17448 15658 17504
rect 15714 17448 20442 17504
rect 20498 17448 20503 17504
rect 15653 17446 20503 17448
rect 15653 17443 15719 17446
rect 20437 17443 20503 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 17401 17370 17467 17373
rect 23197 17370 23263 17373
rect 17401 17368 23263 17370
rect 17401 17312 17406 17368
rect 17462 17312 23202 17368
rect 23258 17312 23263 17368
rect 17401 17310 23263 17312
rect 17401 17307 17467 17310
rect 23197 17307 23263 17310
rect 14273 17234 14339 17237
rect 20713 17234 20779 17237
rect 14273 17232 20779 17234
rect 14273 17176 14278 17232
rect 14334 17176 20718 17232
rect 20774 17176 20779 17232
rect 14273 17174 20779 17176
rect 14273 17171 14339 17174
rect 20713 17171 20779 17174
rect 24945 17234 25011 17237
rect 27520 17234 28000 17264
rect 24945 17232 28000 17234
rect 24945 17176 24950 17232
rect 25006 17176 28000 17232
rect 24945 17174 28000 17176
rect 24945 17171 25011 17174
rect 27520 17144 28000 17174
rect 11421 17098 11487 17101
rect 19333 17098 19399 17101
rect 11421 17096 19399 17098
rect 11421 17040 11426 17096
rect 11482 17040 19338 17096
rect 19394 17040 19399 17096
rect 11421 17038 19399 17040
rect 11421 17035 11487 17038
rect 19333 17035 19399 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 14365 16690 14431 16693
rect 24025 16690 24091 16693
rect 14365 16688 24091 16690
rect 14365 16632 14370 16688
rect 14426 16632 24030 16688
rect 24086 16632 24091 16688
rect 14365 16630 24091 16632
rect 14365 16627 14431 16630
rect 24025 16627 24091 16630
rect 25129 16690 25195 16693
rect 27520 16690 28000 16720
rect 25129 16688 28000 16690
rect 25129 16632 25134 16688
rect 25190 16632 28000 16688
rect 25129 16630 28000 16632
rect 25129 16627 25195 16630
rect 27520 16600 28000 16630
rect 12985 16554 13051 16557
rect 16021 16554 16087 16557
rect 2638 16494 7666 16554
rect 381 16282 447 16285
rect 2638 16282 2698 16494
rect 7606 16418 7666 16494
rect 12985 16552 16087 16554
rect 12985 16496 12990 16552
rect 13046 16496 16026 16552
rect 16082 16496 16087 16552
rect 12985 16494 16087 16496
rect 12985 16491 13051 16494
rect 16021 16491 16087 16494
rect 13445 16418 13511 16421
rect 21265 16418 21331 16421
rect 23197 16418 23263 16421
rect 7606 16416 13511 16418
rect 7606 16360 13450 16416
rect 13506 16360 13511 16416
rect 7606 16358 13511 16360
rect 13445 16355 13511 16358
rect 15334 16416 23263 16418
rect 15334 16360 21270 16416
rect 21326 16360 23202 16416
rect 23258 16360 23263 16416
rect 15334 16358 23263 16360
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 381 16280 2698 16282
rect 381 16224 386 16280
rect 442 16224 2698 16280
rect 381 16222 2698 16224
rect 381 16219 447 16222
rect 15101 16146 15167 16149
rect 15334 16146 15394 16358
rect 21265 16355 21331 16358
rect 23197 16355 23263 16358
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 17769 16282 17835 16285
rect 24117 16282 24183 16285
rect 17769 16280 24183 16282
rect 17769 16224 17774 16280
rect 17830 16224 24122 16280
rect 24178 16224 24183 16280
rect 17769 16222 24183 16224
rect 17769 16219 17835 16222
rect 24117 16219 24183 16222
rect 15101 16144 15394 16146
rect 15101 16088 15106 16144
rect 15162 16088 15394 16144
rect 15101 16086 15394 16088
rect 15101 16083 15167 16086
rect 19057 16010 19123 16013
rect 21449 16010 21515 16013
rect 19057 16008 21515 16010
rect 19057 15952 19062 16008
rect 19118 15952 21454 16008
rect 21510 15952 21515 16008
rect 19057 15950 21515 15952
rect 19057 15947 19123 15950
rect 21449 15947 21515 15950
rect 24761 16010 24827 16013
rect 27520 16010 28000 16040
rect 24761 16008 28000 16010
rect 24761 15952 24766 16008
rect 24822 15952 28000 16008
rect 24761 15950 28000 15952
rect 24761 15947 24827 15950
rect 27520 15920 28000 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 16205 15602 16271 15605
rect 18229 15602 18295 15605
rect 16205 15600 18295 15602
rect 16205 15544 16210 15600
rect 16266 15544 18234 15600
rect 18290 15544 18295 15600
rect 16205 15542 18295 15544
rect 16205 15539 16271 15542
rect 18229 15539 18295 15542
rect 24761 15466 24827 15469
rect 27520 15466 28000 15496
rect 24761 15464 28000 15466
rect 24761 15408 24766 15464
rect 24822 15408 28000 15464
rect 24761 15406 28000 15408
rect 24761 15403 24827 15406
rect 27520 15376 28000 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 15653 15194 15719 15197
rect 23933 15194 23999 15197
rect 15653 15192 23999 15194
rect 15653 15136 15658 15192
rect 15714 15136 23938 15192
rect 23994 15136 23999 15192
rect 15653 15134 23999 15136
rect 15653 15131 15719 15134
rect 23933 15131 23999 15134
rect 13721 15058 13787 15061
rect 24577 15058 24643 15061
rect 13721 15056 24643 15058
rect 13721 15000 13726 15056
rect 13782 15000 24582 15056
rect 24638 15000 24643 15056
rect 13721 14998 24643 15000
rect 13721 14995 13787 14998
rect 24577 14995 24643 14998
rect 17217 14922 17283 14925
rect 24393 14922 24459 14925
rect 17217 14920 24459 14922
rect 17217 14864 17222 14920
rect 17278 14864 24398 14920
rect 24454 14864 24459 14920
rect 17217 14862 24459 14864
rect 17217 14859 17283 14862
rect 24393 14859 24459 14862
rect 24761 14922 24827 14925
rect 27520 14922 28000 14952
rect 24761 14920 28000 14922
rect 24761 14864 24766 14920
rect 24822 14864 28000 14920
rect 24761 14862 28000 14864
rect 24761 14859 24827 14862
rect 27520 14832 28000 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 14181 14514 14247 14517
rect 17953 14514 18019 14517
rect 14181 14512 18019 14514
rect 14181 14456 14186 14512
rect 14242 14456 17958 14512
rect 18014 14456 18019 14512
rect 14181 14454 18019 14456
rect 14181 14451 14247 14454
rect 17953 14451 18019 14454
rect 18597 14514 18663 14517
rect 21909 14514 21975 14517
rect 18597 14512 21975 14514
rect 18597 14456 18602 14512
rect 18658 14456 21914 14512
rect 21970 14456 21975 14512
rect 18597 14454 21975 14456
rect 18597 14451 18663 14454
rect 21909 14451 21975 14454
rect 8201 14378 8267 14381
rect 13629 14378 13695 14381
rect 8201 14376 13695 14378
rect 8201 14320 8206 14376
rect 8262 14320 13634 14376
rect 13690 14320 13695 14376
rect 8201 14318 13695 14320
rect 8201 14315 8267 14318
rect 13629 14315 13695 14318
rect 14273 14378 14339 14381
rect 27520 14378 28000 14408
rect 14273 14376 28000 14378
rect 14273 14320 14278 14376
rect 14334 14320 28000 14376
rect 14273 14318 28000 14320
rect 14273 14315 14339 14318
rect 27520 14288 28000 14318
rect 17401 14242 17467 14245
rect 19241 14242 19307 14245
rect 17401 14240 19307 14242
rect 17401 14184 17406 14240
rect 17462 14184 19246 14240
rect 19302 14184 19307 14240
rect 17401 14182 19307 14184
rect 17401 14179 17467 14182
rect 19241 14179 19307 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10961 14106 11027 14109
rect 14273 14106 14339 14109
rect 10961 14104 14339 14106
rect 10961 14048 10966 14104
rect 11022 14048 14278 14104
rect 14334 14048 14339 14104
rect 10961 14046 14339 14048
rect 10961 14043 11027 14046
rect 14273 14043 14339 14046
rect 0 13970 480 14000
rect 1669 13970 1735 13973
rect 0 13968 1735 13970
rect 0 13912 1674 13968
rect 1730 13912 1735 13968
rect 0 13910 1735 13912
rect 0 13880 480 13910
rect 1669 13907 1735 13910
rect 14825 13970 14891 13973
rect 20897 13970 20963 13973
rect 14825 13968 20963 13970
rect 14825 13912 14830 13968
rect 14886 13912 20902 13968
rect 20958 13912 20963 13968
rect 14825 13910 20963 13912
rect 14825 13907 14891 13910
rect 20897 13907 20963 13910
rect 12065 13834 12131 13837
rect 12985 13834 13051 13837
rect 12065 13832 13051 13834
rect 12065 13776 12070 13832
rect 12126 13776 12990 13832
rect 13046 13776 13051 13832
rect 12065 13774 13051 13776
rect 12065 13771 12131 13774
rect 12985 13771 13051 13774
rect 13261 13834 13327 13837
rect 16481 13834 16547 13837
rect 13261 13832 16547 13834
rect 13261 13776 13266 13832
rect 13322 13776 16486 13832
rect 16542 13776 16547 13832
rect 13261 13774 16547 13776
rect 13261 13771 13327 13774
rect 16481 13771 16547 13774
rect 21081 13834 21147 13837
rect 24669 13834 24735 13837
rect 21081 13832 24735 13834
rect 21081 13776 21086 13832
rect 21142 13776 24674 13832
rect 24730 13776 24735 13832
rect 21081 13774 24735 13776
rect 21081 13771 21147 13774
rect 24669 13771 24735 13774
rect 11053 13698 11119 13701
rect 17769 13698 17835 13701
rect 11053 13696 17835 13698
rect 11053 13640 11058 13696
rect 11114 13640 17774 13696
rect 17830 13640 17835 13696
rect 11053 13638 17835 13640
rect 11053 13635 11119 13638
rect 17769 13635 17835 13638
rect 24761 13698 24827 13701
rect 27520 13698 28000 13728
rect 24761 13696 28000 13698
rect 24761 13640 24766 13696
rect 24822 13640 28000 13696
rect 24761 13638 28000 13640
rect 24761 13635 24827 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 13997 13562 14063 13565
rect 19425 13562 19491 13565
rect 13997 13560 19491 13562
rect 13997 13504 14002 13560
rect 14058 13504 19430 13560
rect 19486 13504 19491 13560
rect 13997 13502 19491 13504
rect 13997 13499 14063 13502
rect 19425 13499 19491 13502
rect 12709 13426 12775 13429
rect 5398 13424 12775 13426
rect 5398 13368 12714 13424
rect 12770 13368 12775 13424
rect 5398 13366 12775 13368
rect 2313 13154 2379 13157
rect 5398 13154 5458 13366
rect 12709 13363 12775 13366
rect 16481 13426 16547 13429
rect 24577 13426 24643 13429
rect 16481 13424 24643 13426
rect 16481 13368 16486 13424
rect 16542 13368 24582 13424
rect 24638 13368 24643 13424
rect 16481 13366 24643 13368
rect 16481 13363 16547 13366
rect 24577 13363 24643 13366
rect 8385 13290 8451 13293
rect 15561 13290 15627 13293
rect 8385 13288 15627 13290
rect 8385 13232 8390 13288
rect 8446 13232 15566 13288
rect 15622 13232 15627 13288
rect 8385 13230 15627 13232
rect 8385 13227 8451 13230
rect 15561 13227 15627 13230
rect 2313 13152 5458 13154
rect 2313 13096 2318 13152
rect 2374 13096 5458 13152
rect 2313 13094 5458 13096
rect 16297 13154 16363 13157
rect 22553 13154 22619 13157
rect 16297 13152 22619 13154
rect 16297 13096 16302 13152
rect 16358 13096 22558 13152
rect 22614 13096 22619 13152
rect 16297 13094 22619 13096
rect 2313 13091 2379 13094
rect 16297 13091 16363 13094
rect 22553 13091 22619 13094
rect 24761 13154 24827 13157
rect 27520 13154 28000 13184
rect 24761 13152 28000 13154
rect 24761 13096 24766 13152
rect 24822 13096 28000 13152
rect 24761 13094 28000 13096
rect 24761 13091 24827 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 20161 13018 20227 13021
rect 22277 13018 22343 13021
rect 20161 13016 22343 13018
rect 20161 12960 20166 13016
rect 20222 12960 22282 13016
rect 22338 12960 22343 13016
rect 20161 12958 22343 12960
rect 20161 12955 20227 12958
rect 22277 12955 22343 12958
rect 13813 12882 13879 12885
rect 24577 12882 24643 12885
rect 13813 12880 24643 12882
rect 13813 12824 13818 12880
rect 13874 12824 24582 12880
rect 24638 12824 24643 12880
rect 13813 12822 24643 12824
rect 13813 12819 13879 12822
rect 24577 12819 24643 12822
rect 12709 12746 12775 12749
rect 18781 12746 18847 12749
rect 12709 12744 18847 12746
rect 12709 12688 12714 12744
rect 12770 12688 18786 12744
rect 18842 12688 18847 12744
rect 12709 12686 18847 12688
rect 12709 12683 12775 12686
rect 18781 12683 18847 12686
rect 19057 12746 19123 12749
rect 22093 12746 22159 12749
rect 19057 12744 22159 12746
rect 19057 12688 19062 12744
rect 19118 12688 22098 12744
rect 22154 12688 22159 12744
rect 19057 12686 22159 12688
rect 19057 12683 19123 12686
rect 22093 12683 22159 12686
rect 12341 12610 12407 12613
rect 16389 12610 16455 12613
rect 12341 12608 16455 12610
rect 12341 12552 12346 12608
rect 12402 12552 16394 12608
rect 16450 12552 16455 12608
rect 12341 12550 16455 12552
rect 12341 12547 12407 12550
rect 16389 12547 16455 12550
rect 24761 12610 24827 12613
rect 27520 12610 28000 12640
rect 24761 12608 28000 12610
rect 24761 12552 24766 12608
rect 24822 12552 28000 12608
rect 24761 12550 28000 12552
rect 24761 12547 24827 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 11881 12474 11947 12477
rect 16297 12474 16363 12477
rect 11881 12472 16363 12474
rect 11881 12416 11886 12472
rect 11942 12416 16302 12472
rect 16358 12416 16363 12472
rect 11881 12414 16363 12416
rect 11881 12411 11947 12414
rect 16297 12411 16363 12414
rect 17125 12474 17191 12477
rect 17493 12474 17559 12477
rect 17125 12472 17559 12474
rect 17125 12416 17130 12472
rect 17186 12416 17498 12472
rect 17554 12416 17559 12472
rect 17125 12414 17559 12416
rect 17125 12411 17191 12414
rect 17493 12411 17559 12414
rect 22185 12338 22251 12341
rect 24577 12338 24643 12341
rect 22185 12336 24643 12338
rect 22185 12280 22190 12336
rect 22246 12280 24582 12336
rect 24638 12280 24643 12336
rect 22185 12278 24643 12280
rect 22185 12275 22251 12278
rect 24577 12275 24643 12278
rect 20069 12066 20135 12069
rect 22461 12066 22527 12069
rect 20069 12064 22527 12066
rect 20069 12008 20074 12064
rect 20130 12008 22466 12064
rect 22522 12008 22527 12064
rect 20069 12006 22527 12008
rect 20069 12003 20135 12006
rect 22461 12003 22527 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 18965 11930 19031 11933
rect 22737 11930 22803 11933
rect 18965 11928 22803 11930
rect 18965 11872 18970 11928
rect 19026 11872 22742 11928
rect 22798 11872 22803 11928
rect 18965 11870 22803 11872
rect 18965 11867 19031 11870
rect 22737 11867 22803 11870
rect 24761 11930 24827 11933
rect 27520 11930 28000 11960
rect 24761 11928 28000 11930
rect 24761 11872 24766 11928
rect 24822 11872 28000 11928
rect 24761 11870 28000 11872
rect 24761 11867 24827 11870
rect 27520 11840 28000 11870
rect 17217 11794 17283 11797
rect 23657 11794 23723 11797
rect 17217 11792 23723 11794
rect 17217 11736 17222 11792
rect 17278 11736 23662 11792
rect 23718 11736 23723 11792
rect 17217 11734 23723 11736
rect 17217 11731 17283 11734
rect 23657 11731 23723 11734
rect 13261 11658 13327 11661
rect 20437 11658 20503 11661
rect 13261 11656 20503 11658
rect 13261 11600 13266 11656
rect 13322 11600 20442 11656
rect 20498 11600 20503 11656
rect 13261 11598 20503 11600
rect 13261 11595 13327 11598
rect 20437 11595 20503 11598
rect 13905 11522 13971 11525
rect 15377 11522 15443 11525
rect 13905 11520 15443 11522
rect 13905 11464 13910 11520
rect 13966 11464 15382 11520
rect 15438 11464 15443 11520
rect 13905 11462 15443 11464
rect 13905 11459 13971 11462
rect 15377 11459 15443 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 24669 11386 24735 11389
rect 27520 11386 28000 11416
rect 24669 11384 28000 11386
rect 24669 11328 24674 11384
rect 24730 11328 28000 11384
rect 24669 11326 28000 11328
rect 24669 11323 24735 11326
rect 27520 11296 28000 11326
rect 19241 11250 19307 11253
rect 20621 11250 20687 11253
rect 19241 11248 20687 11250
rect 19241 11192 19246 11248
rect 19302 11192 20626 11248
rect 20682 11192 20687 11248
rect 19241 11190 20687 11192
rect 19241 11187 19307 11190
rect 20621 11187 20687 11190
rect 4981 11114 5047 11117
rect 12341 11114 12407 11117
rect 4981 11112 12407 11114
rect 4981 11056 4986 11112
rect 5042 11056 12346 11112
rect 12402 11056 12407 11112
rect 4981 11054 12407 11056
rect 4981 11051 5047 11054
rect 12341 11051 12407 11054
rect 19374 11052 19380 11116
rect 19444 11114 19450 11116
rect 19517 11114 19583 11117
rect 19444 11112 19583 11114
rect 19444 11056 19522 11112
rect 19578 11056 19583 11112
rect 19444 11054 19583 11056
rect 19444 11052 19450 11054
rect 19517 11051 19583 11054
rect 21541 11114 21607 11117
rect 24761 11114 24827 11117
rect 21541 11112 24827 11114
rect 21541 11056 21546 11112
rect 21602 11056 24766 11112
rect 24822 11056 24827 11112
rect 21541 11054 24827 11056
rect 21541 11051 21607 11054
rect 24761 11051 24827 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 24761 10842 24827 10845
rect 27520 10842 28000 10872
rect 24761 10840 28000 10842
rect 24761 10784 24766 10840
rect 24822 10784 28000 10840
rect 24761 10782 28000 10784
rect 24761 10779 24827 10782
rect 27520 10752 28000 10782
rect 14457 10706 14523 10709
rect 16665 10706 16731 10709
rect 14457 10704 16731 10706
rect 14457 10648 14462 10704
rect 14518 10648 16670 10704
rect 16726 10648 16731 10704
rect 14457 10646 16731 10648
rect 14457 10643 14523 10646
rect 16665 10643 16731 10646
rect 17033 10706 17099 10709
rect 23197 10706 23263 10709
rect 17033 10704 23263 10706
rect 17033 10648 17038 10704
rect 17094 10648 23202 10704
rect 23258 10648 23263 10704
rect 17033 10646 23263 10648
rect 17033 10643 17099 10646
rect 23197 10643 23263 10646
rect 1485 10570 1551 10573
rect 2865 10570 2931 10573
rect 1485 10568 2931 10570
rect 1485 10512 1490 10568
rect 1546 10512 2870 10568
rect 2926 10512 2931 10568
rect 1485 10510 2931 10512
rect 1485 10507 1551 10510
rect 2865 10507 2931 10510
rect 4337 10570 4403 10573
rect 13537 10570 13603 10573
rect 21265 10570 21331 10573
rect 4337 10568 13603 10570
rect 4337 10512 4342 10568
rect 4398 10512 13542 10568
rect 13598 10512 13603 10568
rect 4337 10510 13603 10512
rect 4337 10507 4403 10510
rect 13537 10507 13603 10510
rect 19382 10568 21331 10570
rect 19382 10512 21270 10568
rect 21326 10512 21331 10568
rect 19382 10510 21331 10512
rect 13353 10434 13419 10437
rect 19382 10434 19442 10510
rect 21265 10507 21331 10510
rect 13353 10432 19442 10434
rect 13353 10376 13358 10432
rect 13414 10376 19442 10432
rect 13353 10374 19442 10376
rect 13353 10371 13419 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 14181 10298 14247 10301
rect 18413 10298 18479 10301
rect 19425 10298 19491 10301
rect 14181 10296 19491 10298
rect 14181 10240 14186 10296
rect 14242 10240 18418 10296
rect 18474 10240 19430 10296
rect 19486 10240 19491 10296
rect 14181 10238 19491 10240
rect 14181 10235 14247 10238
rect 18413 10235 18479 10238
rect 19425 10235 19491 10238
rect 21357 10298 21423 10301
rect 24669 10298 24735 10301
rect 21357 10296 24735 10298
rect 21357 10240 21362 10296
rect 21418 10240 24674 10296
rect 24730 10240 24735 10296
rect 21357 10238 24735 10240
rect 21357 10235 21423 10238
rect 24669 10235 24735 10238
rect 27520 10162 28000 10192
rect 23476 10102 28000 10162
rect 14089 10026 14155 10029
rect 21357 10026 21423 10029
rect 14089 10024 21423 10026
rect 14089 9968 14094 10024
rect 14150 9968 21362 10024
rect 21418 9968 21423 10024
rect 14089 9966 21423 9968
rect 14089 9963 14155 9966
rect 21357 9963 21423 9966
rect 15653 9890 15719 9893
rect 16757 9890 16823 9893
rect 23476 9890 23536 10102
rect 27520 10072 28000 10102
rect 15653 9888 23536 9890
rect 15653 9832 15658 9888
rect 15714 9832 16762 9888
rect 16818 9832 23536 9888
rect 15653 9830 23536 9832
rect 15653 9827 15719 9830
rect 16757 9827 16823 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 2773 9618 2839 9621
rect 9949 9618 10015 9621
rect 2773 9616 10015 9618
rect 2773 9560 2778 9616
rect 2834 9560 9954 9616
rect 10010 9560 10015 9616
rect 2773 9558 10015 9560
rect 2773 9555 2839 9558
rect 9949 9555 10015 9558
rect 18505 9618 18571 9621
rect 27520 9618 28000 9648
rect 18505 9616 28000 9618
rect 18505 9560 18510 9616
rect 18566 9560 28000 9616
rect 18505 9558 28000 9560
rect 18505 9555 18571 9558
rect 27520 9528 28000 9558
rect 17861 9482 17927 9485
rect 18781 9482 18847 9485
rect 24669 9482 24735 9485
rect 17861 9480 24735 9482
rect 17861 9424 17866 9480
rect 17922 9424 18786 9480
rect 18842 9424 24674 9480
rect 24730 9424 24735 9480
rect 17861 9422 24735 9424
rect 17861 9419 17927 9422
rect 18781 9419 18847 9422
rect 24669 9419 24735 9422
rect 2865 9346 2931 9349
rect 9673 9346 9739 9349
rect 2865 9344 9739 9346
rect 2865 9288 2870 9344
rect 2926 9288 9678 9344
rect 9734 9288 9739 9344
rect 2865 9286 9739 9288
rect 2865 9283 2931 9286
rect 9673 9283 9739 9286
rect 12433 9346 12499 9349
rect 13353 9346 13419 9349
rect 12433 9344 13419 9346
rect 12433 9288 12438 9344
rect 12494 9288 13358 9344
rect 13414 9288 13419 9344
rect 12433 9286 13419 9288
rect 12433 9283 12499 9286
rect 13353 9283 13419 9286
rect 15009 9346 15075 9349
rect 16665 9346 16731 9349
rect 15009 9344 16731 9346
rect 15009 9288 15014 9344
rect 15070 9288 16670 9344
rect 16726 9288 16731 9344
rect 15009 9286 16731 9288
rect 15009 9283 15075 9286
rect 16665 9283 16731 9286
rect 20805 9346 20871 9349
rect 24117 9346 24183 9349
rect 20805 9344 24183 9346
rect 20805 9288 20810 9344
rect 20866 9288 24122 9344
rect 24178 9288 24183 9344
rect 20805 9286 24183 9288
rect 20805 9283 20871 9286
rect 24117 9283 24183 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 21081 9210 21147 9213
rect 23933 9210 23999 9213
rect 21081 9208 23999 9210
rect 21081 9152 21086 9208
rect 21142 9152 23938 9208
rect 23994 9152 23999 9208
rect 21081 9150 23999 9152
rect 21081 9147 21147 9150
rect 23933 9147 23999 9150
rect 9121 9074 9187 9077
rect 12157 9074 12223 9077
rect 9121 9072 12223 9074
rect 9121 9016 9126 9072
rect 9182 9016 12162 9072
rect 12218 9016 12223 9072
rect 9121 9014 12223 9016
rect 9121 9011 9187 9014
rect 12157 9011 12223 9014
rect 24209 9074 24275 9077
rect 27520 9074 28000 9104
rect 24209 9072 28000 9074
rect 24209 9016 24214 9072
rect 24270 9016 28000 9072
rect 24209 9014 28000 9016
rect 24209 9011 24275 9014
rect 27520 8984 28000 9014
rect 21081 8938 21147 8941
rect 24669 8938 24735 8941
rect 21081 8936 24735 8938
rect 21081 8880 21086 8936
rect 21142 8880 24674 8936
rect 24730 8880 24735 8936
rect 21081 8878 24735 8880
rect 21081 8875 21147 8878
rect 24669 8875 24735 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 11237 8530 11303 8533
rect 21909 8530 21975 8533
rect 11237 8528 21975 8530
rect 11237 8472 11242 8528
rect 11298 8472 21914 8528
rect 21970 8472 21975 8528
rect 11237 8470 21975 8472
rect 11237 8467 11303 8470
rect 21909 8467 21975 8470
rect 24853 8530 24919 8533
rect 27520 8530 28000 8560
rect 24853 8528 28000 8530
rect 24853 8472 24858 8528
rect 24914 8472 28000 8528
rect 24853 8470 28000 8472
rect 24853 8467 24919 8470
rect 27520 8440 28000 8470
rect 13445 8394 13511 8397
rect 17953 8394 18019 8397
rect 13445 8392 18019 8394
rect 13445 8336 13450 8392
rect 13506 8336 17958 8392
rect 18014 8336 18019 8392
rect 13445 8334 18019 8336
rect 13445 8331 13511 8334
rect 17953 8331 18019 8334
rect 18137 8394 18203 8397
rect 20989 8394 21055 8397
rect 18137 8392 21055 8394
rect 18137 8336 18142 8392
rect 18198 8336 20994 8392
rect 21050 8336 21055 8392
rect 18137 8334 21055 8336
rect 18137 8331 18203 8334
rect 20989 8331 21055 8334
rect 12985 8258 13051 8261
rect 14181 8258 14247 8261
rect 16849 8258 16915 8261
rect 12985 8256 16915 8258
rect 12985 8200 12990 8256
rect 13046 8200 14186 8256
rect 14242 8200 16854 8256
rect 16910 8200 16915 8256
rect 12985 8198 16915 8200
rect 12985 8195 13051 8198
rect 14181 8195 14247 8198
rect 16849 8195 16915 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 12433 8122 12499 8125
rect 18045 8122 18111 8125
rect 12433 8120 18111 8122
rect 12433 8064 12438 8120
rect 12494 8064 18050 8120
rect 18106 8064 18111 8120
rect 12433 8062 18111 8064
rect 12433 8059 12499 8062
rect 18045 8059 18111 8062
rect 11973 7986 12039 7989
rect 12985 7986 13051 7989
rect 11973 7984 13051 7986
rect 11973 7928 11978 7984
rect 12034 7928 12990 7984
rect 13046 7928 13051 7984
rect 11973 7926 13051 7928
rect 11973 7923 12039 7926
rect 12985 7923 13051 7926
rect 13997 7986 14063 7989
rect 18137 7986 18203 7989
rect 13997 7984 18203 7986
rect 13997 7928 14002 7984
rect 14058 7928 18142 7984
rect 18198 7928 18203 7984
rect 13997 7926 18203 7928
rect 13997 7923 14063 7926
rect 18137 7923 18203 7926
rect 12525 7850 12591 7853
rect 16573 7850 16639 7853
rect 12525 7848 16639 7850
rect 12525 7792 12530 7848
rect 12586 7792 16578 7848
rect 16634 7792 16639 7848
rect 12525 7790 16639 7792
rect 12525 7787 12591 7790
rect 16573 7787 16639 7790
rect 18505 7850 18571 7853
rect 19977 7850 20043 7853
rect 24209 7850 24275 7853
rect 18505 7848 24275 7850
rect 18505 7792 18510 7848
rect 18566 7792 19982 7848
rect 20038 7792 24214 7848
rect 24270 7792 24275 7848
rect 18505 7790 24275 7792
rect 18505 7787 18571 7790
rect 19977 7787 20043 7790
rect 24209 7787 24275 7790
rect 24669 7850 24735 7853
rect 25589 7850 25655 7853
rect 27520 7850 28000 7880
rect 24669 7848 28000 7850
rect 24669 7792 24674 7848
rect 24730 7792 25594 7848
rect 25650 7792 28000 7848
rect 24669 7790 28000 7792
rect 24669 7787 24735 7790
rect 25589 7787 25655 7790
rect 27520 7760 28000 7790
rect 10869 7714 10935 7717
rect 13537 7714 13603 7717
rect 10869 7712 13603 7714
rect 10869 7656 10874 7712
rect 10930 7656 13542 7712
rect 13598 7656 13603 7712
rect 10869 7654 13603 7656
rect 10869 7651 10935 7654
rect 13537 7651 13603 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6361 7442 6427 7445
rect 12433 7442 12499 7445
rect 6361 7440 12499 7442
rect 6361 7384 6366 7440
rect 6422 7384 12438 7440
rect 12494 7384 12499 7440
rect 6361 7382 12499 7384
rect 6361 7379 6427 7382
rect 12433 7379 12499 7382
rect 13353 7442 13419 7445
rect 21265 7442 21331 7445
rect 13353 7440 21331 7442
rect 13353 7384 13358 7440
rect 13414 7384 21270 7440
rect 21326 7384 21331 7440
rect 13353 7382 21331 7384
rect 13353 7379 13419 7382
rect 21265 7379 21331 7382
rect 12801 7306 12867 7309
rect 19701 7306 19767 7309
rect 12801 7304 19767 7306
rect 12801 7248 12806 7304
rect 12862 7248 19706 7304
rect 19762 7248 19767 7304
rect 12801 7246 19767 7248
rect 12801 7243 12867 7246
rect 19701 7243 19767 7246
rect 23933 7306 23999 7309
rect 27520 7306 28000 7336
rect 23933 7304 28000 7306
rect 23933 7248 23938 7304
rect 23994 7248 28000 7304
rect 23933 7246 28000 7248
rect 23933 7243 23999 7246
rect 27520 7216 28000 7246
rect 12617 7170 12683 7173
rect 19333 7170 19399 7173
rect 12617 7168 19399 7170
rect 12617 7112 12622 7168
rect 12678 7112 19338 7168
rect 19394 7112 19399 7168
rect 12617 7110 19399 7112
rect 12617 7107 12683 7110
rect 19333 7107 19399 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 11145 6898 11211 6901
rect 15193 6898 15259 6901
rect 11145 6896 15259 6898
rect 11145 6840 11150 6896
rect 11206 6840 15198 6896
rect 15254 6840 15259 6896
rect 11145 6838 15259 6840
rect 11145 6835 11211 6838
rect 15193 6835 15259 6838
rect 16389 6898 16455 6901
rect 18505 6898 18571 6901
rect 16389 6896 18571 6898
rect 16389 6840 16394 6896
rect 16450 6840 18510 6896
rect 18566 6840 18571 6896
rect 16389 6838 18571 6840
rect 16389 6835 16455 6838
rect 18505 6835 18571 6838
rect 22093 6898 22159 6901
rect 25221 6898 25287 6901
rect 22093 6896 25287 6898
rect 22093 6840 22098 6896
rect 22154 6840 25226 6896
rect 25282 6840 25287 6896
rect 22093 6838 25287 6840
rect 22093 6835 22159 6838
rect 25221 6835 25287 6838
rect 3693 6762 3759 6765
rect 13445 6762 13511 6765
rect 3693 6760 13511 6762
rect 3693 6704 3698 6760
rect 3754 6704 13450 6760
rect 13506 6704 13511 6760
rect 3693 6702 13511 6704
rect 3693 6699 3759 6702
rect 13445 6699 13511 6702
rect 13629 6762 13695 6765
rect 15285 6762 15351 6765
rect 13629 6760 15351 6762
rect 13629 6704 13634 6760
rect 13690 6704 15290 6760
rect 15346 6704 15351 6760
rect 13629 6702 15351 6704
rect 13629 6699 13695 6702
rect 15285 6699 15351 6702
rect 18413 6762 18479 6765
rect 19149 6762 19215 6765
rect 27520 6762 28000 6792
rect 18413 6760 28000 6762
rect 18413 6704 18418 6760
rect 18474 6704 19154 6760
rect 19210 6704 28000 6760
rect 18413 6702 28000 6704
rect 18413 6699 18479 6702
rect 19149 6699 19215 6702
rect 27520 6672 28000 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 19057 6490 19123 6493
rect 21357 6490 21423 6493
rect 19057 6488 21423 6490
rect 19057 6432 19062 6488
rect 19118 6432 21362 6488
rect 21418 6432 21423 6488
rect 19057 6430 21423 6432
rect 19057 6427 19123 6430
rect 21357 6427 21423 6430
rect 2313 6354 2379 6357
rect 11789 6354 11855 6357
rect 2313 6352 11855 6354
rect 2313 6296 2318 6352
rect 2374 6296 11794 6352
rect 11850 6296 11855 6352
rect 2313 6294 11855 6296
rect 2313 6291 2379 6294
rect 11789 6291 11855 6294
rect 21633 6354 21699 6357
rect 24117 6354 24183 6357
rect 25313 6354 25379 6357
rect 21633 6352 25379 6354
rect 21633 6296 21638 6352
rect 21694 6296 24122 6352
rect 24178 6296 25318 6352
rect 25374 6296 25379 6352
rect 21633 6294 25379 6296
rect 21633 6291 21699 6294
rect 24117 6291 24183 6294
rect 25313 6291 25379 6294
rect 9029 6218 9095 6221
rect 16849 6218 16915 6221
rect 9029 6216 16915 6218
rect 9029 6160 9034 6216
rect 9090 6160 16854 6216
rect 16910 6160 16915 6216
rect 9029 6158 16915 6160
rect 9029 6155 9095 6158
rect 16849 6155 16915 6158
rect 12249 6082 12315 6085
rect 13629 6082 13695 6085
rect 27520 6082 28000 6112
rect 12249 6080 13695 6082
rect 12249 6024 12254 6080
rect 12310 6024 13634 6080
rect 13690 6024 13695 6080
rect 12249 6022 13695 6024
rect 12249 6019 12315 6022
rect 13629 6019 13695 6022
rect 22096 6022 28000 6082
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 13353 5946 13419 5949
rect 17309 5946 17375 5949
rect 22096 5946 22156 6022
rect 27520 5992 28000 6022
rect 13353 5944 17375 5946
rect 13353 5888 13358 5944
rect 13414 5888 17314 5944
rect 17370 5888 17375 5944
rect 13353 5886 17375 5888
rect 13353 5883 13419 5886
rect 17309 5883 17375 5886
rect 21958 5886 22156 5946
rect 15653 5810 15719 5813
rect 21958 5810 22018 5886
rect 15653 5808 22018 5810
rect 15653 5752 15658 5808
rect 15714 5752 22018 5808
rect 15653 5750 22018 5752
rect 15653 5747 15719 5750
rect 16297 5674 16363 5677
rect 20713 5674 20779 5677
rect 14782 5614 15394 5674
rect 5993 5538 6059 5541
rect 14782 5538 14842 5614
rect 5993 5536 14842 5538
rect 5993 5480 5998 5536
rect 6054 5480 14842 5536
rect 5993 5478 14842 5480
rect 15334 5538 15394 5614
rect 16297 5672 20779 5674
rect 16297 5616 16302 5672
rect 16358 5616 20718 5672
rect 20774 5616 20779 5672
rect 16297 5614 20779 5616
rect 16297 5611 16363 5614
rect 20713 5611 20779 5614
rect 22553 5674 22619 5677
rect 25405 5674 25471 5677
rect 22553 5672 25471 5674
rect 22553 5616 22558 5672
rect 22614 5616 25410 5672
rect 25466 5616 25471 5672
rect 22553 5614 25471 5616
rect 22553 5611 22619 5614
rect 25405 5611 25471 5614
rect 22829 5538 22895 5541
rect 15334 5536 22895 5538
rect 15334 5480 22834 5536
rect 22890 5480 22895 5536
rect 15334 5478 22895 5480
rect 5993 5475 6059 5478
rect 22829 5475 22895 5478
rect 24761 5538 24827 5541
rect 27520 5538 28000 5568
rect 24761 5536 28000 5538
rect 24761 5480 24766 5536
rect 24822 5480 28000 5536
rect 24761 5478 28000 5480
rect 24761 5475 24827 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 27520 5448 28000 5478
rect 24277 5407 24597 5408
rect 15745 5402 15811 5405
rect 16757 5402 16823 5405
rect 15745 5400 16823 5402
rect 15745 5344 15750 5400
rect 15806 5344 16762 5400
rect 16818 5344 16823 5400
rect 15745 5342 16823 5344
rect 15745 5339 15811 5342
rect 16757 5339 16823 5342
rect 15101 5266 15167 5269
rect 15837 5266 15903 5269
rect 16849 5266 16915 5269
rect 15101 5264 16915 5266
rect 15101 5208 15106 5264
rect 15162 5208 15842 5264
rect 15898 5208 16854 5264
rect 16910 5208 16915 5264
rect 15101 5206 16915 5208
rect 15101 5203 15167 5206
rect 15837 5203 15903 5206
rect 16849 5203 16915 5206
rect 19333 5266 19399 5269
rect 21725 5266 21791 5269
rect 19333 5264 21791 5266
rect 19333 5208 19338 5264
rect 19394 5208 21730 5264
rect 21786 5208 21791 5264
rect 19333 5206 21791 5208
rect 19333 5203 19399 5206
rect 21725 5203 21791 5206
rect 9765 5130 9831 5133
rect 16665 5130 16731 5133
rect 9765 5128 16731 5130
rect 9765 5072 9770 5128
rect 9826 5072 16670 5128
rect 16726 5072 16731 5128
rect 9765 5070 16731 5072
rect 9765 5067 9831 5070
rect 16665 5067 16731 5070
rect 17769 4994 17835 4997
rect 21173 4994 21239 4997
rect 27520 4994 28000 5024
rect 16254 4992 17835 4994
rect 16254 4936 17774 4992
rect 17830 4936 17835 4992
rect 16254 4934 17835 4936
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 0 4722 480 4752
rect 2865 4722 2931 4725
rect 0 4720 2931 4722
rect 0 4664 2870 4720
rect 2926 4664 2931 4720
rect 0 4662 2931 4664
rect 0 4632 480 4662
rect 2865 4659 2931 4662
rect 14733 4722 14799 4725
rect 15377 4722 15443 4725
rect 16254 4722 16314 4934
rect 17769 4931 17835 4934
rect 20302 4992 28000 4994
rect 20302 4936 21178 4992
rect 21234 4936 28000 4992
rect 20302 4934 28000 4936
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 16389 4858 16455 4861
rect 16389 4856 16498 4858
rect 16389 4800 16394 4856
rect 16450 4800 16498 4856
rect 16389 4795 16498 4800
rect 14733 4720 16314 4722
rect 14733 4664 14738 4720
rect 14794 4664 15382 4720
rect 15438 4664 16314 4720
rect 14733 4662 16314 4664
rect 14733 4659 14799 4662
rect 15377 4659 15443 4662
rect 10777 4586 10843 4589
rect 16297 4586 16363 4589
rect 10777 4584 16363 4586
rect 10777 4528 10782 4584
rect 10838 4528 16302 4584
rect 16358 4528 16363 4584
rect 10777 4526 16363 4528
rect 16438 4586 16498 4795
rect 18781 4722 18847 4725
rect 20302 4722 20362 4934
rect 21173 4931 21239 4934
rect 27520 4904 28000 4934
rect 18781 4720 20362 4722
rect 18781 4664 18786 4720
rect 18842 4664 20362 4720
rect 18781 4662 20362 4664
rect 18781 4659 18847 4662
rect 23565 4586 23631 4589
rect 16438 4584 23631 4586
rect 16438 4528 23570 4584
rect 23626 4528 23631 4584
rect 16438 4526 23631 4528
rect 10777 4523 10843 4526
rect 16297 4523 16363 4526
rect 23565 4523 23631 4526
rect 17493 4450 17559 4453
rect 19517 4450 19583 4453
rect 17493 4448 19583 4450
rect 17493 4392 17498 4448
rect 17554 4392 19522 4448
rect 19578 4392 19583 4448
rect 17493 4390 19583 4392
rect 17493 4387 17559 4390
rect 19517 4387 19583 4390
rect 19885 4450 19951 4453
rect 22277 4450 22343 4453
rect 19885 4448 22343 4450
rect 19885 4392 19890 4448
rect 19946 4392 22282 4448
rect 22338 4392 22343 4448
rect 19885 4390 22343 4392
rect 19885 4387 19951 4390
rect 22277 4387 22343 4390
rect 25221 4450 25287 4453
rect 27520 4450 28000 4480
rect 25221 4448 28000 4450
rect 25221 4392 25226 4448
rect 25282 4392 28000 4448
rect 25221 4390 28000 4392
rect 25221 4387 25287 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 16941 4314 17007 4317
rect 18689 4314 18755 4317
rect 16941 4312 18755 4314
rect 16941 4256 16946 4312
rect 17002 4256 18694 4312
rect 18750 4256 18755 4312
rect 16941 4254 18755 4256
rect 16941 4251 17007 4254
rect 18689 4251 18755 4254
rect 11697 4178 11763 4181
rect 14825 4178 14891 4181
rect 11697 4176 14891 4178
rect 11697 4120 11702 4176
rect 11758 4120 14830 4176
rect 14886 4120 14891 4176
rect 11697 4118 14891 4120
rect 11697 4115 11763 4118
rect 14825 4115 14891 4118
rect 17677 4178 17743 4181
rect 18413 4178 18479 4181
rect 21357 4178 21423 4181
rect 17677 4176 17970 4178
rect 17677 4120 17682 4176
rect 17738 4120 17970 4176
rect 17677 4118 17970 4120
rect 17677 4115 17743 4118
rect 7097 4042 7163 4045
rect 11237 4042 11303 4045
rect 7097 4040 11303 4042
rect 7097 3984 7102 4040
rect 7158 3984 11242 4040
rect 11298 3984 11303 4040
rect 7097 3982 11303 3984
rect 17910 4042 17970 4118
rect 18413 4176 21423 4178
rect 18413 4120 18418 4176
rect 18474 4120 21362 4176
rect 21418 4120 21423 4176
rect 18413 4118 21423 4120
rect 18413 4115 18479 4118
rect 21357 4115 21423 4118
rect 21541 4178 21607 4181
rect 21541 4176 24778 4178
rect 21541 4120 21546 4176
rect 21602 4120 24778 4176
rect 21541 4118 24778 4120
rect 21541 4115 21607 4118
rect 20989 4042 21055 4045
rect 17910 4040 21055 4042
rect 17910 3984 20994 4040
rect 21050 3984 21055 4040
rect 17910 3982 21055 3984
rect 7097 3979 7163 3982
rect 11237 3979 11303 3982
rect 20989 3979 21055 3982
rect 21541 4042 21607 4045
rect 23749 4042 23815 4045
rect 21541 4040 23815 4042
rect 21541 3984 21546 4040
rect 21602 3984 23754 4040
rect 23810 3984 23815 4040
rect 21541 3982 23815 3984
rect 24718 4042 24778 4118
rect 25313 4042 25379 4045
rect 24718 4040 25379 4042
rect 24718 3984 25318 4040
rect 25374 3984 25379 4040
rect 24718 3982 25379 3984
rect 21541 3979 21607 3982
rect 23749 3979 23815 3982
rect 25313 3979 25379 3982
rect 12433 3906 12499 3909
rect 15929 3906 15995 3909
rect 12433 3904 15995 3906
rect 12433 3848 12438 3904
rect 12494 3848 15934 3904
rect 15990 3848 15995 3904
rect 12433 3846 15995 3848
rect 12433 3843 12499 3846
rect 15929 3843 15995 3846
rect 24117 3906 24183 3909
rect 24117 3904 25514 3906
rect 24117 3848 24122 3904
rect 24178 3848 25514 3904
rect 24117 3846 25514 3848
rect 24117 3843 24183 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 15101 3770 15167 3773
rect 18137 3770 18203 3773
rect 15101 3768 18203 3770
rect 15101 3712 15106 3768
rect 15162 3712 18142 3768
rect 18198 3712 18203 3768
rect 15101 3710 18203 3712
rect 15101 3707 15167 3710
rect 18137 3707 18203 3710
rect 20897 3770 20963 3773
rect 25221 3770 25287 3773
rect 20897 3768 25287 3770
rect 20897 3712 20902 3768
rect 20958 3712 25226 3768
rect 25282 3712 25287 3768
rect 20897 3710 25287 3712
rect 25454 3770 25514 3846
rect 27520 3770 28000 3800
rect 25454 3710 28000 3770
rect 20897 3707 20963 3710
rect 25221 3707 25287 3710
rect 27520 3680 28000 3710
rect 14273 3634 14339 3637
rect 17769 3634 17835 3637
rect 7606 3632 17835 3634
rect 7606 3576 14278 3632
rect 14334 3576 17774 3632
rect 17830 3576 17835 3632
rect 7606 3574 17835 3576
rect 933 3498 999 3501
rect 1945 3498 2011 3501
rect 7606 3498 7666 3574
rect 14273 3571 14339 3574
rect 17769 3571 17835 3574
rect 20989 3634 21055 3637
rect 22093 3634 22159 3637
rect 20989 3632 22159 3634
rect 20989 3576 20994 3632
rect 21050 3576 22098 3632
rect 22154 3576 22159 3632
rect 20989 3574 22159 3576
rect 20989 3571 21055 3574
rect 22093 3571 22159 3574
rect 933 3496 2011 3498
rect 933 3440 938 3496
rect 994 3440 1950 3496
rect 2006 3440 2011 3496
rect 933 3438 2011 3440
rect 933 3435 999 3438
rect 1945 3435 2011 3438
rect 2086 3438 7666 3498
rect 12249 3498 12315 3501
rect 15377 3498 15443 3501
rect 12249 3496 15443 3498
rect 12249 3440 12254 3496
rect 12310 3440 15382 3496
rect 15438 3440 15443 3496
rect 12249 3438 15443 3440
rect 289 3362 355 3365
rect 2086 3362 2146 3438
rect 12249 3435 12315 3438
rect 15377 3435 15443 3438
rect 17217 3498 17283 3501
rect 19333 3498 19399 3501
rect 17217 3496 19399 3498
rect 17217 3440 17222 3496
rect 17278 3440 19338 3496
rect 19394 3440 19399 3496
rect 17217 3438 19399 3440
rect 17217 3435 17283 3438
rect 19333 3435 19399 3438
rect 22277 3498 22343 3501
rect 24117 3498 24183 3501
rect 22277 3496 24183 3498
rect 22277 3440 22282 3496
rect 22338 3440 24122 3496
rect 24178 3440 24183 3496
rect 22277 3438 24183 3440
rect 22277 3435 22343 3438
rect 24117 3435 24183 3438
rect 289 3360 2146 3362
rect 289 3304 294 3360
rect 350 3304 2146 3360
rect 289 3302 2146 3304
rect 18505 3362 18571 3365
rect 23657 3362 23723 3365
rect 18505 3360 23723 3362
rect 18505 3304 18510 3360
rect 18566 3304 23662 3360
rect 23718 3304 23723 3360
rect 18505 3302 23723 3304
rect 289 3299 355 3302
rect 18505 3299 18571 3302
rect 23657 3299 23723 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 15561 3226 15627 3229
rect 20713 3226 20779 3229
rect 23933 3226 23999 3229
rect 27520 3226 28000 3256
rect 15561 3224 20779 3226
rect 15561 3168 15566 3224
rect 15622 3168 20718 3224
rect 20774 3168 20779 3224
rect 15561 3166 20779 3168
rect 15561 3163 15627 3166
rect 20713 3163 20779 3166
rect 21958 3224 23999 3226
rect 21958 3168 23938 3224
rect 23994 3168 23999 3224
rect 21958 3166 23999 3168
rect 13537 3090 13603 3093
rect 16573 3090 16639 3093
rect 13537 3088 16639 3090
rect 13537 3032 13542 3088
rect 13598 3032 16578 3088
rect 16634 3032 16639 3088
rect 13537 3030 16639 3032
rect 13537 3027 13603 3030
rect 16573 3027 16639 3030
rect 16757 3090 16823 3093
rect 21958 3090 22018 3166
rect 23933 3163 23999 3166
rect 24718 3166 28000 3226
rect 16757 3088 22018 3090
rect 16757 3032 16762 3088
rect 16818 3032 22018 3088
rect 16757 3030 22018 3032
rect 24209 3090 24275 3093
rect 24718 3090 24778 3166
rect 27520 3136 28000 3166
rect 24209 3088 24778 3090
rect 24209 3032 24214 3088
rect 24270 3032 24778 3088
rect 24209 3030 24778 3032
rect 16757 3027 16823 3030
rect 24209 3027 24275 3030
rect 13629 2954 13695 2957
rect 17953 2954 18019 2957
rect 21541 2954 21607 2957
rect 13629 2952 18019 2954
rect 13629 2896 13634 2952
rect 13690 2896 17958 2952
rect 18014 2896 18019 2952
rect 13629 2894 18019 2896
rect 13629 2891 13695 2894
rect 17953 2891 18019 2894
rect 19382 2952 21607 2954
rect 19382 2896 21546 2952
rect 21602 2896 21607 2952
rect 19382 2894 21607 2896
rect 11421 2818 11487 2821
rect 15285 2818 15351 2821
rect 11421 2816 15351 2818
rect 11421 2760 11426 2816
rect 11482 2760 15290 2816
rect 15346 2760 15351 2816
rect 11421 2758 15351 2760
rect 11421 2755 11487 2758
rect 15285 2755 15351 2758
rect 15469 2818 15535 2821
rect 19382 2818 19442 2894
rect 21541 2891 21607 2894
rect 24761 2954 24827 2957
rect 27521 2954 27587 2957
rect 24761 2952 27587 2954
rect 24761 2896 24766 2952
rect 24822 2896 27526 2952
rect 27582 2896 27587 2952
rect 24761 2894 27587 2896
rect 24761 2891 24827 2894
rect 27521 2891 27587 2894
rect 15469 2816 19442 2818
rect 15469 2760 15474 2816
rect 15530 2760 19442 2816
rect 15469 2758 19442 2760
rect 23197 2818 23263 2821
rect 25497 2818 25563 2821
rect 23197 2816 25563 2818
rect 23197 2760 23202 2816
rect 23258 2760 25502 2816
rect 25558 2760 25563 2816
rect 23197 2758 25563 2760
rect 15469 2755 15535 2758
rect 23197 2755 23263 2758
rect 25497 2755 25563 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 23657 2682 23723 2685
rect 27520 2682 28000 2712
rect 23657 2680 28000 2682
rect 23657 2624 23662 2680
rect 23718 2624 28000 2680
rect 23657 2622 28000 2624
rect 23657 2619 23723 2622
rect 27520 2592 28000 2622
rect 12433 2546 12499 2549
rect 15929 2546 15995 2549
rect 12433 2544 15995 2546
rect 12433 2488 12438 2544
rect 12494 2488 15934 2544
rect 15990 2488 15995 2544
rect 12433 2486 15995 2488
rect 12433 2483 12499 2486
rect 15929 2483 15995 2486
rect 16205 2546 16271 2549
rect 22829 2546 22895 2549
rect 16205 2544 22895 2546
rect 16205 2488 16210 2544
rect 16266 2488 22834 2544
rect 22890 2488 22895 2544
rect 16205 2486 22895 2488
rect 16205 2483 16271 2486
rect 22829 2483 22895 2486
rect 4061 2410 4127 2413
rect 9029 2410 9095 2413
rect 4061 2408 9095 2410
rect 4061 2352 4066 2408
rect 4122 2352 9034 2408
rect 9090 2352 9095 2408
rect 4061 2350 9095 2352
rect 4061 2347 4127 2350
rect 9029 2347 9095 2350
rect 13629 2410 13695 2413
rect 16389 2410 16455 2413
rect 18321 2410 18387 2413
rect 13629 2408 16314 2410
rect 13629 2352 13634 2408
rect 13690 2352 16314 2408
rect 13629 2350 16314 2352
rect 13629 2347 13695 2350
rect 16254 2274 16314 2350
rect 16389 2408 18387 2410
rect 16389 2352 16394 2408
rect 16450 2352 18326 2408
rect 18382 2352 18387 2408
rect 16389 2350 18387 2352
rect 16389 2347 16455 2350
rect 18321 2347 18387 2350
rect 17217 2274 17283 2277
rect 16254 2272 17283 2274
rect 16254 2216 17222 2272
rect 17278 2216 17283 2272
rect 16254 2214 17283 2216
rect 17217 2211 17283 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 23565 2002 23631 2005
rect 27520 2002 28000 2032
rect 23565 2000 28000 2002
rect 23565 1944 23570 2000
rect 23626 1944 28000 2000
rect 23565 1942 28000 1944
rect 23565 1939 23631 1942
rect 27520 1912 28000 1942
rect 14457 1866 14523 1869
rect 21357 1866 21423 1869
rect 14457 1864 21423 1866
rect 14457 1808 14462 1864
rect 14518 1808 21362 1864
rect 21418 1808 21423 1864
rect 14457 1806 21423 1808
rect 14457 1803 14523 1806
rect 21357 1803 21423 1806
rect 13353 1730 13419 1733
rect 19425 1730 19491 1733
rect 13353 1728 19491 1730
rect 13353 1672 13358 1728
rect 13414 1672 19430 1728
rect 19486 1672 19491 1728
rect 13353 1670 19491 1672
rect 13353 1667 13419 1670
rect 19425 1667 19491 1670
rect 11605 1594 11671 1597
rect 15929 1594 15995 1597
rect 11605 1592 15995 1594
rect 11605 1536 11610 1592
rect 11666 1536 15934 1592
rect 15990 1536 15995 1592
rect 11605 1534 15995 1536
rect 11605 1531 11671 1534
rect 15929 1531 15995 1534
rect 19333 1594 19399 1597
rect 19333 1592 26986 1594
rect 19333 1536 19338 1592
rect 19394 1536 26986 1592
rect 19333 1534 26986 1536
rect 19333 1531 19399 1534
rect 10501 1458 10567 1461
rect 14549 1458 14615 1461
rect 10501 1456 14615 1458
rect 10501 1400 10506 1456
rect 10562 1400 14554 1456
rect 14610 1400 14615 1456
rect 10501 1398 14615 1400
rect 10501 1395 10567 1398
rect 14549 1395 14615 1398
rect 21909 1458 21975 1461
rect 26785 1458 26851 1461
rect 21909 1456 26851 1458
rect 21909 1400 21914 1456
rect 21970 1400 26790 1456
rect 26846 1400 26851 1456
rect 21909 1398 26851 1400
rect 26926 1458 26986 1534
rect 27520 1458 28000 1488
rect 26926 1398 28000 1458
rect 21909 1395 21975 1398
rect 26785 1395 26851 1398
rect 27520 1368 28000 1398
rect 21265 914 21331 917
rect 27520 914 28000 944
rect 21265 912 28000 914
rect 21265 856 21270 912
rect 21326 856 28000 912
rect 21265 854 28000 856
rect 21265 851 21331 854
rect 27520 824 28000 854
rect 25313 370 25379 373
rect 27520 370 28000 400
rect 25313 368 28000 370
rect 25313 312 25318 368
rect 25374 312 28000 368
rect 25313 310 28000 312
rect 25313 307 25379 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 14780 21796 14844 21860
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 14780 19408 14844 19412
rect 14780 19352 14830 19408
rect 14830 19352 14844 19408
rect 14780 19348 14844 19352
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 19380 18668 19444 18732
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 19380 11052 19444 11116
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14779 21860 14845 21861
rect 14779 21796 14780 21860
rect 14844 21796 14845 21860
rect 14779 21795 14845 21796
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 14782 19413 14842 21795
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14779 19412 14845 19413
rect 14779 19348 14780 19412
rect 14844 19348 14845 19412
rect 14779 19347 14845 19348
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 18528 15264 19552
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19379 18732 19445 18733
rect 19379 18668 19380 18732
rect 19444 18668 19445 18732
rect 19379 18667 19445 18668
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 19382 11117 19442 18667
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19379 11116 19445 11117
rect 19379 11052 19380 11116
rect 19444 11052 19445 11116
rect 19379 11051 19445 11052
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__buf_2  _059_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604666999
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604666999
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604666999
transform 1 0 5520 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604666999
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1604666999
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604666999
transform 1 0 8096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1604666999
transform 1 0 8004 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604666999
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604666999
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1604666999
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84
timestamp 1604666999
transform 1 0 8832 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1604666999
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604666999
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604666999
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1604666999
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604666999
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604666999
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1604666999
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604666999
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604666999
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604666999
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604666999
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604666999
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604666999
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1604666999
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604666999
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_130
timestamp 1604666999
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604666999
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604666999
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1604666999
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1604666999
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604666999
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604666999
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604666999
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604666999
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_139
timestamp 1604666999
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604666999
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604666999
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604666999
transform 1 0 15640 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 14536 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1604666999
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_160
timestamp 1604666999
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 15916 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170
timestamp 1604666999
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1604666999
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1604666999
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_174
timestamp 1604666999
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604666999
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1604666999
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604666999
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604666999
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18308 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_206
timestamp 1604666999
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1604666999
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_200
timestamp 1604666999
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604666999
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1604666999
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1604666999
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_212
timestamp 1604666999
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604666999
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20792 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_223
timestamp 1604666999
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1604666999
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1604666999
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604666999
transform 1 0 21712 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp 1604666999
transform 1 0 22356 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_232
timestamp 1604666999
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_228
timestamp 1604666999
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604666999
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_236
timestamp 1604666999
transform 1 0 22816 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604666999
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604666999
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_240
timestamp 1604666999
transform 1 0 23184 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604666999
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604666999
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1604666999
transform 1 0 24012 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23828 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604666999
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604666999
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604666999
transform 1 0 24564 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_267
timestamp 1604666999
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_263
timestamp 1604666999
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_259
timestamp 1604666999
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1604666999
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604666999
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_271
timestamp 1604666999
transform 1 0 26036 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_275
timestamp 1604666999
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_263
timestamp 1604666999
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 11500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1604666999
transform 1 0 10396 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_116
timestamp 1604666999
transform 1 0 11776 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604666999
transform 1 0 12512 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1604666999
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_132
timestamp 1604666999
transform 1 0 13248 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1604666999
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604666999
transform 1 0 15364 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604666999
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604666999
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16468 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1604666999
transform 1 0 15732 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_165
timestamp 1604666999
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18952 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1604666999
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1604666999
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp 1604666999
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1604666999
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 21988 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604666999
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_224
timestamp 1604666999
transform 1 0 21712 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_229
timestamp 1604666999
transform 1 0 22172 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_234
timestamp 1604666999
transform 1 0 22632 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23276 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24288 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_240
timestamp 1604666999
transform 1 0 23184 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1604666999
transform 1 0 24104 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_254
timestamp 1604666999
transform 1 0 24472 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604666999
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604666999
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604666999
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13340 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1604666999
transform 1 0 12788 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1604666999
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_156
timestamp 1604666999
transform 1 0 15456 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1604666999
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1604666999
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_180
timestamp 1604666999
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604666999
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604666999
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19596 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604666999
transform 1 0 22080 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604666999
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1604666999
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_224
timestamp 1604666999
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_232
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604666999
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604666999
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1604666999
transform 1 0 25392 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604666999
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1604666999
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1604666999
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12236 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604666999
transform 1 0 15548 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604666999
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_140
timestamp 1604666999
transform 1 0 13984 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_146
timestamp 1604666999
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604666999
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_161
timestamp 1604666999
transform 1 0 15916 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_165
timestamp 1604666999
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604666999
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_182
timestamp 1604666999
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1604666999
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1604666999
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1604666999
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604666999
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_234
timestamp 1604666999
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_238
timestamp 1604666999
transform 1 0 23000 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23368 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_261
timestamp 1604666999
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_273
timestamp 1604666999
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604666999
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604666999
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604666999
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604666999
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604666999
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604666999
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1604666999
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1604666999
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13984 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604666999
transform 1 0 16744 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604666999
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1604666999
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_163
timestamp 1604666999
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_167
timestamp 1604666999
transform 1 0 16468 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1604666999
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp 1604666999
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18400 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604666999
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604666999
transform 1 0 19964 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604666999
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_201
timestamp 1604666999
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_214
timestamp 1604666999
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1604666999
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604666999
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_222
timestamp 1604666999
transform 1 0 21528 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604666999
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23736 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604666999
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_265
timestamp 1604666999
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604666999
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604666999
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 1604666999
transform 1 0 11868 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604666999
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12144 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 13156 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1604666999
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_148
timestamp 1604666999
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_144
timestamp 1604666999
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1604666999
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1604666999
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_139
timestamp 1604666999
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_152
timestamp 1604666999
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15456 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 17020 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1604666999
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_167
timestamp 1604666999
transform 1 0 16468 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604666999
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604666999
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604666999
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604666999
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_196
timestamp 1604666999
transform 1 0 19136 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1604666999
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 19320 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18952 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19596 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_200
timestamp 1604666999
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604666999
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1604666999
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_224
timestamp 1604666999
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604666999
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1604666999
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604666999
transform 1 0 22080 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604666999
transform 1 0 22448 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1604666999
transform 1 0 22908 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_236
timestamp 1604666999
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1604666999
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_240
timestamp 1604666999
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23368 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23552 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1604666999
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1604666999
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 24196 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_260
timestamp 1604666999
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_264
timestamp 1604666999
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604666999
transform 1 0 25116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604666999
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_272
timestamp 1604666999
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_264
timestamp 1604666999
transform 1 0 25392 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604666999
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604666999
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_121
timestamp 1604666999
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1604666999
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1604666999
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604666999
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604666999
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_163
timestamp 1604666999
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_168
timestamp 1604666999
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_181
timestamp 1604666999
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp 1604666999
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_198
timestamp 1604666999
transform 1 0 19320 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21160 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1604666999
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_207
timestamp 1604666999
transform 1 0 20148 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_211
timestamp 1604666999
transform 1 0 20516 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 22724 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604666999
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_227
timestamp 1604666999
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1604666999
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_254
timestamp 1604666999
transform 1 0 24472 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25208 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1604666999
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_273
timestamp 1604666999
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604666999
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604666999
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604666999
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1604666999
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604666999
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604666999
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604666999
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1604666999
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1604666999
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_153
timestamp 1604666999
transform 1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1604666999
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1604666999
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604666999
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604666999
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_187
timestamp 1604666999
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_191
timestamp 1604666999
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_195
timestamp 1604666999
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 19412 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_218
timestamp 1604666999
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_222
timestamp 1604666999
transform 1 0 21528 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604666999
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604666999
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604666999
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604666999
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604666999
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1604666999
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604666999
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604666999
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1604666999
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1604666999
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_145
timestamp 1604666999
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_149
timestamp 1604666999
transform 1 0 14812 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604666999
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1604666999
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16560 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604666999
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1604666999
transform 1 0 16284 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1604666999
transform 1 0 17388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18124 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_183
timestamp 1604666999
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_194
timestamp 1604666999
transform 1 0 18952 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_198
timestamp 1604666999
transform 1 0 19320 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604666999
transform 1 0 19688 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1604666999
transform 1 0 19596 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_205
timestamp 1604666999
transform 1 0 19964 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_211
timestamp 1604666999
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 22632 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22448 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 1604666999
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_230
timestamp 1604666999
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1604666999
transform 1 0 24380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_257
timestamp 1604666999
transform 1 0 24748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 24932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_261
timestamp 1604666999
transform 1 0 25116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_273
timestamp 1604666999
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604666999
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604666999
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604666999
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604666999
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604666999
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_98
timestamp 1604666999
transform 1 0 10120 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604666999
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_104
timestamp 1604666999
transform 1 0 10672 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_107
timestamp 1604666999
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604666999
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604666999
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14904 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1604666999
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_146
timestamp 1604666999
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1604666999
transform 1 0 16652 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604666999
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604666999
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1604666999
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1604666999
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19964 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_201
timestamp 1604666999
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_224
timestamp 1604666999
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_228
timestamp 1604666999
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_235
timestamp 1604666999
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 24104 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_239
timestamp 1604666999
transform 1 0 23092 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604666999
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604666999
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604666999
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604666999
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604666999
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1604666999
transform 1 0 10028 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11132 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1604666999
transform 1 0 12880 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_145
timestamp 1604666999
transform 1 0 14444 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1604666999
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1604666999
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1604666999
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_190
timestamp 1604666999
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_194
timestamp 1604666999
transform 1 0 18952 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_198
timestamp 1604666999
transform 1 0 19320 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21068 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_202
timestamp 1604666999
transform 1 0 19688 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_207
timestamp 1604666999
transform 1 0 20148 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_211
timestamp 1604666999
transform 1 0 20516 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 22632 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_226
timestamp 1604666999
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_230
timestamp 1604666999
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24196 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_243
timestamp 1604666999
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_247
timestamp 1604666999
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_260
timestamp 1604666999
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_264
timestamp 1604666999
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_272
timestamp 1604666999
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_7
timestamp 1604666999
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_19
timestamp 1604666999
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604666999
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604666999
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604666999
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604666999
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9844 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1604666999
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604666999
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 11592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604666999
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1604666999
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_110
timestamp 1604666999
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_127
timestamp 1604666999
transform 1 0 12788 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1604666999
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1604666999
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1604666999
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1604666999
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14720 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_142
timestamp 1604666999
transform 1 0 14168 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_145
timestamp 1604666999
transform 1 0 14444 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1604666999
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1604666999
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1604666999
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1604666999
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604666999
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1604666999
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1604666999
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1604666999
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604666999
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1604666999
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604666999
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1604666999
transform 1 0 19228 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1604666999
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1604666999
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604666999
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1604666999
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1604666999
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20700 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604666999
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_226
timestamp 1604666999
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1604666999
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_235
timestamp 1604666999
transform 1 0 22724 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1604666999
transform 1 0 22080 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1604666999
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_230
timestamp 1604666999
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604666999
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23460 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 24104 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604666999
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604666999
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_262
timestamp 1604666999
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_266
timestamp 1604666999
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604666999
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_22
timestamp 1604666999
transform 1 0 3128 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_34
timestamp 1604666999
transform 1 0 4232 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_46
timestamp 1604666999
transform 1 0 5336 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1604666999
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604666999
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604666999
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_106
timestamp 1604666999
transform 1 0 10856 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604666999
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604666999
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604666999
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604666999
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15548 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1604666999
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1604666999
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_166
timestamp 1604666999
transform 1 0 16376 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_170
timestamp 1604666999
transform 1 0 16744 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1604666999
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18860 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_188
timestamp 1604666999
transform 1 0 18400 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1604666999
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1604666999
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21344 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1604666999
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_233
timestamp 1604666999
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1604666999
transform 1 0 22908 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1604666999
transform 1 0 23276 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604666999
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604666999
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_272
timestamp 1604666999
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604666999
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1604666999
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_19
timestamp 1604666999
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604666999
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604666999
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604666999
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604666999
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_105
timestamp 1604666999
transform 1 0 10764 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_113
timestamp 1604666999
transform 1 0 11500 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_117
timestamp 1604666999
transform 1 0 11868 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1604666999
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1604666999
transform 1 0 12604 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 1604666999
transform 1 0 12972 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1604666999
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604666999
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16836 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604666999
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1604666999
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_190
timestamp 1604666999
transform 1 0 18584 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_195
timestamp 1604666999
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1604666999
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604666999
transform 1 0 19780 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1604666999
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_210
timestamp 1604666999
transform 1 0 20424 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 20516 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604666999
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 22264 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_222
timestamp 1604666999
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_226
timestamp 1604666999
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24748 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_249
timestamp 1604666999
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1604666999
transform 1 0 24380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_266
timestamp 1604666999
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604666999
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604666999
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604666999
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604666999
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604666999
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604666999
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604666999
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_110
timestamp 1604666999
transform 1 0 11224 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1604666999
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1604666999
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13524 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604666999
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1604666999
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1604666999
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_154
timestamp 1604666999
transform 1 0 15272 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1604666999
transform 1 0 15732 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_163
timestamp 1604666999
transform 1 0 16100 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20516 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1604666999
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_207
timestamp 1604666999
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1604666999
transform 1 0 22264 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604666999
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604666999
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604666999
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_254
timestamp 1604666999
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_258
timestamp 1604666999
transform 1 0 24840 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_270
timestamp 1604666999
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604666999
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604666999
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604666999
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604666999
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604666999
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604666999
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_117
timestamp 1604666999
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_128
timestamp 1604666999
transform 1 0 12880 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15548 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604666999
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604666999
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1604666999
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604666999
transform 1 0 18032 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1604666999
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_187
timestamp 1604666999
transform 1 0 18308 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1604666999
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_196
timestamp 1604666999
transform 1 0 19136 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21068 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20516 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_206
timestamp 1604666999
transform 1 0 20056 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_210
timestamp 1604666999
transform 1 0 20424 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604666999
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 23000 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_236
timestamp 1604666999
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604666999
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1604666999
transform 1 0 23184 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_247
timestamp 1604666999
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_251
timestamp 1604666999
transform 1 0 24196 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_259
timestamp 1604666999
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1604666999
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604666999
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604666999
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604666999
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604666999
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604666999
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604666999
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604666999
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604666999
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604666999
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604666999
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604666999
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604666999
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604666999
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604666999
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1604666999
transform 1 0 12972 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 1604666999
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_137
timestamp 1604666999
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604666999
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 14076 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1604666999
transform 1 0 14076 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604666999
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1604666999
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1604666999
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1604666999
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 1604666999
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_176
timestamp 1604666999
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_171
timestamp 1604666999
transform 1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 17112 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1604666999
transform 1 0 18308 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_183
timestamp 1604666999
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1604666999
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1604666999
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1604666999
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18952 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1604666999
transform 1 0 20056 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1604666999
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1604666999
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604666999
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1604666999
transform 1 0 20424 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 20516 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20516 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_228
timestamp 1604666999
transform 1 0 22080 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_224
timestamp 1604666999
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_224
timestamp 1604666999
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_220
timestamp 1604666999
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22080 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_232
timestamp 1604666999
transform 1 0 22448 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_237
timestamp 1604666999
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_231
timestamp 1604666999
transform 1 0 22356 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22264 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604666999
transform 1 0 22724 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_244
timestamp 1604666999
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_241
timestamp 1604666999
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23736 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23092 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_254
timestamp 1604666999
transform 1 0 24472 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_248
timestamp 1604666999
transform 1 0 23920 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604666999
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604666999
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604666999
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1604666999
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604666999
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604666999
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_275
timestamp 1604666999
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604666999
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_263
timestamp 1604666999
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604666999
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604666999
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604666999
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604666999
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604666999
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604666999
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604666999
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1604666999
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1604666999
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1604666999
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14628 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1604666999
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1604666999
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15640 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1604666999
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1604666999
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_175
timestamp 1604666999
transform 1 0 17204 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1604666999
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1604666999
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19596 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604666999
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604666999
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_220
timestamp 1604666999
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_224
timestamp 1604666999
transform 1 0 21712 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_229
timestamp 1604666999
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604666999
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604666999
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604666999
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1604666999
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_268
timestamp 1604666999
transform 1 0 25760 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604666999
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604666999
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604666999
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604666999
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604666999
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604666999
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604666999
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604666999
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 13064 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_129
timestamp 1604666999
transform 1 0 12972 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_133
timestamp 1604666999
transform 1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604666999
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_145
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16008 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_160
timestamp 1604666999
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19044 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_181
timestamp 1604666999
transform 1 0 17756 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_186
timestamp 1604666999
transform 1 0 18216 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1604666999
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_204
timestamp 1604666999
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1604666999
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21988 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1604666999
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1604666999
transform 1 0 21620 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_230
timestamp 1604666999
transform 1 0 22264 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604666999
transform 1 0 24748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604666999
transform 1 0 23184 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_249
timestamp 1604666999
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_261
timestamp 1604666999
transform 1 0 25116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_273
timestamp 1604666999
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604666999
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604666999
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604666999
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604666999
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604666999
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604666999
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12972 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604666999
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_136
timestamp 1604666999
transform 1 0 13616 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604666999
transform 1 0 15180 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1604666999
transform 1 0 14168 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1604666999
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1604666999
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1604666999
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_160
timestamp 1604666999
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_173
timestamp 1604666999
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1604666999
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18492 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_208
timestamp 1604666999
transform 1 0 20240 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_216
timestamp 1604666999
transform 1 0 20976 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604666999
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21436 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604666999
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1604666999
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_228
timestamp 1604666999
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604666999
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604666999
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604666999
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1604666999
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604666999
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1604666999
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_263
timestamp 1604666999
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_275
timestamp 1604666999
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604666999
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604666999
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604666999
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604666999
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604666999
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604666999
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604666999
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604666999
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1604666999
transform 1 0 14076 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_144
timestamp 1604666999
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1604666999
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 17112 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_166
timestamp 1604666999
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1604666999
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604666999
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1604666999
transform 1 0 19228 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604666999
transform 1 0 19596 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_204
timestamp 1604666999
transform 1 0 19872 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1604666999
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1604666999
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21344 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1604666999
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604666999
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604666999
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_251
timestamp 1604666999
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_259
timestamp 1604666999
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604666999
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604666999
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604666999
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604666999
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604666999
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_98
timestamp 1604666999
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604666999
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_106
timestamp 1604666999
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604666999
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604666999
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_126
timestamp 1604666999
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_130
timestamp 1604666999
transform 1 0 13064 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_136
timestamp 1604666999
transform 1 0 13616 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1604666999
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1604666999
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_160
timestamp 1604666999
transform 1 0 15824 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604666999
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18584 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604666999
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20148 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_199
timestamp 1604666999
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1604666999
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_216
timestamp 1604666999
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21712 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1604666999
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1604666999
transform 1 0 22540 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1604666999
transform 1 0 22908 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604666999
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_241
timestamp 1604666999
transform 1 0 23276 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_249
timestamp 1604666999
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_253
timestamp 1604666999
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604666999
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604666999
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_259
timestamp 1604666999
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_263
timestamp 1604666999
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_267
timestamp 1604666999
transform 1 0 25668 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1604666999
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604666999
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604666999
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604666999
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604666999
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604666999
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604666999
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604666999
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_98
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1604666999
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_107
timestamp 1604666999
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604666999
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604666999
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1604666999
transform 1 0 11316 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_120
timestamp 1604666999
transform 1 0 12144 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1604666999
transform 1 0 12604 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_137
timestamp 1604666999
transform 1 0 13708 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1604666999
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1604666999
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_145
timestamp 1604666999
transform 1 0 14444 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1604666999
transform 1 0 14076 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604666999
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1604666999
transform 1 0 14812 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14904 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16836 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1604666999
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_168
timestamp 1604666999
transform 1 0 16560 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1604666999
transform 1 0 16652 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_174
timestamp 1604666999
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1604666999
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 18584 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1604666999
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_194
timestamp 1604666999
transform 1 0 18952 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604666999
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1604666999
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_202
timestamp 1604666999
transform 1 0 19688 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604666999
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1604666999
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1604666999
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604666999
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 21068 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_226
timestamp 1604666999
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1604666999
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_234
timestamp 1604666999
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_234
timestamp 1604666999
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1604666999
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_238
timestamp 1604666999
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23368 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_251
timestamp 1604666999
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_255
timestamp 1604666999
transform 1 0 24564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1604666999
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604666999
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604666999
transform 1 0 24932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604666999
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_268
timestamp 1604666999
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604666999
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604666999
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604666999
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11224 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_107
timestamp 1604666999
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_129
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_135
timestamp 1604666999
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_138
timestamp 1604666999
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604666999
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604666999
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1604666999
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16928 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1604666999
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1604666999
transform 1 0 16468 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_171
timestamp 1604666999
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_191
timestamp 1604666999
transform 1 0 18676 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_196
timestamp 1604666999
transform 1 0 19136 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19780 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_202
timestamp 1604666999
transform 1 0 19688 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604666999
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1604666999
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 22264 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1604666999
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1604666999
transform 1 0 22080 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_232
timestamp 1604666999
transform 1 0 22448 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604666999
transform 1 0 24748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23184 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1604666999
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1604666999
transform 1 0 24380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_261
timestamp 1604666999
transform 1 0 25116 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1604666999
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604666999
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604666999
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_86
timestamp 1604666999
transform 1 0 9016 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_94
timestamp 1604666999
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604666999
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604666999
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12788 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604666999
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 14352 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_140
timestamp 1604666999
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1604666999
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_167
timestamp 1604666999
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_174
timestamp 1604666999
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_178
timestamp 1604666999
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18952 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18768 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17664 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604666999
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1604666999
transform 1 0 18400 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1604666999
transform 1 0 20700 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1604666999
transform 1 0 21068 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21436 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_220
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_230
timestamp 1604666999
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_234
timestamp 1604666999
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_238
timestamp 1604666999
transform 1 0 23000 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1604666999
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604666999
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604666999
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1604666999
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1604666999
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_270
timestamp 1604666999
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604666999
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604666999
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604666999
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_99
timestamp 1604666999
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10672 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604666999
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1604666999
transform 1 0 12420 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_129
timestamp 1604666999
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_133
timestamp 1604666999
transform 1 0 13340 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1604666999
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1604666999
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 17112 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_164
timestamp 1604666999
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1604666999
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1604666999
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1604666999
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1604666999
transform 1 0 19228 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 21160 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19412 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1604666999
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_206
timestamp 1604666999
transform 1 0 20056 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604666999
transform 1 0 22816 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 22540 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_227
timestamp 1604666999
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1604666999
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_235
timestamp 1604666999
transform 1 0 22724 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23828 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_239
timestamp 1604666999
transform 1 0 23092 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_266
timestamp 1604666999
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604666999
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604666999
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604666999
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604666999
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_86
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1604666999
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_96
timestamp 1604666999
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1604666999
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1604666999
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604666999
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_136
timestamp 1604666999
transform 1 0 13616 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14168 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16652 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1604666999
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_165
timestamp 1604666999
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1604666999
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_176
timestamp 1604666999
transform 1 0 17296 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604666999
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1604666999
transform 1 0 18860 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1604666999
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19688 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1604666999
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp 1604666999
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21252 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_228
timestamp 1604666999
transform 1 0 22080 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_232
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604666999
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23920 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604666999
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_257
timestamp 1604666999
transform 1 0 24748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604666999
transform 1 0 25484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604666999
transform 1 0 26036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1604666999
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_269
timestamp 1604666999
transform 1 0 25852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_273
timestamp 1604666999
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A
timestamp 1604666999
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1604666999
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_19
timestamp 1604666999
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604666999
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604666999
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10212 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604666999
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_118
timestamp 1604666999
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12696 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_122
timestamp 1604666999
transform 1 0 12328 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1604666999
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15456 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14720 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_145
timestamp 1604666999
transform 1 0 14444 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1604666999
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_154
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1604666999
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18676 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1604666999
transform 1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1604666999
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_186
timestamp 1604666999
transform 1 0 18216 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_200
timestamp 1604666999
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_204
timestamp 1604666999
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_208
timestamp 1604666999
transform 1 0 20240 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604666999
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_234
timestamp 1604666999
transform 1 0 22632 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23920 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604666999
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A
timestamp 1604666999
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604666999
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_11
timestamp 1604666999
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_7
timestamp 1604666999
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_19
timestamp 1604666999
transform 1 0 2852 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_23
timestamp 1604666999
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_35
timestamp 1604666999
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_47
timestamp 1604666999
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604666999
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604666999
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604666999
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604666999
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604666999
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_98
timestamp 1604666999
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_107
timestamp 1604666999
transform 1 0 10948 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_103
timestamp 1604666999
transform 1 0 10580 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604666999
transform 1 0 10304 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_111
timestamp 1604666999
transform 1 0 11316 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604666999
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604666999
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604666999
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11408 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_135
timestamp 1604666999
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_131
timestamp 1604666999
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1604666999
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604666999
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_142
timestamp 1604666999
transform 1 0 14168 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1604666999
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp 1604666999
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604666999
transform 1 0 13892 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1604666999
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14904 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15364 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14720 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_34_164
timestamp 1604666999
transform 1 0 16192 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_167
timestamp 1604666999
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_172
timestamp 1604666999
transform 1 0 16928 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604666999
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1604666999
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17112 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 17296 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18860 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604666999
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1604666999
transform 1 0 18124 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1604666999
transform 1 0 18492 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_192
timestamp 1604666999
transform 1 0 18768 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1604666999
transform 1 0 20056 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_202
timestamp 1604666999
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1604666999
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1604666999
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19872 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604666999
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1604666999
transform 1 0 20424 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20516 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604666999
transform 1 0 20516 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_227
timestamp 1604666999
transform 1 0 21988 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_224
timestamp 1604666999
transform 1 0 21712 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1604666999
transform 1 0 21344 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_236
timestamp 1604666999
transform 1 0 22816 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_231
timestamp 1604666999
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22172 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604666999
transform 1 0 22540 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21804 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_244
timestamp 1604666999
transform 1 0 23552 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23736 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_248
timestamp 1604666999
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1604666999
transform 1 0 24104 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24288 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_267
timestamp 1604666999
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_263
timestamp 1604666999
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_259
timestamp 1604666999
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1604666999
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_271
timestamp 1604666999
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_261
timestamp 1604666999
transform 1 0 25116 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604666999
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604666999
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604666999
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604666999
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604666999
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_98
timestamp 1604666999
transform 1 0 10120 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_102
timestamp 1604666999
transform 1 0 10488 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604666999
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1604666999
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1604666999
transform 1 0 13616 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604666999
transform 1 0 14904 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_142
timestamp 1604666999
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_146
timestamp 1604666999
transform 1 0 14536 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604666999
transform 1 0 16928 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_159
timestamp 1604666999
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_163
timestamp 1604666999
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_167
timestamp 1604666999
transform 1 0 16468 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604666999
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 19044 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604666999
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_187
timestamp 1604666999
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_191
timestamp 1604666999
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_214
timestamp 1604666999
transform 1 0 20792 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1604666999
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_223
timestamp 1604666999
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_236
timestamp 1604666999
transform 1 0 22816 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 24104 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23920 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23092 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_241
timestamp 1604666999
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_245
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604666999
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604666999
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604666999
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604666999
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604666999
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604666999
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604666999
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 12052 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_107
timestamp 1604666999
transform 1 0 10948 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12880 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1604666999
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_125
timestamp 1604666999
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_137
timestamp 1604666999
transform 1 0 13708 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 15364 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 14904 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1604666999
transform 1 0 14076 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1604666999
transform 1 0 14812 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1604666999
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_154
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16928 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_164
timestamp 1604666999
transform 1 0 16192 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18584 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18400 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_181
timestamp 1604666999
transform 1 0 17756 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_186
timestamp 1604666999
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21068 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20148 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_199
timestamp 1604666999
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1604666999
transform 1 0 19780 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_209
timestamp 1604666999
transform 1 0 20332 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22080 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21528 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22908 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 22540 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_220
timestamp 1604666999
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_224
timestamp 1604666999
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_231
timestamp 1604666999
transform 1 0 22356 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_235
timestamp 1604666999
transform 1 0 22724 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23092 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1604666999
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1604666999
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1604666999
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604666999
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604666999
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604666999
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604666999
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604666999
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604666999
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_98
timestamp 1604666999
transform 1 0 10120 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_102
timestamp 1604666999
transform 1 0 10488 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_105
timestamp 1604666999
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_109
timestamp 1604666999
transform 1 0 11132 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_117
timestamp 1604666999
transform 1 0 11868 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604666999
transform 1 0 14904 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1604666999
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1604666999
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604666999
transform 1 0 16836 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604666999
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_159
timestamp 1604666999
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_163
timestamp 1604666999
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_167
timestamp 1604666999
transform 1 0 16468 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604666999
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604666999
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_193
timestamp 1604666999
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1604666999
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20148 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19964 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1604666999
transform 1 0 19596 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 22080 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_226
timestamp 1604666999
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1604666999
transform 1 0 22264 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1604666999
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604666999
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604666999
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_254
timestamp 1604666999
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604666999
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_258
timestamp 1604666999
transform 1 0 24840 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_266
timestamp 1604666999
transform 1 0 25576 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_274
timestamp 1604666999
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604666999
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604666999
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604666999
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604666999
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604666999
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604666999
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_93
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10580 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_38_101
timestamp 1604666999
transform 1 0 10396 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13064 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_122
timestamp 1604666999
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1604666999
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_143
timestamp 1604666999
transform 1 0 14260 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_139
timestamp 1604666999
transform 1 0 13892 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14076 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1604666999
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_149
timestamp 1604666999
transform 1 0 14812 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 14904 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_158
timestamp 1604666999
transform 1 0 15640 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15732 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_38_178
timestamp 1604666999
transform 1 0 17480 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 18216 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 17664 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_182
timestamp 1604666999
transform 1 0 17848 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1604666999
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1604666999
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23000 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_224
timestamp 1604666999
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_228
timestamp 1604666999
transform 1 0 22080 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_236
timestamp 1604666999
transform 1 0 22816 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604666999
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 24012 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_247
timestamp 1604666999
transform 1 0 23828 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_251
timestamp 1604666999
transform 1 0 24196 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1604666999
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1604666999
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604666999
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604666999
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604666999
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604666999
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604666999
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604666999
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604666999
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_98
timestamp 1604666999
transform 1 0 10120 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604666999
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_109
timestamp 1604666999
transform 1 0 11132 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_105
timestamp 1604666999
transform 1 0 10764 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_106
timestamp 1604666999
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_112
timestamp 1604666999
transform 1 0 11408 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604666999
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604666999
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604666999
transform 1 0 11224 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11776 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604666999
transform 1 0 11224 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604666999
transform 1 0 13340 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13156 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_125
timestamp 1604666999
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_129
timestamp 1604666999
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_142
timestamp 1604666999
transform 1 0 14168 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_146
timestamp 1604666999
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1604666999
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_158
timestamp 1604666999
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1604666999
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 14904 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15456 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1604666999
transform 1 0 14904 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_39_167
timestamp 1604666999
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_163
timestamp 1604666999
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1604666999
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15824 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1604666999
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_169
timestamp 1604666999
transform 1 0 16652 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_175
timestamp 1604666999
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604666999
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604666999
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_184
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604666999
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 17572 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18308 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 17756 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_40_195
timestamp 1604666999
transform 1 0 19044 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_190
timestamp 1604666999
transform 1 0 18584 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_189
timestamp 1604666999
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18860 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604666999
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18860 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604666999
transform 1 0 19596 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604666999
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1604666999
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1604666999
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_205
timestamp 1604666999
transform 1 0 19964 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1604666999
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_227
timestamp 1604666999
transform 1 0 21988 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_223
timestamp 1604666999
transform 1 0 21620 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 21804 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21344 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604666999
transform 1 0 21252 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_235
timestamp 1604666999
transform 1 0 22724 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_233
timestamp 1604666999
transform 1 0 22540 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_229
timestamp 1604666999
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604666999
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604666999
transform 1 0 22356 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_245
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_241
timestamp 1604666999
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604666999
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_247
timestamp 1604666999
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1604666999
transform 1 0 24012 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604666999
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604666999
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604666999
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604666999
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604666999
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604666999
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604666999
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604666999
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604666999
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604666999
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604666999
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604666999
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604666999
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604666999
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604666999
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604666999
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604666999
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604666999
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604666999
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604666999
transform 1 0 13156 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604666999
transform 1 0 13708 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_135
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604666999
transform 1 0 14260 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15364 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604666999
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604666999
transform 1 0 14076 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_139
timestamp 1604666999
transform 1 0 13892 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_147
timestamp 1604666999
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_151
timestamp 1604666999
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604666999
transform 1 0 16928 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604666999
transform 1 0 16652 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1604666999
transform 1 0 16192 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_168
timestamp 1604666999
transform 1 0 16560 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_171
timestamp 1604666999
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_175
timestamp 1604666999
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_179
timestamp 1604666999
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_193
timestamp 1604666999
transform 1 0 18860 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604666999
transform 1 0 20976 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604666999
transform 1 0 19872 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604666999
transform 1 0 20424 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604666999
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_201
timestamp 1604666999
transform 1 0 19596 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_208
timestamp 1604666999
transform 1 0 20240 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_212
timestamp 1604666999
transform 1 0 20608 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604666999
transform 1 0 22172 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604666999
transform 1 0 21528 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604666999
transform 1 0 22724 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604666999
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_220
timestamp 1604666999
transform 1 0 21344 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_224
timestamp 1604666999
transform 1 0 21712 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_233
timestamp 1604666999
transform 1 0 22540 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_237
timestamp 1604666999
transform 1 0 22908 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1604666999
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_248
timestamp 1604666999
transform 1 0 23920 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_260
timestamp 1604666999
transform 1 0 25024 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_272
timestamp 1604666999
transform 1 0 26128 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_276
timestamp 1604666999
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604666999
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604666999
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604666999
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604666999
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604666999
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604666999
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604666999
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604666999
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604666999
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_137
timestamp 1604666999
transform 1 0 13708 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604666999
transform 1 0 15548 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604666999
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604666999
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_147
timestamp 1604666999
transform 1 0 14628 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_156
timestamp 1604666999
transform 1 0 15456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604666999
transform 1 0 16652 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16100 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_161
timestamp 1604666999
transform 1 0 15916 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1604666999
transform 1 0 16284 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_173
timestamp 1604666999
transform 1 0 17020 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_181
timestamp 1604666999
transform 1 0 17756 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604666999
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604666999
transform 1 0 19412 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_203
timestamp 1604666999
transform 1 0 19780 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_215
timestamp 1604666999
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_218
timestamp 1604666999
transform 1 0 21160 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604666999
transform 1 0 21988 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_226
timestamp 1604666999
transform 1 0 21896 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_231
timestamp 1604666999
transform 1 0 22356 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_243
timestamp 1604666999
transform 1 0 23460 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_247
timestamp 1604666999
transform 1 0 23828 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604666999
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604666999
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604666999
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 13880 480 14000 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 23264 480 23384 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 280 28000 400 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 824 28000 944 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 7746 27520 7802 28000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2962 27520 3018 28000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 5722 27520 5778 28000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 25502 27520 25558 28000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 26146 27520 26202 28000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 15290 27520 15346 28000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 17314 27520 17370 28000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 20718 27520 20774 28000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 prog_clk
port 123 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 right_top_grid_pin_42_
port 124 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 right_top_grid_pin_43_
port 125 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 126 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 127 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_top_grid_pin_46_
port 128 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 129 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 130 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 131 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
