magic
tech EFS8A
magscale 1 2
timestamp 1602269554
<< locali >>
rect 12173 18207 12207 18309
rect 14473 18207 14507 18377
rect 6319 17697 6354 17731
rect 8619 17697 8654 17731
rect 16347 17697 16382 17731
rect 18647 17697 18682 17731
rect 19107 17085 19142 17119
rect 8033 16031 8067 16201
rect 8953 14263 8987 14569
rect 13093 13855 13127 14025
rect 8947 13719 8981 13787
rect 8947 13685 8953 13719
rect 9999 13413 10044 13447
rect 6009 12835 6043 12937
rect 15853 12631 15887 12869
rect 4439 12393 4445 12427
rect 6187 12393 6193 12427
rect 4439 12325 4473 12393
rect 6187 12325 6221 12393
rect 6016 11237 6088 11271
rect 10091 11169 10218 11203
rect 1547 10217 1685 10251
rect 3007 8993 3042 9027
rect 5675 8993 5710 9027
rect 5175 8041 5181 8075
rect 5175 7973 5209 8041
rect 17240 7973 17312 8007
rect 12449 7327 12483 7497
rect 1771 7191 1805 7259
rect 14283 7191 14317 7259
rect 1771 7157 1777 7191
rect 14283 7157 14289 7191
rect 2783 6103 2817 6171
rect 2783 6069 2789 6103
rect 18423 5015 18457 5083
rect 18423 4981 18429 5015
rect 2973 4063 3007 4233
rect 14743 3927 14777 3995
rect 14743 3893 14749 3927
rect 17332 3621 17404 3655
rect 2697 2975 2731 3145
rect 12081 2907 12115 3145
rect 1547 2533 1685 2567
rect 6101 2363 6135 2601
rect 16037 2295 16071 2465
<< viali >>
rect 10287 19397 10321 19431
rect 10216 19261 10250 19295
rect 11228 19261 11262 19295
rect 13160 19261 13194 19295
rect 14156 19261 14190 19295
rect 10701 19125 10735 19159
rect 11299 19125 11333 19159
rect 11621 19125 11655 19159
rect 13231 19125 13265 19159
rect 13553 19125 13587 19159
rect 14243 19125 14277 19159
rect 14657 19125 14691 19159
rect 8620 18785 8654 18819
rect 10676 18785 10710 18819
rect 11656 18785 11690 18819
rect 13496 18785 13530 18819
rect 15368 18785 15402 18819
rect 8723 18581 8757 18615
rect 10747 18581 10781 18615
rect 11759 18581 11793 18615
rect 13599 18581 13633 18615
rect 15439 18581 15473 18615
rect 7481 18377 7515 18411
rect 10701 18377 10735 18411
rect 11989 18377 12023 18411
rect 14473 18377 14507 18411
rect 14749 18377 14783 18411
rect 8999 18309 9033 18343
rect 12173 18309 12207 18343
rect 15347 18309 15381 18343
rect 7297 18173 7331 18207
rect 8928 18173 8962 18207
rect 10184 18173 10218 18207
rect 10977 18173 11011 18207
rect 11212 18173 11246 18207
rect 11621 18173 11655 18207
rect 12173 18173 12207 18207
rect 14248 18173 14282 18207
rect 14473 18173 14507 18207
rect 15244 18173 15278 18207
rect 15669 18173 15703 18207
rect 18128 18173 18162 18207
rect 7941 18105 7975 18139
rect 10287 18105 10321 18139
rect 11299 18105 11333 18139
rect 14335 18105 14369 18139
rect 18521 18105 18555 18139
rect 8585 18037 8619 18071
rect 9413 18037 9447 18071
rect 12449 18037 12483 18071
rect 13461 18037 13495 18071
rect 16037 18037 16071 18071
rect 18199 18037 18233 18071
rect 13185 17833 13219 17867
rect 6285 17697 6319 17731
rect 7640 17697 7674 17731
rect 8585 17697 8619 17731
rect 11504 17697 11538 17731
rect 13369 17697 13403 17731
rect 13553 17697 13587 17731
rect 16313 17697 16347 17731
rect 17636 17697 17670 17731
rect 18613 17697 18647 17731
rect 19660 17697 19694 17731
rect 9689 17629 9723 17663
rect 15301 17629 15335 17663
rect 19763 17561 19797 17595
rect 6423 17493 6457 17527
rect 7711 17493 7745 17527
rect 8723 17493 8757 17527
rect 11575 17493 11609 17527
rect 12541 17493 12575 17527
rect 12817 17493 12851 17527
rect 14105 17493 14139 17527
rect 16451 17493 16485 17527
rect 17739 17493 17773 17527
rect 18061 17493 18095 17527
rect 18751 17493 18785 17527
rect 19073 17493 19107 17527
rect 6377 17289 6411 17323
rect 8677 17289 8711 17323
rect 10609 17289 10643 17323
rect 19211 17289 19245 17323
rect 19717 17289 19751 17323
rect 9275 17221 9309 17255
rect 11805 17221 11839 17255
rect 16313 17221 16347 17255
rect 7481 17153 7515 17187
rect 13001 17153 13035 17187
rect 17141 17153 17175 17187
rect 6996 17085 7030 17119
rect 8160 17085 8194 17119
rect 8953 17085 8987 17119
rect 9204 17085 9238 17119
rect 9597 17085 9631 17119
rect 10216 17085 10250 17119
rect 11380 17085 11414 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 14013 17085 14047 17119
rect 14473 17085 14507 17119
rect 16732 17085 16766 17119
rect 18096 17085 18130 17119
rect 19073 17085 19107 17119
rect 7757 17017 7791 17051
rect 8263 17017 8297 17051
rect 13921 17017 13955 17051
rect 16819 17017 16853 17051
rect 7067 16949 7101 16983
rect 10287 16949 10321 16983
rect 11483 16949 11517 16983
rect 13461 16949 13495 16983
rect 14289 16949 14323 16983
rect 15577 16949 15611 16983
rect 17601 16949 17635 16983
rect 18199 16949 18233 16983
rect 18705 16949 18739 16983
rect 8677 16745 8711 16779
rect 12357 16745 12391 16779
rect 13921 16745 13955 16779
rect 19257 16745 19291 16779
rect 10425 16677 10459 16711
rect 5248 16609 5282 16643
rect 6260 16609 6294 16643
rect 7272 16609 7306 16643
rect 8493 16609 8527 16643
rect 9689 16609 9723 16643
rect 12357 16609 12391 16643
rect 12633 16609 12667 16643
rect 13737 16609 13771 16643
rect 14105 16609 14139 16643
rect 15945 16609 15979 16643
rect 19073 16609 19107 16643
rect 10057 16541 10091 16575
rect 15301 16541 15335 16575
rect 16865 16541 16899 16575
rect 17877 16541 17911 16575
rect 9413 16473 9447 16507
rect 9827 16473 9861 16507
rect 5319 16405 5353 16439
rect 6331 16405 6365 16439
rect 7343 16405 7377 16439
rect 8309 16405 8343 16439
rect 9045 16405 9079 16439
rect 9965 16405 9999 16439
rect 13185 16405 13219 16439
rect 13461 16405 13495 16439
rect 6285 16201 6319 16235
rect 8033 16201 8067 16235
rect 8309 16201 8343 16235
rect 14841 16201 14875 16235
rect 19625 16201 19659 16235
rect 3663 16133 3697 16167
rect 1547 16065 1581 16099
rect 1961 16065 1995 16099
rect 4859 16065 4893 16099
rect 7297 16065 7331 16099
rect 8907 16133 8941 16167
rect 9045 16133 9079 16167
rect 9137 16065 9171 16099
rect 10241 16065 10275 16099
rect 13277 16065 13311 16099
rect 1460 15997 1494 16031
rect 2580 15997 2614 16031
rect 3592 15997 3626 16031
rect 4756 15997 4790 16031
rect 5181 15997 5215 16031
rect 5784 15997 5818 16031
rect 7824 15997 7858 16031
rect 8033 15997 8067 16031
rect 9873 15997 9907 16031
rect 10793 15997 10827 16031
rect 11345 15997 11379 16031
rect 12516 15997 12550 16031
rect 12909 15997 12943 16031
rect 13461 15997 13495 16031
rect 14013 15997 14047 16031
rect 16221 15997 16255 16031
rect 16497 15997 16531 16031
rect 19200 15997 19234 16031
rect 19993 15997 20027 16031
rect 5871 15929 5905 15963
rect 7665 15929 7699 15963
rect 8769 15929 8803 15963
rect 9505 15929 9539 15963
rect 10701 15929 10735 15963
rect 11529 15929 11563 15963
rect 14197 15929 14231 15963
rect 15393 15929 15427 15963
rect 16681 15929 16715 15963
rect 19303 15929 19337 15963
rect 2651 15861 2685 15895
rect 3065 15861 3099 15895
rect 4077 15861 4111 15895
rect 5549 15861 5583 15895
rect 6653 15861 6687 15895
rect 7895 15861 7929 15895
rect 8585 15861 8619 15895
rect 12081 15861 12115 15895
rect 12587 15861 12621 15895
rect 14473 15861 14507 15895
rect 15853 15861 15887 15895
rect 18153 15861 18187 15895
rect 5089 15657 5123 15691
rect 10793 15657 10827 15691
rect 15439 15657 15473 15691
rect 19257 15657 19291 15691
rect 8033 15589 8067 15623
rect 3008 15521 3042 15555
rect 5089 15521 5123 15555
rect 5365 15521 5399 15555
rect 6561 15521 6595 15555
rect 8217 15521 8251 15555
rect 9781 15521 9815 15555
rect 11437 15521 11471 15555
rect 13737 15521 13771 15555
rect 14013 15521 14047 15555
rect 15368 15521 15402 15555
rect 16313 15521 16347 15555
rect 16865 15521 16899 15555
rect 18096 15521 18130 15555
rect 19073 15521 19107 15555
rect 1409 15453 1443 15487
rect 9689 15453 9723 15487
rect 11345 15453 11379 15487
rect 14197 15453 14231 15487
rect 17049 15453 17083 15487
rect 9413 15385 9447 15419
rect 12449 15385 12483 15419
rect 3111 15317 3145 15351
rect 6929 15317 6963 15351
rect 9137 15317 9171 15351
rect 14473 15317 14507 15351
rect 16037 15317 16071 15351
rect 18199 15317 18233 15351
rect 2053 15113 2087 15147
rect 2605 15113 2639 15147
rect 8125 15113 8159 15147
rect 9781 15113 9815 15147
rect 14197 15113 14231 15147
rect 17417 15113 17451 15147
rect 17785 15113 17819 15147
rect 19165 15113 19199 15147
rect 13921 15045 13955 15079
rect 6469 14977 6503 15011
rect 8953 14977 8987 15011
rect 10977 14977 11011 15011
rect 14473 14977 14507 15011
rect 1409 14909 1443 14943
rect 2973 14909 3007 14943
rect 3157 14909 3191 14943
rect 4077 14909 4111 14943
rect 5273 14909 5307 14943
rect 5457 14909 5491 14943
rect 7113 14909 7147 14943
rect 7297 14909 7331 14943
rect 8677 14909 8711 14943
rect 8861 14909 8895 14943
rect 10149 14909 10183 14943
rect 10517 14909 10551 14943
rect 13553 14909 13587 14943
rect 15117 14909 15151 14943
rect 15853 14909 15887 14943
rect 16037 14909 16071 14943
rect 18061 14909 18095 14943
rect 18521 14909 18555 14943
rect 19660 14909 19694 14943
rect 20085 14909 20119 14943
rect 3065 14841 3099 14875
rect 6101 14841 6135 14875
rect 12909 14841 12943 14875
rect 13001 14841 13035 14875
rect 14565 14841 14599 14875
rect 15945 14841 15979 14875
rect 19763 14841 19797 14875
rect 1593 14773 1627 14807
rect 4537 14773 4571 14807
rect 4813 14773 4847 14807
rect 5089 14773 5123 14807
rect 6929 14773 6963 14807
rect 10057 14773 10091 14807
rect 11345 14773 11379 14807
rect 12725 14773 12759 14807
rect 15485 14773 15519 14807
rect 17049 14773 17083 14807
rect 18153 14773 18187 14807
rect 1685 14569 1719 14603
rect 6561 14569 6595 14603
rect 7941 14569 7975 14603
rect 8953 14569 8987 14603
rect 11345 14569 11379 14603
rect 12909 14569 12943 14603
rect 14473 14569 14507 14603
rect 16957 14569 16991 14603
rect 18521 14569 18555 14603
rect 2237 14433 2271 14467
rect 4813 14433 4847 14467
rect 5181 14433 5215 14467
rect 5365 14433 5399 14467
rect 6745 14433 6779 14467
rect 6929 14433 6963 14467
rect 8309 14433 8343 14467
rect 8585 14433 8619 14467
rect 5457 14365 5491 14399
rect 7481 14365 7515 14399
rect 8769 14365 8803 14399
rect 9873 14501 9907 14535
rect 13185 14501 13219 14535
rect 13737 14501 13771 14535
rect 15485 14501 15519 14535
rect 18153 14501 18187 14535
rect 11253 14433 11287 14467
rect 11713 14433 11747 14467
rect 16865 14433 16899 14467
rect 17417 14433 17451 14467
rect 18429 14433 18463 14467
rect 18981 14433 19015 14467
rect 9781 14365 9815 14399
rect 10057 14365 10091 14399
rect 13093 14365 13127 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 9045 14297 9079 14331
rect 10701 14297 10735 14331
rect 16313 14297 16347 14331
rect 2605 14229 2639 14263
rect 3157 14229 3191 14263
rect 8953 14229 8987 14263
rect 11161 14229 11195 14263
rect 3801 14025 3835 14059
rect 10149 14025 10183 14059
rect 12587 14025 12621 14059
rect 13001 14025 13035 14059
rect 13093 14025 13127 14059
rect 14381 14025 14415 14059
rect 15117 14025 15151 14059
rect 16589 14025 16623 14059
rect 2881 13957 2915 13991
rect 8125 13957 8159 13991
rect 9873 13957 9907 13991
rect 10977 13957 11011 13991
rect 12265 13957 12299 13991
rect 8493 13889 8527 13923
rect 10425 13889 10459 13923
rect 11437 13889 11471 13923
rect 14749 13957 14783 13991
rect 16911 13957 16945 13991
rect 1409 13821 1443 13855
rect 2789 13821 2823 13855
rect 3065 13821 3099 13855
rect 3525 13821 3559 13855
rect 4353 13821 4387 13855
rect 5273 13821 5307 13855
rect 5641 13821 5675 13855
rect 7297 13821 7331 13855
rect 7573 13821 7607 13855
rect 8585 13821 8619 13855
rect 12516 13821 12550 13855
rect 13093 13821 13127 13855
rect 13461 13821 13495 13855
rect 15853 13821 15887 13855
rect 16221 13821 16255 13855
rect 16819 13821 16853 13855
rect 18061 13821 18095 13855
rect 18521 13821 18555 13855
rect 19073 13821 19107 13855
rect 19660 13821 19694 13855
rect 20085 13821 20119 13855
rect 2237 13753 2271 13787
rect 5089 13753 5123 13787
rect 7757 13753 7791 13787
rect 10517 13753 10551 13787
rect 13782 13753 13816 13787
rect 15209 13753 15243 13787
rect 1593 13685 1627 13719
rect 2605 13685 2639 13719
rect 4629 13685 4663 13719
rect 5457 13685 5491 13719
rect 6469 13685 6503 13719
rect 8953 13685 8987 13719
rect 9505 13685 9539 13719
rect 11805 13685 11839 13719
rect 13277 13685 13311 13719
rect 17233 13685 17267 13719
rect 17785 13685 17819 13719
rect 18153 13685 18187 13719
rect 19763 13685 19797 13719
rect 1961 13481 1995 13515
rect 5181 13481 5215 13515
rect 5733 13481 5767 13515
rect 9505 13481 9539 13515
rect 12909 13481 12943 13515
rect 14335 13481 14369 13515
rect 18613 13481 18647 13515
rect 1409 13413 1443 13447
rect 3893 13413 3927 13447
rect 4261 13413 4295 13447
rect 8769 13413 8803 13447
rect 9045 13413 9079 13447
rect 9965 13413 9999 13447
rect 12310 13413 12344 13447
rect 13185 13413 13219 13447
rect 15117 13413 15151 13447
rect 15485 13413 15519 13447
rect 17411 13413 17445 13447
rect 18981 13413 19015 13447
rect 2421 13345 2455 13379
rect 2973 13345 3007 13379
rect 5733 13345 5767 13379
rect 6101 13345 6135 13379
rect 8309 13345 8343 13379
rect 8585 13345 8619 13379
rect 14232 13345 14266 13379
rect 17969 13345 18003 13379
rect 3157 13277 3191 13311
rect 4169 13277 4203 13311
rect 4445 13277 4479 13311
rect 6653 13277 6687 13311
rect 9689 13277 9723 13311
rect 11989 13277 12023 13311
rect 15393 13277 15427 13311
rect 16037 13277 16071 13311
rect 16773 13277 16807 13311
rect 17049 13277 17083 13311
rect 18889 13277 18923 13311
rect 19165 13277 19199 13311
rect 7389 13209 7423 13243
rect 2237 13141 2271 13175
rect 3433 13141 3467 13175
rect 7021 13141 7055 13175
rect 10609 13141 10643 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 18245 13141 18279 13175
rect 3985 12937 4019 12971
rect 4261 12937 4295 12971
rect 5917 12937 5951 12971
rect 6009 12937 6043 12971
rect 10149 12937 10183 12971
rect 13921 12937 13955 12971
rect 15301 12937 15335 12971
rect 17509 12937 17543 12971
rect 19625 12937 19659 12971
rect 10793 12869 10827 12903
rect 11253 12869 11287 12903
rect 15853 12869 15887 12903
rect 19993 12869 20027 12903
rect 2605 12801 2639 12835
rect 3065 12801 3099 12835
rect 5181 12801 5215 12835
rect 6009 12801 6043 12835
rect 6929 12801 6963 12835
rect 8493 12801 8527 12835
rect 12541 12801 12575 12835
rect 12817 12801 12851 12835
rect 13461 12801 13495 12835
rect 14381 12801 14415 12835
rect 1777 12733 1811 12767
rect 2053 12733 2087 12767
rect 9229 12733 9263 12767
rect 11412 12733 11446 12767
rect 15577 12733 15611 12767
rect 2973 12665 3007 12699
rect 3386 12665 3420 12699
rect 4905 12665 4939 12699
rect 4997 12665 5031 12699
rect 7021 12665 7055 12699
rect 7573 12665 7607 12699
rect 9550 12665 9584 12699
rect 11897 12665 11931 12699
rect 12633 12665 12667 12699
rect 14702 12665 14736 12699
rect 18705 12801 18739 12835
rect 18981 12801 19015 12835
rect 16129 12733 16163 12767
rect 16589 12733 16623 12767
rect 16865 12665 16899 12699
rect 18797 12665 18831 12699
rect 1593 12597 1627 12631
rect 4629 12597 4663 12631
rect 6285 12597 6319 12631
rect 6653 12597 6687 12631
rect 8125 12597 8159 12631
rect 9045 12597 9079 12631
rect 10425 12597 10459 12631
rect 11483 12597 11517 12631
rect 12173 12597 12207 12631
rect 14197 12597 14231 12631
rect 15853 12597 15887 12631
rect 15945 12597 15979 12631
rect 17141 12597 17175 12631
rect 18521 12597 18555 12631
rect 2237 12393 2271 12427
rect 3801 12393 3835 12427
rect 4445 12393 4479 12427
rect 5641 12393 5675 12427
rect 6193 12393 6227 12427
rect 6745 12393 6779 12427
rect 12909 12393 12943 12427
rect 14289 12393 14323 12427
rect 15117 12393 15151 12427
rect 17141 12393 17175 12427
rect 18245 12393 18279 12427
rect 1961 12325 1995 12359
rect 3157 12325 3191 12359
rect 8769 12325 8803 12359
rect 9229 12325 9263 12359
rect 9965 12325 9999 12359
rect 11707 12325 11741 12359
rect 15485 12325 15519 12359
rect 17647 12325 17681 12359
rect 18797 12325 18831 12359
rect 19257 12325 19291 12359
rect 1476 12257 1510 12291
rect 2421 12257 2455 12291
rect 2973 12257 3007 12291
rect 4077 12257 4111 12291
rect 5825 12257 5859 12291
rect 7021 12257 7055 12291
rect 8033 12257 8067 12291
rect 8585 12257 8619 12291
rect 10517 12257 10551 12291
rect 13185 12257 13219 12291
rect 13645 12257 13679 12291
rect 17325 12257 17359 12291
rect 9873 12189 9907 12223
rect 11345 12189 11379 12223
rect 13553 12189 13587 12223
rect 15393 12189 15427 12223
rect 16037 12189 16071 12223
rect 19165 12189 19199 12223
rect 19441 12189 19475 12223
rect 1547 12121 1581 12155
rect 3433 12053 3467 12087
rect 4997 12053 5031 12087
rect 5273 12053 5307 12087
rect 12265 12053 12299 12087
rect 12633 12053 12667 12087
rect 3157 11849 3191 11883
rect 4169 11849 4203 11883
rect 4905 11849 4939 11883
rect 6653 11849 6687 11883
rect 8861 11849 8895 11883
rect 9321 11849 9355 11883
rect 11253 11849 11287 11883
rect 13461 11849 13495 11883
rect 17325 11849 17359 11883
rect 17785 11849 17819 11883
rect 19257 11849 19291 11883
rect 4537 11781 4571 11815
rect 2421 11713 2455 11747
rect 3249 11713 3283 11747
rect 5365 11713 5399 11747
rect 6929 11713 6963 11747
rect 9873 11713 9907 11747
rect 10885 11713 10919 11747
rect 12541 11713 12575 11747
rect 14197 11713 14231 11747
rect 15669 11713 15703 11747
rect 18061 11713 18095 11747
rect 1961 11645 1995 11679
rect 2237 11645 2271 11679
rect 8125 11645 8159 11679
rect 11380 11645 11414 11679
rect 11805 11645 11839 11679
rect 16405 11645 16439 11679
rect 16589 11645 16623 11679
rect 19625 11645 19659 11679
rect 3570 11577 3604 11611
rect 5089 11577 5123 11611
rect 5181 11577 5215 11611
rect 7021 11577 7055 11611
rect 7573 11577 7607 11611
rect 9689 11577 9723 11611
rect 9965 11577 9999 11611
rect 10517 11577 10551 11611
rect 12633 11577 12667 11611
rect 13185 11577 13219 11611
rect 14518 11577 14552 11611
rect 16037 11577 16071 11611
rect 16865 11577 16899 11611
rect 18382 11577 18416 11611
rect 2697 11509 2731 11543
rect 6101 11509 6135 11543
rect 8401 11509 8435 11543
rect 11483 11509 11517 11543
rect 12173 11509 12207 11543
rect 14105 11509 14139 11543
rect 15117 11509 15151 11543
rect 18981 11509 19015 11543
rect 1593 11305 1627 11339
rect 2421 11305 2455 11339
rect 6929 11305 6963 11339
rect 9965 11305 9999 11339
rect 12541 11305 12575 11339
rect 13921 11305 13955 11339
rect 14289 11305 14323 11339
rect 15025 11305 15059 11339
rect 18061 11305 18095 11339
rect 18337 11305 18371 11339
rect 18705 11305 18739 11339
rect 4261 11237 4295 11271
rect 5982 11237 6016 11271
rect 7665 11237 7699 11271
rect 9505 11237 9539 11271
rect 11482 11237 11516 11271
rect 13093 11237 13127 11271
rect 15485 11237 15519 11271
rect 16037 11237 16071 11271
rect 17462 11237 17496 11271
rect 19073 11237 19107 11271
rect 2605 11169 2639 11203
rect 2789 11169 2823 11203
rect 7297 11169 7331 11203
rect 10057 11169 10091 11203
rect 11161 11169 11195 11203
rect 17141 11169 17175 11203
rect 4169 11101 4203 11135
rect 4813 11101 4847 11135
rect 5733 11101 5767 11135
rect 7573 11101 7607 11135
rect 7849 11101 7883 11135
rect 10701 11101 10735 11135
rect 13001 11101 13035 11135
rect 13277 11101 13311 11135
rect 15393 11101 15427 11135
rect 18981 11101 19015 11135
rect 19257 11101 19291 11135
rect 5181 11033 5215 11067
rect 2053 10965 2087 10999
rect 3433 10965 3467 10999
rect 3709 10965 3743 10999
rect 5457 10965 5491 10999
rect 6653 10965 6687 10999
rect 10287 10965 10321 10999
rect 12081 10965 12115 10999
rect 14657 10965 14691 10999
rect 2605 10761 2639 10795
rect 2973 10761 3007 10795
rect 4629 10761 4663 10795
rect 6653 10761 6687 10795
rect 9873 10761 9907 10795
rect 10517 10761 10551 10795
rect 12265 10761 12299 10795
rect 15393 10761 15427 10795
rect 17877 10761 17911 10795
rect 18337 10761 18371 10795
rect 19533 10761 19567 10795
rect 5825 10693 5859 10727
rect 8217 10693 8251 10727
rect 11345 10693 11379 10727
rect 13093 10693 13127 10727
rect 17049 10693 17083 10727
rect 3065 10625 3099 10659
rect 5089 10625 5123 10659
rect 5273 10625 5307 10659
rect 6929 10625 6963 10659
rect 7297 10625 7331 10659
rect 8953 10625 8987 10659
rect 10793 10625 10827 10659
rect 12541 10625 12575 10659
rect 14197 10625 14231 10659
rect 16497 10625 16531 10659
rect 18613 10625 18647 10659
rect 18889 10625 18923 10659
rect 19901 10625 19935 10659
rect 1685 10557 1719 10591
rect 2053 10557 2087 10591
rect 6285 10557 6319 10591
rect 15117 10557 15151 10591
rect 2237 10489 2271 10523
rect 3386 10489 3420 10523
rect 5365 10489 5399 10523
rect 7021 10489 7055 10523
rect 9274 10489 9308 10523
rect 10885 10489 10919 10523
rect 12633 10489 12667 10523
rect 14518 10489 14552 10523
rect 16313 10489 16347 10523
rect 16589 10489 16623 10523
rect 18705 10489 18739 10523
rect 3985 10421 4019 10455
rect 4261 10421 4295 10455
rect 7849 10421 7883 10455
rect 8861 10421 8895 10455
rect 10149 10421 10183 10455
rect 11713 10421 11747 10455
rect 13461 10421 13495 10455
rect 14105 10421 14139 10455
rect 15761 10421 15795 10455
rect 17417 10421 17451 10455
rect 1685 10217 1719 10251
rect 5733 10217 5767 10251
rect 7757 10217 7791 10251
rect 8953 10217 8987 10251
rect 11253 10217 11287 10251
rect 12541 10217 12575 10251
rect 12817 10217 12851 10251
rect 15577 10217 15611 10251
rect 16497 10217 16531 10251
rect 1961 10149 1995 10183
rect 3157 10149 3191 10183
rect 3433 10149 3467 10183
rect 4261 10149 4295 10183
rect 4813 10149 4847 10183
rect 6469 10149 6503 10183
rect 8033 10149 8067 10183
rect 9873 10149 9907 10183
rect 9965 10149 9999 10183
rect 11529 10149 11563 10183
rect 13185 10149 13219 10183
rect 13823 10149 13857 10183
rect 17094 10149 17128 10183
rect 18705 10149 18739 10183
rect 1476 10081 1510 10115
rect 2697 10081 2731 10115
rect 2973 10081 3007 10115
rect 13461 10081 13495 10115
rect 15669 10081 15703 10115
rect 16773 10081 16807 10115
rect 17693 10081 17727 10115
rect 2329 10013 2363 10047
rect 4169 10013 4203 10047
rect 6377 10013 6411 10047
rect 6653 10013 6687 10047
rect 7941 10013 7975 10047
rect 8217 10013 8251 10047
rect 10149 10013 10183 10047
rect 11437 10013 11471 10047
rect 11713 10013 11747 10047
rect 18613 10013 18647 10047
rect 18889 10013 18923 10047
rect 3801 9945 3835 9979
rect 15853 9945 15887 9979
rect 5273 9877 5307 9911
rect 6101 9877 6135 9911
rect 14381 9877 14415 9911
rect 4445 9673 4479 9707
rect 5917 9673 5951 9707
rect 9045 9673 9079 9707
rect 10425 9673 10459 9707
rect 11161 9673 11195 9707
rect 15761 9673 15795 9707
rect 16313 9673 16347 9707
rect 19073 9673 19107 9707
rect 6377 9605 6411 9639
rect 8585 9605 8619 9639
rect 10793 9605 10827 9639
rect 11437 9605 11471 9639
rect 13829 9605 13863 9639
rect 17049 9605 17083 9639
rect 19441 9605 19475 9639
rect 4997 9537 5031 9571
rect 7205 9537 7239 9571
rect 9505 9537 9539 9571
rect 12541 9537 12575 9571
rect 14565 9537 14599 9571
rect 16497 9537 16531 9571
rect 18153 9537 18187 9571
rect 18797 9537 18831 9571
rect 2145 9469 2179 9503
rect 2421 9469 2455 9503
rect 3249 9469 3283 9503
rect 3433 9469 3467 9503
rect 3893 9469 3927 9503
rect 7665 9469 7699 9503
rect 11253 9469 11287 9503
rect 11805 9469 11839 9503
rect 19692 9469 19726 9503
rect 20085 9469 20119 9503
rect 1777 9401 1811 9435
rect 2605 9401 2639 9435
rect 4169 9401 4203 9435
rect 4905 9401 4939 9435
rect 5359 9401 5393 9435
rect 7573 9401 7607 9435
rect 8027 9401 8061 9435
rect 9413 9401 9447 9435
rect 9867 9401 9901 9435
rect 12265 9401 12299 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 14657 9401 14691 9435
rect 15209 9401 15243 9435
rect 16589 9401 16623 9435
rect 18245 9401 18279 9435
rect 2973 9333 3007 9367
rect 13461 9333 13495 9367
rect 14381 9333 14415 9367
rect 17417 9333 17451 9367
rect 17785 9333 17819 9367
rect 19763 9333 19797 9367
rect 3433 9129 3467 9163
rect 5089 9129 5123 9163
rect 5549 9129 5583 9163
rect 7941 9129 7975 9163
rect 9965 9129 9999 9163
rect 11621 9129 11655 9163
rect 13553 9129 13587 9163
rect 14749 9129 14783 9163
rect 16497 9129 16531 9163
rect 17785 9129 17819 9163
rect 18153 9129 18187 9163
rect 1501 9061 1535 9095
rect 1593 9061 1627 9095
rect 2145 9061 2179 9095
rect 4261 9061 4295 9095
rect 4813 9061 4847 9095
rect 7383 9061 7417 9095
rect 10241 9061 10275 9095
rect 10609 9061 10643 9095
rect 10701 9061 10735 9095
rect 12265 9061 12299 9095
rect 12817 9061 12851 9095
rect 13737 9061 13771 9095
rect 13829 9061 13863 9095
rect 15025 9061 15059 9095
rect 15485 9061 15519 9095
rect 17227 9061 17261 9095
rect 18797 9061 18831 9095
rect 2973 8993 3007 9027
rect 5641 8993 5675 9027
rect 7021 8993 7055 9027
rect 8217 8993 8251 9027
rect 16865 8993 16899 9027
rect 3801 8925 3835 8959
rect 4169 8925 4203 8959
rect 11897 8925 11931 8959
rect 12173 8925 12207 8959
rect 15393 8925 15427 8959
rect 16037 8925 16071 8959
rect 18705 8925 18739 8959
rect 2881 8857 2915 8891
rect 6653 8857 6687 8891
rect 11161 8857 11195 8891
rect 14289 8857 14323 8891
rect 19257 8857 19291 8891
rect 2421 8789 2455 8823
rect 3111 8789 3145 8823
rect 5779 8789 5813 8823
rect 6377 8789 6411 8823
rect 1593 8585 1627 8619
rect 2697 8585 2731 8619
rect 3709 8585 3743 8619
rect 4169 8585 4203 8619
rect 6653 8585 6687 8619
rect 10241 8585 10275 8619
rect 10609 8585 10643 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 15393 8585 15427 8619
rect 17233 8585 17267 8619
rect 17877 8585 17911 8619
rect 18429 8585 18463 8619
rect 19625 8585 19659 8619
rect 8309 8517 8343 8551
rect 2789 8449 2823 8483
rect 4629 8449 4663 8483
rect 5273 8449 5307 8483
rect 7757 8449 7791 8483
rect 8677 8449 8711 8483
rect 9321 8449 9355 8483
rect 9965 8449 9999 8483
rect 10885 8449 10919 8483
rect 11161 8449 11195 8483
rect 15761 8449 15795 8483
rect 16037 8449 16071 8483
rect 18613 8449 18647 8483
rect 1409 8381 1443 8415
rect 5641 8381 5675 8415
rect 12817 8381 12851 8415
rect 13369 8381 13403 8415
rect 13921 8381 13955 8415
rect 3151 8313 3185 8347
rect 4721 8313 4755 8347
rect 7113 8313 7147 8347
rect 7849 8313 7883 8347
rect 9413 8313 9447 8347
rect 10977 8313 11011 8347
rect 14242 8313 14276 8347
rect 15853 8313 15887 8347
rect 18705 8313 18739 8347
rect 19257 8313 19291 8347
rect 2053 8245 2087 8279
rect 6009 8245 6043 8279
rect 7481 8245 7515 8279
rect 9045 8245 9079 8279
rect 12081 8245 12115 8279
rect 13737 8245 13771 8279
rect 14841 8245 14875 8279
rect 16957 8245 16991 8279
rect 1961 8041 1995 8075
rect 3433 8041 3467 8075
rect 4629 8041 4663 8075
rect 5181 8041 5215 8075
rect 9229 8041 9263 8075
rect 10057 8041 10091 8075
rect 12081 8041 12115 8075
rect 14657 8041 14691 8075
rect 15117 8041 15151 8075
rect 16405 8041 16439 8075
rect 1685 7973 1719 8007
rect 2599 7973 2633 8007
rect 7475 7973 7509 8007
rect 11523 7973 11557 8007
rect 13553 7973 13587 8007
rect 13829 7973 13863 8007
rect 15485 7973 15519 8007
rect 17206 7973 17240 8007
rect 18889 7973 18923 8007
rect 2237 7905 2271 7939
rect 3157 7905 3191 7939
rect 4813 7905 4847 7939
rect 9781 7905 9815 7939
rect 9965 7905 9999 7939
rect 10701 7905 10735 7939
rect 16957 7905 16991 7939
rect 17877 7905 17911 7939
rect 3801 7837 3835 7871
rect 7113 7837 7147 7871
rect 11161 7837 11195 7871
rect 13185 7837 13219 7871
rect 13737 7837 13771 7871
rect 15393 7837 15427 7871
rect 15669 7837 15703 7871
rect 18797 7837 18831 7871
rect 19073 7837 19107 7871
rect 6009 7769 6043 7803
rect 14289 7769 14323 7803
rect 5733 7701 5767 7735
rect 6377 7701 6411 7735
rect 6929 7701 6963 7735
rect 8033 7701 8067 7735
rect 8585 7701 8619 7735
rect 11069 7701 11103 7735
rect 12357 7701 12391 7735
rect 18521 7701 18555 7735
rect 2329 7497 2363 7531
rect 2697 7497 2731 7531
rect 6193 7497 6227 7531
rect 12449 7497 12483 7531
rect 12817 7497 12851 7531
rect 14841 7497 14875 7531
rect 15393 7497 15427 7531
rect 15669 7497 15703 7531
rect 16221 7497 16255 7531
rect 17693 7497 17727 7531
rect 18429 7497 18463 7531
rect 19533 7497 19567 7531
rect 5825 7429 5859 7463
rect 11529 7429 11563 7463
rect 1409 7361 1443 7395
rect 3893 7361 3927 7395
rect 5273 7361 5307 7395
rect 7205 7361 7239 7395
rect 10609 7361 10643 7395
rect 19901 7429 19935 7463
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 8493 7293 8527 7327
rect 12449 7293 12483 7327
rect 12725 7293 12759 7327
rect 13369 7293 13403 7327
rect 13921 7293 13955 7327
rect 16497 7293 16531 7327
rect 16773 7293 16807 7327
rect 3249 7225 3283 7259
rect 3341 7225 3375 7259
rect 4537 7225 4571 7259
rect 5365 7225 5399 7259
rect 6929 7225 6963 7259
rect 7021 7225 7055 7259
rect 7941 7225 7975 7259
rect 8401 7225 8435 7259
rect 8855 7225 8889 7259
rect 10517 7225 10551 7259
rect 10971 7225 11005 7259
rect 12541 7225 12575 7259
rect 17049 7225 17083 7259
rect 18705 7225 18739 7259
rect 1777 7157 1811 7191
rect 3065 7157 3099 7191
rect 4905 7157 4939 7191
rect 6561 7157 6595 7191
rect 9413 7157 9447 7191
rect 9781 7157 9815 7191
rect 11897 7157 11931 7191
rect 12265 7157 12299 7191
rect 13737 7157 13771 7191
rect 14289 7157 14323 7191
rect 17325 7157 17359 7191
rect 1547 6953 1581 6987
rect 6745 6953 6779 6987
rect 9045 6953 9079 6987
rect 11069 6953 11103 6987
rect 13921 6953 13955 6987
rect 14381 6953 14415 6987
rect 17877 6953 17911 6987
rect 18613 6953 18647 6987
rect 1961 6885 1995 6919
rect 2237 6885 2271 6919
rect 2605 6885 2639 6919
rect 4721 6885 4755 6919
rect 5549 6885 5583 6919
rect 7113 6885 7147 6919
rect 12909 6885 12943 6919
rect 17319 6885 17353 6919
rect 18889 6885 18923 6919
rect 1476 6817 1510 6851
rect 3157 6817 3191 6851
rect 4077 6817 4111 6851
rect 6101 6817 6135 6851
rect 8493 6817 8527 6851
rect 9873 6817 9907 6851
rect 10977 6817 11011 6851
rect 11805 6817 11839 6851
rect 13461 6817 13495 6851
rect 15393 6817 15427 6851
rect 15945 6817 15979 6851
rect 2513 6749 2547 6783
rect 5457 6749 5491 6783
rect 7021 6749 7055 6783
rect 7297 6749 7331 6783
rect 10517 6749 10551 6783
rect 11713 6749 11747 6783
rect 16129 6749 16163 6783
rect 16957 6749 16991 6783
rect 18797 6749 18831 6783
rect 19073 6749 19107 6783
rect 7941 6681 7975 6715
rect 8677 6681 8711 6715
rect 16405 6681 16439 6715
rect 3433 6613 3467 6647
rect 3801 6613 3835 6647
rect 4261 6613 4295 6647
rect 4997 6613 5031 6647
rect 6377 6613 6411 6647
rect 10057 6613 10091 6647
rect 10793 6613 10827 6647
rect 12541 6613 12575 6647
rect 14841 6613 14875 6647
rect 16773 6613 16807 6647
rect 1547 6409 1581 6443
rect 3341 6409 3375 6443
rect 5457 6409 5491 6443
rect 5825 6409 5859 6443
rect 6653 6409 6687 6443
rect 8585 6409 8619 6443
rect 9873 6409 9907 6443
rect 13461 6409 13495 6443
rect 16221 6409 16255 6443
rect 17785 6409 17819 6443
rect 18521 6409 18555 6443
rect 6193 6341 6227 6375
rect 7941 6341 7975 6375
rect 11161 6341 11195 6375
rect 13829 6341 13863 6375
rect 15945 6341 15979 6375
rect 2329 6273 2363 6307
rect 4537 6273 4571 6307
rect 7389 6273 7423 6307
rect 8953 6273 8987 6307
rect 9229 6273 9263 6307
rect 14749 6273 14783 6307
rect 17141 6273 17175 6307
rect 18705 6273 18739 6307
rect 19993 6273 20027 6307
rect 1476 6205 1510 6239
rect 2421 6205 2455 6239
rect 3709 6205 3743 6239
rect 10425 6205 10459 6239
rect 11253 6205 11287 6239
rect 11437 6205 11471 6239
rect 12541 6205 12575 6239
rect 13001 6205 13035 6239
rect 14841 6205 14875 6239
rect 15393 6205 15427 6239
rect 4899 6137 4933 6171
rect 7481 6137 7515 6171
rect 9045 6137 9079 6171
rect 10241 6137 10275 6171
rect 15577 6137 15611 6171
rect 16497 6137 16531 6171
rect 16598 6137 16632 6171
rect 18797 6137 18831 6171
rect 19349 6137 19383 6171
rect 1869 6069 1903 6103
rect 2789 6069 2823 6103
rect 4169 6069 4203 6103
rect 7205 6069 7239 6103
rect 11805 6069 11839 6103
rect 12265 6069 12299 6103
rect 12541 6069 12575 6103
rect 17417 6069 17451 6103
rect 19625 6069 19659 6103
rect 3433 5865 3467 5899
rect 3893 5865 3927 5899
rect 5181 5865 5215 5899
rect 6101 5865 6135 5899
rect 6561 5865 6595 5899
rect 8493 5865 8527 5899
rect 9045 5865 9079 5899
rect 9781 5865 9815 5899
rect 10977 5865 11011 5899
rect 11437 5865 11471 5899
rect 12817 5865 12851 5899
rect 13553 5865 13587 5899
rect 15025 5865 15059 5899
rect 15945 5865 15979 5899
rect 16865 5865 16899 5899
rect 17969 5865 18003 5899
rect 18245 5865 18279 5899
rect 2973 5797 3007 5831
rect 4813 5797 4847 5831
rect 6745 5797 6779 5831
rect 6837 5797 6871 5831
rect 13093 5797 13127 5831
rect 15301 5797 15335 5831
rect 16497 5797 16531 5831
rect 17411 5797 17445 5831
rect 18981 5797 19015 5831
rect 2237 5729 2271 5763
rect 2789 5729 2823 5763
rect 4077 5729 4111 5763
rect 4537 5729 4571 5763
rect 5708 5729 5742 5763
rect 8217 5729 8251 5763
rect 8401 5729 8435 5763
rect 9689 5729 9723 5763
rect 10149 5729 10183 5763
rect 11345 5729 11379 5763
rect 12173 5729 12207 5763
rect 13277 5729 13311 5763
rect 14105 5729 14139 5763
rect 17049 5729 17083 5763
rect 8033 5661 8067 5695
rect 12265 5661 12299 5695
rect 14013 5661 14047 5695
rect 15669 5661 15703 5695
rect 18889 5661 18923 5695
rect 19349 5661 19383 5695
rect 5457 5593 5491 5627
rect 7297 5593 7331 5627
rect 15577 5593 15611 5627
rect 1961 5525 1995 5559
rect 5779 5525 5813 5559
rect 7665 5525 7699 5559
rect 9413 5525 9447 5559
rect 14657 5525 14691 5559
rect 15466 5525 15500 5559
rect 18705 5525 18739 5559
rect 2973 5321 3007 5355
rect 4537 5321 4571 5355
rect 4905 5321 4939 5355
rect 10057 5321 10091 5355
rect 10701 5321 10735 5355
rect 12173 5321 12207 5355
rect 12587 5321 12621 5355
rect 14473 5321 14507 5355
rect 15117 5321 15151 5355
rect 16865 5321 16899 5355
rect 18981 5321 19015 5355
rect 6653 5253 6687 5287
rect 9045 5253 9079 5287
rect 11437 5253 11471 5287
rect 16037 5253 16071 5287
rect 19625 5253 19659 5287
rect 2605 5185 2639 5219
rect 4997 5185 5031 5219
rect 6929 5185 6963 5219
rect 7297 5185 7331 5219
rect 7849 5185 7883 5219
rect 8493 5185 8527 5219
rect 10885 5185 10919 5219
rect 13277 5185 13311 5219
rect 13553 5185 13587 5219
rect 18061 5185 18095 5219
rect 1869 5117 1903 5151
rect 1961 5117 1995 5151
rect 2145 5117 2179 5151
rect 3341 5117 3375 5151
rect 3433 5117 3467 5151
rect 3525 5117 3559 5151
rect 3709 5117 3743 5151
rect 6285 5117 6319 5151
rect 8217 5117 8251 5151
rect 12516 5117 12550 5151
rect 15025 5117 15059 5151
rect 15761 5117 15795 5151
rect 16773 5117 16807 5151
rect 17509 5117 17543 5151
rect 1777 5049 1811 5083
rect 5318 5049 5352 5083
rect 7021 5049 7055 5083
rect 8585 5049 8619 5083
rect 9689 5049 9723 5083
rect 10977 5049 11011 5083
rect 13645 5049 13679 5083
rect 14197 5049 14231 5083
rect 16405 5049 16439 5083
rect 16589 5049 16623 5083
rect 3893 4981 3927 5015
rect 5917 4981 5951 5015
rect 11805 4981 11839 5015
rect 13001 4981 13035 5015
rect 14841 4981 14875 5015
rect 17877 4981 17911 5015
rect 18429 4981 18463 5015
rect 19257 4981 19291 5015
rect 1547 4777 1581 4811
rect 1869 4777 1903 4811
rect 3801 4777 3835 4811
rect 5089 4777 5123 4811
rect 5457 4777 5491 4811
rect 6561 4777 6595 4811
rect 7205 4777 7239 4811
rect 8493 4777 8527 4811
rect 10885 4777 10919 4811
rect 12081 4777 12115 4811
rect 15117 4777 15151 4811
rect 15945 4777 15979 4811
rect 16589 4777 16623 4811
rect 18337 4777 18371 4811
rect 2421 4709 2455 4743
rect 3157 4709 3191 4743
rect 4813 4709 4847 4743
rect 6003 4709 6037 4743
rect 7573 4709 7607 4743
rect 8125 4709 8159 4743
rect 9689 4709 9723 4743
rect 11253 4709 11287 4743
rect 11805 4709 11839 4743
rect 12995 4709 13029 4743
rect 17779 4709 17813 4743
rect 19165 4709 19199 4743
rect 1476 4641 1510 4675
rect 2568 4641 2602 4675
rect 3525 4641 3559 4675
rect 4077 4641 4111 4675
rect 4169 4641 4203 4675
rect 4353 4641 4387 4675
rect 5641 4641 5675 4675
rect 6837 4641 6871 4675
rect 9873 4641 9907 4675
rect 12633 4641 12667 4675
rect 13921 4641 13955 4675
rect 15301 4641 15335 4675
rect 19349 4641 19383 4675
rect 2789 4573 2823 4607
rect 7481 4573 7515 4607
rect 11161 4573 11195 4607
rect 12541 4573 12575 4607
rect 14749 4573 14783 4607
rect 15669 4573 15703 4607
rect 17417 4573 17451 4607
rect 2329 4505 2363 4539
rect 14197 4505 14231 4539
rect 15577 4505 15611 4539
rect 2697 4437 2731 4471
rect 8769 4437 8803 4471
rect 9229 4437 9263 4471
rect 9965 4437 9999 4471
rect 13553 4437 13587 4471
rect 15466 4437 15500 4471
rect 17049 4437 17083 4471
rect 19441 4437 19475 4471
rect 2973 4233 3007 4267
rect 4629 4233 4663 4267
rect 6561 4233 6595 4267
rect 7021 4233 7055 4267
rect 9045 4233 9079 4267
rect 9505 4233 9539 4267
rect 12173 4233 12207 4267
rect 13461 4233 13495 4267
rect 15577 4233 15611 4267
rect 19165 4233 19199 4267
rect 19763 4233 19797 4267
rect 20085 4233 20119 4267
rect 1685 4097 1719 4131
rect 3157 4165 3191 4199
rect 5089 4165 5123 4199
rect 7757 4165 7791 4199
rect 10241 4165 10275 4199
rect 11069 4165 11103 4199
rect 3801 4097 3835 4131
rect 4353 4097 4387 4131
rect 5917 4097 5951 4131
rect 7481 4097 7515 4131
rect 9689 4097 9723 4131
rect 10609 4097 10643 4131
rect 12541 4097 12575 4131
rect 13921 4097 13955 4131
rect 14381 4097 14415 4131
rect 17877 4097 17911 4131
rect 2329 4029 2363 4063
rect 2789 4029 2823 4063
rect 2973 4029 3007 4063
rect 3249 4029 3283 4063
rect 3341 4029 3375 4063
rect 3525 4029 3559 4063
rect 5457 4029 5491 4063
rect 5641 4029 5675 4063
rect 6837 4029 6871 4063
rect 11161 4029 11195 4063
rect 11713 4029 11747 4063
rect 16221 4029 16255 4063
rect 16773 4029 16807 4063
rect 18245 4029 18279 4063
rect 18521 4029 18555 4063
rect 19692 4029 19726 4063
rect 8033 3961 8067 3995
rect 8125 3961 8159 3995
rect 8677 3961 8711 3995
rect 9781 3961 9815 3995
rect 12633 3961 12667 3995
rect 13185 3961 13219 3995
rect 16957 3961 16991 3995
rect 18797 3961 18831 3995
rect 20453 3961 20487 3995
rect 6285 3893 6319 3927
rect 11345 3893 11379 3927
rect 14197 3893 14231 3927
rect 14749 3893 14783 3927
rect 15301 3893 15335 3927
rect 16037 3893 16071 3927
rect 17417 3893 17451 3927
rect 1409 3689 1443 3723
rect 5549 3689 5583 3723
rect 5917 3689 5951 3723
rect 8585 3689 8619 3723
rect 9229 3689 9263 3723
rect 10241 3689 10275 3723
rect 11805 3689 11839 3723
rect 12633 3689 12667 3723
rect 13001 3689 13035 3723
rect 15025 3689 15059 3723
rect 16405 3689 16439 3723
rect 18245 3689 18279 3723
rect 18705 3689 18739 3723
rect 2329 3621 2363 3655
rect 3157 3621 3191 3655
rect 6193 3621 6227 3655
rect 6285 3621 6319 3655
rect 7986 3621 8020 3655
rect 11247 3621 11281 3655
rect 13553 3621 13587 3655
rect 14105 3621 14139 3655
rect 14749 3621 14783 3655
rect 15393 3621 15427 3655
rect 15485 3621 15519 3655
rect 16037 3621 16071 3655
rect 17298 3621 17332 3655
rect 18981 3621 19015 3655
rect 1961 3553 1995 3587
rect 2421 3553 2455 3587
rect 2697 3553 2731 3587
rect 3893 3553 3927 3587
rect 4261 3553 4295 3587
rect 4813 3553 4847 3587
rect 5089 3553 5123 3587
rect 6837 3553 6871 3587
rect 9689 3553 9723 3587
rect 12081 3553 12115 3587
rect 16681 3553 16715 3587
rect 17969 3553 18003 3587
rect 5273 3485 5307 3519
rect 7665 3485 7699 3519
rect 10885 3485 10919 3519
rect 13461 3485 13495 3519
rect 17049 3485 17083 3519
rect 18889 3485 18923 3519
rect 19165 3485 19199 3519
rect 2513 3417 2547 3451
rect 3433 3349 3467 3383
rect 7389 3349 7423 3383
rect 9873 3349 9907 3383
rect 10701 3349 10735 3383
rect 2421 3145 2455 3179
rect 2697 3145 2731 3179
rect 2881 3145 2915 3179
rect 4537 3145 4571 3179
rect 6193 3145 6227 3179
rect 10057 3145 10091 3179
rect 10425 3145 10459 3179
rect 10977 3145 11011 3179
rect 12081 3145 12115 3179
rect 12173 3145 12207 3179
rect 13553 3145 13587 3179
rect 15117 3145 15151 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 19441 3145 19475 3179
rect 2145 3009 2179 3043
rect 3065 3077 3099 3111
rect 3985 3077 4019 3111
rect 11437 3077 11471 3111
rect 4997 3009 5031 3043
rect 7389 3009 7423 3043
rect 8033 3009 8067 3043
rect 9137 3009 9171 3043
rect 1685 2941 1719 2975
rect 1961 2941 1995 2975
rect 2697 2941 2731 2975
rect 2973 2941 3007 2975
rect 3249 2941 3283 2975
rect 3709 2941 3743 2975
rect 4905 2941 4939 2975
rect 11253 2941 11287 2975
rect 11805 2941 11839 2975
rect 19073 3077 19107 3111
rect 12541 3009 12575 3043
rect 13185 3009 13219 3043
rect 14105 3009 14139 3043
rect 14749 3009 14783 3043
rect 19763 3009 19797 3043
rect 15577 2941 15611 2975
rect 18061 2941 18095 2975
rect 18521 2941 18555 2975
rect 19676 2941 19710 2975
rect 20085 2941 20119 2975
rect 5318 2873 5352 2907
rect 6561 2873 6595 2907
rect 7021 2873 7055 2907
rect 7481 2873 7515 2907
rect 8401 2873 8435 2907
rect 9045 2873 9079 2907
rect 9499 2873 9533 2907
rect 12081 2873 12115 2907
rect 12633 2873 12667 2907
rect 14197 2873 14231 2907
rect 15393 2873 15427 2907
rect 15898 2873 15932 2907
rect 17049 2873 17083 2907
rect 5917 2805 5951 2839
rect 13921 2805 13955 2839
rect 16497 2805 16531 2839
rect 18153 2805 18187 2839
rect 2329 2601 2363 2635
rect 3801 2601 3835 2635
rect 4261 2601 4295 2635
rect 5089 2601 5123 2635
rect 6101 2601 6135 2635
rect 6377 2601 6411 2635
rect 6745 2601 6779 2635
rect 7849 2601 7883 2635
rect 8815 2601 8849 2635
rect 9919 2601 9953 2635
rect 10701 2601 10735 2635
rect 11713 2601 11747 2635
rect 12357 2601 12391 2635
rect 13093 2601 13127 2635
rect 13461 2601 13495 2635
rect 14565 2601 14599 2635
rect 14841 2601 14875 2635
rect 15301 2601 15335 2635
rect 16129 2601 16163 2635
rect 17325 2601 17359 2635
rect 18061 2601 18095 2635
rect 1685 2533 1719 2567
rect 5457 2533 5491 2567
rect 6009 2533 6043 2567
rect 1476 2465 1510 2499
rect 2421 2465 2455 2499
rect 2697 2465 2731 2499
rect 3157 2465 3191 2499
rect 4102 2465 4136 2499
rect 4629 2397 4663 2431
rect 5365 2397 5399 2431
rect 7291 2533 7325 2567
rect 8125 2533 8159 2567
rect 11114 2533 11148 2567
rect 13966 2533 14000 2567
rect 15853 2533 15887 2567
rect 16497 2533 16531 2567
rect 17693 2533 17727 2567
rect 6929 2465 6963 2499
rect 8493 2465 8527 2499
rect 8744 2465 8778 2499
rect 9137 2465 9171 2499
rect 9848 2465 9882 2499
rect 10241 2465 10275 2499
rect 12700 2465 12734 2499
rect 16037 2465 16071 2499
rect 18337 2465 18371 2499
rect 18797 2465 18831 2499
rect 10793 2397 10827 2431
rect 13645 2397 13679 2431
rect 2513 2329 2547 2363
rect 6101 2329 6135 2363
rect 9505 2329 9539 2363
rect 12081 2329 12115 2363
rect 16405 2397 16439 2431
rect 18889 2397 18923 2431
rect 16957 2329 16991 2363
rect 1961 2261 1995 2295
rect 3525 2261 3559 2295
rect 12771 2261 12805 2295
rect 16037 2261 16071 2295
rect 19349 2261 19383 2295
<< metal1 >>
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17310 21536 17316 21548
rect 16632 21508 17316 21536
rect 16632 21496 16638 21508
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 1104 19610 20884 19632
rect 1104 19558 4648 19610
rect 4700 19558 4712 19610
rect 4764 19558 4776 19610
rect 4828 19558 4840 19610
rect 4892 19558 11982 19610
rect 12034 19558 12046 19610
rect 12098 19558 12110 19610
rect 12162 19558 12174 19610
rect 12226 19558 19315 19610
rect 19367 19558 19379 19610
rect 19431 19558 19443 19610
rect 19495 19558 19507 19610
rect 19559 19558 20884 19610
rect 1104 19536 20884 19558
rect 10275 19431 10333 19437
rect 10275 19397 10287 19431
rect 10321 19428 10333 19431
rect 11054 19428 11060 19440
rect 10321 19400 11060 19428
rect 10321 19397 10333 19400
rect 10275 19391 10333 19397
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 10204 19295 10262 19301
rect 10204 19261 10216 19295
rect 10250 19292 10262 19295
rect 11216 19295 11274 19301
rect 10250 19264 10732 19292
rect 10250 19261 10262 19264
rect 10204 19255 10262 19261
rect 10704 19168 10732 19264
rect 11216 19261 11228 19295
rect 11262 19292 11274 19295
rect 13148 19295 13206 19301
rect 11262 19264 11652 19292
rect 11262 19261 11274 19264
rect 11216 19255 11274 19261
rect 11624 19168 11652 19264
rect 13148 19261 13160 19295
rect 13194 19292 13206 19295
rect 14144 19295 14202 19301
rect 13194 19264 13400 19292
rect 13194 19261 13206 19264
rect 13148 19255 13206 19261
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11287 19159 11345 19165
rect 11287 19156 11299 19159
rect 11020 19128 11299 19156
rect 11020 19116 11026 19128
rect 11287 19125 11299 19128
rect 11333 19125 11345 19159
rect 11606 19156 11612 19168
rect 11567 19128 11612 19156
rect 11287 19119 11345 19125
rect 11606 19116 11612 19128
rect 11664 19116 11670 19168
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 13219 19159 13277 19165
rect 13219 19156 13231 19159
rect 12676 19128 13231 19156
rect 12676 19116 12682 19128
rect 13219 19125 13231 19128
rect 13265 19125 13277 19159
rect 13372 19156 13400 19264
rect 14144 19261 14156 19295
rect 14190 19292 14202 19295
rect 14190 19264 14688 19292
rect 14190 19261 14202 19264
rect 14144 19255 14202 19261
rect 14660 19168 14688 19264
rect 13538 19156 13544 19168
rect 13372 19128 13544 19156
rect 13219 19119 13277 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14231 19159 14289 19165
rect 14231 19156 14243 19159
rect 13872 19128 14243 19156
rect 13872 19116 13878 19128
rect 14231 19125 14243 19128
rect 14277 19125 14289 19159
rect 14642 19156 14648 19168
rect 14603 19128 14648 19156
rect 14231 19119 14289 19125
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 1104 19066 20884 19088
rect 1104 19014 8315 19066
rect 8367 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 15648 19066
rect 15700 19014 15712 19066
rect 15764 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 20884 19066
rect 1104 18992 20884 19014
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 19150 18952 19156 18964
rect 10744 18924 19156 18952
rect 10744 18912 10750 18924
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 6546 18844 6552 18896
rect 6604 18884 6610 18896
rect 10502 18884 10508 18896
rect 6604 18856 10508 18884
rect 6604 18844 6610 18856
rect 10502 18844 10508 18856
rect 10560 18884 10566 18896
rect 10560 18856 11652 18884
rect 10560 18844 10566 18856
rect 8202 18776 8208 18828
rect 8260 18816 8266 18828
rect 10686 18825 10692 18828
rect 8608 18819 8666 18825
rect 8608 18816 8620 18819
rect 8260 18788 8620 18816
rect 8260 18776 8266 18788
rect 8608 18785 8620 18788
rect 8654 18785 8666 18819
rect 10664 18819 10692 18825
rect 10664 18816 10676 18819
rect 10599 18788 10676 18816
rect 8608 18779 8666 18785
rect 10664 18785 10676 18788
rect 10744 18816 10750 18828
rect 11514 18816 11520 18828
rect 10744 18788 11520 18816
rect 10664 18779 10692 18785
rect 10686 18776 10692 18779
rect 10744 18776 10750 18788
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 11624 18825 11652 18856
rect 11624 18819 11702 18825
rect 11624 18788 11656 18819
rect 11644 18785 11656 18788
rect 11690 18816 11702 18819
rect 11790 18816 11796 18828
rect 11690 18788 11796 18816
rect 11690 18785 11702 18788
rect 11644 18779 11702 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 13484 18819 13542 18825
rect 13484 18816 13496 18819
rect 13412 18788 13496 18816
rect 13412 18776 13418 18788
rect 13484 18785 13496 18788
rect 13530 18785 13542 18819
rect 13484 18779 13542 18785
rect 15356 18819 15414 18825
rect 15356 18785 15368 18819
rect 15402 18816 15414 18819
rect 16022 18816 16028 18828
rect 15402 18788 16028 18816
rect 15402 18785 15414 18788
rect 15356 18779 15414 18785
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 8711 18615 8769 18621
rect 8711 18581 8723 18615
rect 8757 18612 8769 18615
rect 8846 18612 8852 18624
rect 8757 18584 8852 18612
rect 8757 18581 8769 18584
rect 8711 18575 8769 18581
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 10735 18615 10793 18621
rect 10735 18581 10747 18615
rect 10781 18612 10793 18615
rect 10870 18612 10876 18624
rect 10781 18584 10876 18612
rect 10781 18581 10793 18584
rect 10735 18575 10793 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11514 18572 11520 18624
rect 11572 18612 11578 18624
rect 11747 18615 11805 18621
rect 11747 18612 11759 18615
rect 11572 18584 11759 18612
rect 11572 18572 11578 18584
rect 11747 18581 11759 18584
rect 11793 18581 11805 18615
rect 11747 18575 11805 18581
rect 13587 18615 13645 18621
rect 13587 18581 13599 18615
rect 13633 18612 13645 18615
rect 13722 18612 13728 18624
rect 13633 18584 13728 18612
rect 13633 18581 13645 18584
rect 13587 18575 13645 18581
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 14826 18572 14832 18624
rect 14884 18612 14890 18624
rect 15427 18615 15485 18621
rect 15427 18612 15439 18615
rect 14884 18584 15439 18612
rect 14884 18572 14890 18584
rect 15427 18581 15439 18584
rect 15473 18581 15485 18615
rect 15427 18575 15485 18581
rect 1104 18522 20884 18544
rect 1104 18470 4648 18522
rect 4700 18470 4712 18522
rect 4764 18470 4776 18522
rect 4828 18470 4840 18522
rect 4892 18470 11982 18522
rect 12034 18470 12046 18522
rect 12098 18470 12110 18522
rect 12162 18470 12174 18522
rect 12226 18470 19315 18522
rect 19367 18470 19379 18522
rect 19431 18470 19443 18522
rect 19495 18470 19507 18522
rect 19559 18470 20884 18522
rect 1104 18448 20884 18470
rect 7469 18411 7527 18417
rect 7469 18377 7481 18411
rect 7515 18408 7527 18411
rect 7742 18408 7748 18420
rect 7515 18380 7748 18408
rect 7515 18377 7527 18380
rect 7469 18371 7527 18377
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 10686 18408 10692 18420
rect 10647 18380 10692 18408
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 11790 18368 11796 18420
rect 11848 18408 11854 18420
rect 11977 18411 12035 18417
rect 11977 18408 11989 18411
rect 11848 18380 11989 18408
rect 11848 18368 11854 18380
rect 11977 18377 11989 18380
rect 12023 18377 12035 18411
rect 11977 18371 12035 18377
rect 14461 18411 14519 18417
rect 14461 18377 14473 18411
rect 14507 18408 14519 18411
rect 14737 18411 14795 18417
rect 14737 18408 14749 18411
rect 14507 18380 14749 18408
rect 14507 18377 14519 18380
rect 14461 18371 14519 18377
rect 14737 18377 14749 18380
rect 14783 18408 14795 18411
rect 15194 18408 15200 18420
rect 14783 18380 15200 18408
rect 14783 18377 14795 18380
rect 14737 18371 14795 18377
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 8987 18343 9045 18349
rect 8987 18340 8999 18343
rect 7432 18312 8999 18340
rect 7432 18300 7438 18312
rect 8987 18309 8999 18312
rect 9033 18309 9045 18343
rect 8987 18303 9045 18309
rect 4430 18232 4436 18284
rect 4488 18272 4494 18284
rect 11992 18272 12020 18371
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 12161 18343 12219 18349
rect 12161 18309 12173 18343
rect 12207 18340 12219 18343
rect 14366 18340 14372 18352
rect 12207 18312 14372 18340
rect 12207 18309 12219 18312
rect 12161 18303 12219 18309
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 14550 18300 14556 18352
rect 14608 18340 14614 18352
rect 15335 18343 15393 18349
rect 15335 18340 15347 18343
rect 14608 18312 15347 18340
rect 14608 18300 14614 18312
rect 15335 18309 15347 18312
rect 15381 18309 15393 18343
rect 15335 18303 15393 18309
rect 4488 18244 10215 18272
rect 4488 18232 4494 18244
rect 10187 18213 10215 18244
rect 10980 18244 11928 18272
rect 11992 18244 15056 18272
rect 10980 18213 11008 18244
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18204 7343 18207
rect 8916 18207 8974 18213
rect 7331 18176 7972 18204
rect 7331 18173 7343 18176
rect 7285 18167 7343 18173
rect 7944 18145 7972 18176
rect 8916 18173 8928 18207
rect 8962 18204 8974 18207
rect 10172 18207 10230 18213
rect 8962 18176 9444 18204
rect 8962 18173 8974 18176
rect 8916 18167 8974 18173
rect 7929 18139 7987 18145
rect 7929 18105 7941 18139
rect 7975 18136 7987 18139
rect 8754 18136 8760 18148
rect 7975 18108 8760 18136
rect 7975 18105 7987 18108
rect 7929 18099 7987 18105
rect 8754 18096 8760 18108
rect 8812 18096 8818 18148
rect 9416 18080 9444 18176
rect 10172 18173 10184 18207
rect 10218 18204 10230 18207
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10218 18176 10977 18204
rect 10218 18173 10230 18176
rect 10172 18167 10230 18173
rect 10965 18173 10977 18176
rect 11011 18173 11023 18207
rect 11146 18204 11152 18216
rect 11110 18176 11152 18204
rect 10965 18167 11023 18173
rect 11146 18164 11152 18176
rect 11204 18213 11210 18216
rect 11204 18207 11258 18213
rect 11204 18173 11212 18207
rect 11246 18204 11258 18207
rect 11606 18204 11612 18216
rect 11246 18176 11612 18204
rect 11246 18173 11258 18176
rect 11204 18167 11258 18173
rect 11204 18164 11210 18167
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 11900 18204 11928 18244
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 11900 18176 12173 18204
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 12161 18167 12219 18173
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 13538 18204 13544 18216
rect 13320 18176 13544 18204
rect 13320 18164 13326 18176
rect 13538 18164 13544 18176
rect 13596 18204 13602 18216
rect 14236 18207 14294 18213
rect 14236 18204 14248 18207
rect 13596 18176 14248 18204
rect 13596 18164 13602 18176
rect 14236 18173 14248 18176
rect 14282 18204 14294 18207
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 14282 18176 14473 18204
rect 14282 18173 14294 18176
rect 14236 18167 14294 18173
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 15028 18204 15056 18244
rect 15232 18207 15290 18213
rect 15232 18204 15244 18207
rect 15028 18176 15244 18204
rect 14461 18167 14519 18173
rect 15232 18173 15244 18176
rect 15278 18204 15290 18207
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15278 18176 15669 18204
rect 15278 18173 15290 18176
rect 15232 18167 15290 18173
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 18116 18207 18174 18213
rect 18116 18173 18128 18207
rect 18162 18173 18174 18207
rect 18116 18167 18174 18173
rect 10275 18139 10333 18145
rect 10275 18105 10287 18139
rect 10321 18136 10333 18139
rect 10686 18136 10692 18148
rect 10321 18108 10692 18136
rect 10321 18105 10333 18108
rect 10275 18099 10333 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 11287 18139 11345 18145
rect 11287 18105 11299 18139
rect 11333 18136 11345 18139
rect 11882 18136 11888 18148
rect 11333 18108 11888 18136
rect 11333 18105 11345 18108
rect 11287 18099 11345 18105
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 14323 18139 14381 18145
rect 14323 18105 14335 18139
rect 14369 18136 14381 18139
rect 14734 18136 14740 18148
rect 14369 18108 14740 18136
rect 14369 18105 14381 18108
rect 14323 18099 14381 18105
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 18131 18136 18159 18167
rect 18506 18136 18512 18148
rect 18131 18108 18512 18136
rect 18506 18096 18512 18108
rect 18564 18096 18570 18148
rect 8202 18028 8208 18080
rect 8260 18068 8266 18080
rect 8573 18071 8631 18077
rect 8573 18068 8585 18071
rect 8260 18040 8585 18068
rect 8260 18028 8266 18040
rect 8573 18037 8585 18040
rect 8619 18037 8631 18071
rect 9398 18068 9404 18080
rect 9359 18040 9404 18068
rect 8573 18031 8631 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 12434 18068 12440 18080
rect 12395 18040 12440 18068
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 13354 18068 13360 18080
rect 12860 18040 13360 18068
rect 12860 18028 12866 18040
rect 13354 18028 13360 18040
rect 13412 18068 13418 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 13412 18040 13461 18068
rect 13412 18028 13418 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 16022 18068 16028 18080
rect 15983 18040 16028 18068
rect 13449 18031 13507 18037
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 18187 18071 18245 18077
rect 18187 18068 18199 18071
rect 16448 18040 18199 18068
rect 16448 18028 16454 18040
rect 18187 18037 18199 18040
rect 18233 18037 18245 18071
rect 18187 18031 18245 18037
rect 1104 17978 20884 18000
rect 1104 17926 8315 17978
rect 8367 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 15648 17978
rect 15700 17926 15712 17978
rect 15764 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 20884 17978
rect 1104 17904 20884 17926
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 13136 17836 13185 17864
rect 13136 17824 13142 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 16758 17796 16764 17808
rect 9456 17768 16764 17796
rect 9456 17756 9462 17768
rect 16758 17756 16764 17768
rect 16816 17756 16822 17808
rect 6273 17731 6331 17737
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 6362 17728 6368 17740
rect 6319 17700 6368 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 7628 17731 7686 17737
rect 7628 17697 7640 17731
rect 7674 17728 7686 17731
rect 7742 17728 7748 17740
rect 7674 17700 7748 17728
rect 7674 17697 7686 17700
rect 7628 17691 7686 17697
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 8662 17728 8668 17740
rect 8619 17700 8668 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 8662 17688 8668 17700
rect 8720 17688 8726 17740
rect 11492 17731 11550 17737
rect 11492 17697 11504 17731
rect 11538 17728 11550 17731
rect 11698 17728 11704 17740
rect 11538 17700 11704 17728
rect 11538 17697 11550 17700
rect 11492 17691 11550 17697
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17697 13415 17731
rect 13538 17728 13544 17740
rect 13499 17700 13544 17728
rect 13357 17691 13415 17697
rect 9674 17660 9680 17672
rect 9635 17632 9680 17660
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 13372 17660 13400 17691
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 16298 17728 16304 17740
rect 16259 17700 16304 17728
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 17402 17688 17408 17740
rect 17460 17728 17466 17740
rect 17624 17731 17682 17737
rect 17624 17728 17636 17731
rect 17460 17700 17636 17728
rect 17460 17688 17466 17700
rect 17624 17697 17636 17700
rect 17670 17697 17682 17731
rect 17624 17691 17682 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17728 18659 17731
rect 18690 17728 18696 17740
rect 18647 17700 18696 17728
rect 18647 17697 18659 17700
rect 18601 17691 18659 17697
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 19150 17688 19156 17740
rect 19208 17728 19214 17740
rect 19702 17737 19708 17740
rect 19648 17731 19708 17737
rect 19648 17728 19660 17731
rect 19208 17700 19660 17728
rect 19208 17688 19214 17700
rect 19648 17697 19660 17700
rect 19694 17697 19708 17731
rect 19648 17691 19708 17697
rect 19702 17688 19708 17691
rect 19760 17688 19766 17740
rect 13446 17660 13452 17672
rect 13372 17632 13452 17660
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 15378 17660 15384 17672
rect 15335 17632 15384 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 17218 17552 17224 17604
rect 17276 17592 17282 17604
rect 19751 17595 19809 17601
rect 19751 17592 19763 17595
rect 17276 17564 19763 17592
rect 17276 17552 17282 17564
rect 19751 17561 19763 17564
rect 19797 17561 19809 17595
rect 19751 17555 19809 17561
rect 6411 17527 6469 17533
rect 6411 17493 6423 17527
rect 6457 17524 6469 17527
rect 6546 17524 6552 17536
rect 6457 17496 6552 17524
rect 6457 17493 6469 17496
rect 6411 17487 6469 17493
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 7699 17527 7757 17533
rect 7699 17524 7711 17527
rect 7616 17496 7711 17524
rect 7616 17484 7622 17496
rect 7699 17493 7711 17496
rect 7745 17493 7757 17527
rect 7699 17487 7757 17493
rect 8711 17527 8769 17533
rect 8711 17493 8723 17527
rect 8757 17524 8769 17527
rect 9122 17524 9128 17536
rect 8757 17496 9128 17524
rect 8757 17493 8769 17496
rect 8711 17487 8769 17493
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 11563 17527 11621 17533
rect 11563 17493 11575 17527
rect 11609 17524 11621 17527
rect 11790 17524 11796 17536
rect 11609 17496 11796 17524
rect 11609 17493 11621 17496
rect 11563 17487 11621 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12768 17496 12817 17524
rect 12768 17484 12774 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 14090 17524 14096 17536
rect 14051 17496 14096 17524
rect 12805 17487 12863 17493
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 16439 17527 16497 17533
rect 16439 17524 16451 17527
rect 16080 17496 16451 17524
rect 16080 17484 16086 17496
rect 16439 17493 16451 17496
rect 16485 17493 16497 17527
rect 16439 17487 16497 17493
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 17727 17527 17785 17533
rect 17727 17524 17739 17527
rect 17644 17496 17739 17524
rect 17644 17484 17650 17496
rect 17727 17493 17739 17496
rect 17773 17493 17785 17527
rect 18046 17524 18052 17536
rect 18007 17496 18052 17524
rect 17727 17487 17785 17493
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 18739 17527 18797 17533
rect 18739 17524 18751 17527
rect 18656 17496 18751 17524
rect 18656 17484 18662 17496
rect 18739 17493 18751 17496
rect 18785 17493 18797 17527
rect 19058 17524 19064 17536
rect 19019 17496 19064 17524
rect 18739 17487 18797 17493
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 1104 17434 20884 17456
rect 1104 17382 4648 17434
rect 4700 17382 4712 17434
rect 4764 17382 4776 17434
rect 4828 17382 4840 17434
rect 4892 17382 11982 17434
rect 12034 17382 12046 17434
rect 12098 17382 12110 17434
rect 12162 17382 12174 17434
rect 12226 17382 19315 17434
rect 19367 17382 19379 17434
rect 19431 17382 19443 17434
rect 19495 17382 19507 17434
rect 19559 17382 20884 17434
rect 1104 17360 20884 17382
rect 6362 17320 6368 17332
rect 6323 17292 6368 17320
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 8662 17320 8668 17332
rect 8575 17292 8668 17320
rect 8662 17280 8668 17292
rect 8720 17320 8726 17332
rect 9582 17320 9588 17332
rect 8720 17292 9588 17320
rect 8720 17280 8726 17292
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 10560 17292 10609 17320
rect 10560 17280 10566 17292
rect 10597 17289 10609 17292
rect 10643 17289 10655 17323
rect 10597 17283 10655 17289
rect 19199 17323 19257 17329
rect 19199 17289 19211 17323
rect 19245 17320 19257 17323
rect 19610 17320 19616 17332
rect 19245 17292 19616 17320
rect 19245 17289 19257 17292
rect 19199 17283 19257 17289
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 19702 17280 19708 17332
rect 19760 17320 19766 17332
rect 19760 17292 19805 17320
rect 19760 17280 19766 17292
rect 106 17212 112 17264
rect 164 17252 170 17264
rect 9263 17255 9321 17261
rect 9263 17252 9275 17255
rect 164 17224 9275 17252
rect 164 17212 170 17224
rect 9263 17221 9275 17224
rect 9309 17221 9321 17255
rect 9263 17215 9321 17221
rect 11330 17212 11336 17264
rect 11388 17252 11394 17264
rect 11388 17212 11411 17252
rect 11698 17212 11704 17264
rect 11756 17252 11762 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11756 17224 11805 17252
rect 11756 17212 11762 17224
rect 11793 17221 11805 17224
rect 11839 17252 11851 17255
rect 13354 17252 13360 17264
rect 11839 17224 13360 17252
rect 11839 17221 11851 17224
rect 11793 17215 11851 17221
rect 13354 17212 13360 17224
rect 13412 17252 13418 17264
rect 16298 17252 16304 17264
rect 13412 17224 16304 17252
rect 13412 17212 13418 17224
rect 16298 17212 16304 17224
rect 16356 17212 16362 17264
rect 7469 17187 7527 17193
rect 7469 17184 7481 17187
rect 6999 17156 7481 17184
rect 6999 17125 7027 17156
rect 7469 17153 7481 17156
rect 7515 17184 7527 17187
rect 9398 17184 9404 17196
rect 7515 17156 9404 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 9398 17144 9404 17156
rect 9456 17184 9462 17196
rect 10594 17184 10600 17196
rect 9456 17156 10600 17184
rect 9456 17144 9462 17156
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 11383 17184 11411 17212
rect 12710 17184 12716 17196
rect 11383 17156 12716 17184
rect 6984 17119 7042 17125
rect 6984 17085 6996 17119
rect 7030 17085 7042 17119
rect 6984 17079 7042 17085
rect 8018 17076 8024 17128
rect 8076 17116 8082 17128
rect 8148 17119 8206 17125
rect 8148 17116 8160 17119
rect 8076 17088 8160 17116
rect 8076 17076 8082 17088
rect 8148 17085 8160 17088
rect 8194 17116 8206 17119
rect 8941 17119 8999 17125
rect 8941 17116 8953 17119
rect 8194 17088 8953 17116
rect 8194 17085 8206 17088
rect 8148 17079 8206 17085
rect 8941 17085 8953 17088
rect 8987 17085 8999 17119
rect 8941 17079 8999 17085
rect 9192 17119 9250 17125
rect 9192 17085 9204 17119
rect 9238 17116 9250 17119
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9238 17088 9597 17116
rect 9238 17085 9250 17088
rect 9192 17079 9250 17085
rect 9585 17085 9597 17088
rect 9631 17116 9643 17119
rect 9950 17116 9956 17128
rect 9631 17088 9956 17116
rect 9631 17085 9643 17088
rect 9585 17079 9643 17085
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10204 17119 10262 17125
rect 10204 17085 10216 17119
rect 10250 17116 10262 17119
rect 10502 17116 10508 17128
rect 10250 17088 10508 17116
rect 10250 17085 10262 17088
rect 10204 17079 10262 17085
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 12452 17125 12480 17156
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 14090 17184 14096 17196
rect 14016 17156 14096 17184
rect 11368 17119 11426 17125
rect 11368 17116 11380 17119
rect 11231 17088 11380 17116
rect 7742 17048 7748 17060
rect 7703 17020 7748 17048
rect 7742 17008 7748 17020
rect 7800 17008 7806 17060
rect 8251 17051 8309 17057
rect 8251 17017 8263 17051
rect 8297 17048 8309 17051
rect 8297 17020 9260 17048
rect 8297 17017 8309 17020
rect 8251 17011 8309 17017
rect 9232 16992 9260 17020
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 11231 17048 11259 17088
rect 11368 17085 11380 17088
rect 11414 17116 11426 17119
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 11414 17088 12173 17116
rect 11414 17085 11426 17088
rect 11368 17079 11426 17085
rect 12161 17085 12173 17088
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 10836 17020 11259 17048
rect 12176 17048 12204 17079
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12584 17088 12909 17116
rect 12584 17076 12590 17088
rect 12897 17085 12909 17088
rect 12943 17116 12955 17119
rect 13814 17116 13820 17128
rect 12943 17088 13820 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 14016 17125 14044 17156
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 14424 17156 17141 17184
rect 14424 17144 14430 17156
rect 16735 17125 16763 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14001 17079 14059 17085
rect 14159 17088 14473 17116
rect 12802 17048 12808 17060
rect 12176 17020 12808 17048
rect 10836 17008 10842 17020
rect 12802 17008 12808 17020
rect 12860 17008 12866 17060
rect 13909 17051 13967 17057
rect 13909 17048 13921 17051
rect 13786 17020 13921 17048
rect 7055 16983 7113 16989
rect 7055 16949 7067 16983
rect 7101 16980 7113 16983
rect 7282 16980 7288 16992
rect 7101 16952 7288 16980
rect 7101 16949 7113 16952
rect 7055 16943 7113 16949
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 9214 16940 9220 16992
rect 9272 16940 9278 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10275 16983 10333 16989
rect 10275 16980 10287 16983
rect 10100 16952 10287 16980
rect 10100 16940 10106 16952
rect 10275 16949 10287 16952
rect 10321 16949 10333 16983
rect 10275 16943 10333 16949
rect 11471 16983 11529 16989
rect 11471 16949 11483 16983
rect 11517 16980 11529 16983
rect 11698 16980 11704 16992
rect 11517 16952 11704 16980
rect 11517 16949 11529 16952
rect 11471 16943 11529 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 12768 16952 13461 16980
rect 12768 16940 12774 16952
rect 13449 16949 13461 16952
rect 13495 16980 13507 16983
rect 13538 16980 13544 16992
rect 13495 16952 13544 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 13538 16940 13544 16952
rect 13596 16980 13602 16992
rect 13786 16980 13814 17020
rect 13909 17017 13921 17020
rect 13955 17048 13967 17051
rect 14159 17048 14187 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 16720 17119 16778 17125
rect 16720 17085 16732 17119
rect 16766 17085 16778 17119
rect 16720 17079 16778 17085
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18046 17116 18052 17128
rect 18104 17125 18110 17128
rect 18104 17119 18142 17125
rect 17828 17088 18052 17116
rect 17828 17076 17834 17088
rect 18046 17076 18052 17088
rect 18130 17085 18142 17119
rect 19058 17116 19064 17128
rect 19019 17088 19064 17116
rect 18104 17079 18142 17085
rect 18104 17076 18110 17079
rect 19058 17076 19064 17088
rect 19116 17076 19122 17128
rect 13955 17020 14187 17048
rect 16807 17051 16865 17057
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 16807 17017 16819 17051
rect 16853 17048 16865 17051
rect 18414 17048 18420 17060
rect 16853 17020 18420 17048
rect 16853 17017 16865 17020
rect 16807 17011 16865 17017
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 13596 16952 13814 16980
rect 14277 16983 14335 16989
rect 13596 16940 13602 16952
rect 14277 16949 14289 16983
rect 14323 16980 14335 16983
rect 14366 16980 14372 16992
rect 14323 16952 14372 16980
rect 14323 16949 14335 16952
rect 14277 16943 14335 16949
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 15286 16940 15292 16992
rect 15344 16980 15350 16992
rect 15565 16983 15623 16989
rect 15565 16980 15577 16983
rect 15344 16952 15577 16980
rect 15344 16940 15350 16952
rect 15565 16949 15577 16952
rect 15611 16949 15623 16983
rect 15565 16943 15623 16949
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 17589 16983 17647 16989
rect 17589 16980 17601 16983
rect 17460 16952 17601 16980
rect 17460 16940 17466 16952
rect 17589 16949 17601 16952
rect 17635 16949 17647 16983
rect 17589 16943 17647 16949
rect 18187 16983 18245 16989
rect 18187 16949 18199 16983
rect 18233 16980 18245 16983
rect 18506 16980 18512 16992
rect 18233 16952 18512 16980
rect 18233 16949 18245 16952
rect 18187 16943 18245 16949
rect 18506 16940 18512 16952
rect 18564 16940 18570 16992
rect 18690 16980 18696 16992
rect 18651 16952 18696 16980
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 1104 16890 20884 16912
rect 1104 16838 8315 16890
rect 8367 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 15648 16890
rect 15700 16838 15712 16890
rect 15764 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 20884 16890
rect 1104 16816 20884 16838
rect 8665 16779 8723 16785
rect 8665 16745 8677 16779
rect 8711 16776 8723 16779
rect 9766 16776 9772 16788
rect 8711 16748 9772 16776
rect 8711 16745 8723 16748
rect 8665 16739 8723 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 12342 16776 12348 16788
rect 12303 16748 12348 16776
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 13906 16776 13912 16788
rect 13867 16748 13912 16776
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 19245 16779 19303 16785
rect 19245 16745 19257 16779
rect 19291 16776 19303 16779
rect 19518 16776 19524 16788
rect 19291 16748 19524 16776
rect 19291 16745 19303 16748
rect 19245 16739 19303 16745
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 10413 16711 10471 16717
rect 10413 16708 10425 16711
rect 2096 16680 10425 16708
rect 2096 16668 2102 16680
rect 10413 16677 10425 16680
rect 10459 16677 10471 16711
rect 10413 16671 10471 16677
rect 5236 16643 5294 16649
rect 5236 16609 5248 16643
rect 5282 16640 5294 16643
rect 5534 16640 5540 16652
rect 5282 16612 5540 16640
rect 5282 16609 5294 16612
rect 5236 16603 5294 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 6248 16643 6306 16649
rect 6248 16609 6260 16643
rect 6294 16640 6306 16643
rect 6638 16640 6644 16652
rect 6294 16612 6644 16640
rect 6294 16609 6306 16612
rect 6248 16603 6306 16609
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 7260 16643 7318 16649
rect 7260 16609 7272 16643
rect 7306 16640 7318 16643
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 7306 16612 8493 16640
rect 7306 16609 7318 16612
rect 7260 16603 7318 16609
rect 8481 16609 8493 16612
rect 8527 16640 8539 16643
rect 8754 16640 8760 16652
rect 8527 16612 8760 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10134 16640 10140 16652
rect 9723 16612 10140 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 12710 16640 12716 16652
rect 12667 16612 12716 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16572 10103 16575
rect 10226 16572 10232 16584
rect 10091 16544 10232 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 12360 16572 12388 16603
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 13722 16640 13728 16652
rect 13683 16612 13728 16640
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 13998 16600 14004 16652
rect 14056 16640 14062 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 14056 16612 14105 16640
rect 14056 16600 14062 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16114 16640 16120 16652
rect 15979 16612 16120 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 18690 16600 18696 16652
rect 18748 16640 18754 16652
rect 19061 16643 19119 16649
rect 19061 16640 19073 16643
rect 18748 16612 19073 16640
rect 18748 16600 18754 16612
rect 19061 16609 19073 16612
rect 19107 16640 19119 16643
rect 19610 16640 19616 16652
rect 19107 16612 19616 16640
rect 19107 16609 19119 16612
rect 19061 16603 19119 16609
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 12894 16572 12900 16584
rect 12360 16544 12900 16572
rect 12894 16532 12900 16544
rect 12952 16532 12958 16584
rect 14918 16532 14924 16584
rect 14976 16572 14982 16584
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 14976 16544 15301 16572
rect 14976 16532 14982 16544
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 16850 16572 16856 16584
rect 16811 16544 16856 16572
rect 15289 16535 15347 16541
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 17126 16532 17132 16584
rect 17184 16572 17190 16584
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 17184 16544 17877 16572
rect 17184 16532 17190 16544
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 9401 16507 9459 16513
rect 9401 16504 9413 16507
rect 8312 16476 9413 16504
rect 5307 16439 5365 16445
rect 5307 16405 5319 16439
rect 5353 16436 5365 16439
rect 5442 16436 5448 16448
rect 5353 16408 5448 16436
rect 5353 16405 5365 16408
rect 5307 16399 5365 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6319 16439 6377 16445
rect 6319 16405 6331 16439
rect 6365 16436 6377 16439
rect 6730 16436 6736 16448
rect 6365 16408 6736 16436
rect 6365 16405 6377 16408
rect 6319 16399 6377 16405
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7331 16439 7389 16445
rect 7331 16436 7343 16439
rect 6972 16408 7343 16436
rect 6972 16396 6978 16408
rect 7331 16405 7343 16408
rect 7377 16405 7389 16439
rect 7331 16399 7389 16405
rect 7926 16396 7932 16448
rect 7984 16436 7990 16448
rect 8312 16445 8340 16476
rect 9401 16473 9413 16476
rect 9447 16504 9459 16507
rect 9815 16507 9873 16513
rect 9815 16504 9827 16507
rect 9447 16476 9827 16504
rect 9447 16473 9459 16476
rect 9401 16467 9459 16473
rect 9815 16473 9827 16476
rect 9861 16473 9873 16507
rect 9815 16467 9873 16473
rect 8297 16439 8355 16445
rect 8297 16436 8309 16439
rect 7984 16408 8309 16436
rect 7984 16396 7990 16408
rect 8297 16405 8309 16408
rect 8343 16405 8355 16439
rect 9030 16436 9036 16448
rect 8991 16408 9036 16436
rect 8297 16399 8355 16405
rect 9030 16396 9036 16408
rect 9088 16436 9094 16448
rect 9953 16439 10011 16445
rect 9953 16436 9965 16439
rect 9088 16408 9965 16436
rect 9088 16396 9094 16408
rect 9953 16405 9965 16408
rect 9999 16405 10011 16439
rect 9953 16399 10011 16405
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 13446 16436 13452 16448
rect 13219 16408 13452 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 1104 16346 20884 16368
rect 1104 16294 4648 16346
rect 4700 16294 4712 16346
rect 4764 16294 4776 16346
rect 4828 16294 4840 16346
rect 4892 16294 11982 16346
rect 12034 16294 12046 16346
rect 12098 16294 12110 16346
rect 12162 16294 12174 16346
rect 12226 16294 19315 16346
rect 19367 16294 19379 16346
rect 19431 16294 19443 16346
rect 19495 16294 19507 16346
rect 19559 16294 20884 16346
rect 1104 16272 20884 16294
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6638 16232 6644 16244
rect 6319 16204 6644 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 8021 16235 8079 16241
rect 8021 16201 8033 16235
rect 8067 16232 8079 16235
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 8067 16204 8309 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8297 16201 8309 16204
rect 8343 16232 8355 16235
rect 9306 16232 9312 16244
rect 8343 16204 9312 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 13722 16232 13728 16244
rect 10652 16204 13728 16232
rect 10652 16192 10658 16204
rect 13722 16192 13728 16204
rect 13780 16232 13786 16244
rect 14829 16235 14887 16241
rect 14829 16232 14841 16235
rect 13780 16204 14841 16232
rect 13780 16192 13786 16204
rect 14829 16201 14841 16204
rect 14875 16232 14887 16235
rect 16758 16232 16764 16244
rect 14875 16204 16764 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 19610 16232 19616 16244
rect 19571 16204 19616 16232
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 106 16124 112 16176
rect 164 16164 170 16176
rect 3651 16167 3709 16173
rect 3651 16164 3663 16167
rect 164 16136 3663 16164
rect 164 16124 170 16136
rect 3651 16133 3663 16136
rect 3697 16133 3709 16167
rect 5902 16164 5908 16176
rect 3651 16127 3709 16133
rect 4126 16136 5908 16164
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1535 16099 1593 16105
rect 1535 16096 1547 16099
rect 1360 16068 1547 16096
rect 1360 16056 1366 16068
rect 1535 16065 1547 16068
rect 1581 16065 1593 16099
rect 1535 16059 1593 16065
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16096 2007 16099
rect 4126 16096 4154 16136
rect 5902 16124 5908 16136
rect 5960 16124 5966 16176
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 8895 16167 8953 16173
rect 8895 16164 8907 16167
rect 7984 16136 8907 16164
rect 7984 16124 7990 16136
rect 8895 16133 8907 16136
rect 8941 16133 8953 16167
rect 9030 16164 9036 16176
rect 8991 16136 9036 16164
rect 8895 16127 8953 16133
rect 9030 16124 9036 16136
rect 9088 16124 9094 16176
rect 13280 16136 14044 16164
rect 1995 16068 4154 16096
rect 4847 16099 4905 16105
rect 1995 16065 2007 16068
rect 1949 16059 2007 16065
rect 4847 16065 4859 16099
rect 4893 16096 4905 16099
rect 6178 16096 6184 16108
rect 4893 16068 6184 16096
rect 4893 16065 4905 16068
rect 4847 16059 4905 16065
rect 1448 16031 1506 16037
rect 1448 15997 1460 16031
rect 1494 16028 1506 16031
rect 1964 16028 1992 16059
rect 6178 16056 6184 16068
rect 6236 16056 6242 16108
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16096 7343 16099
rect 8754 16096 8760 16108
rect 7331 16068 8760 16096
rect 7331 16065 7343 16068
rect 7285 16059 7343 16065
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9306 16096 9312 16108
rect 9171 16068 9312 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9306 16056 9312 16068
rect 9364 16096 9370 16108
rect 10226 16096 10232 16108
rect 9364 16068 10232 16096
rect 9364 16056 9370 16068
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 13280 16105 13308 16136
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 11348 16068 13277 16096
rect 1494 16000 1992 16028
rect 2568 16031 2626 16037
rect 1494 15997 1506 16000
rect 1448 15991 1506 15997
rect 2568 15997 2580 16031
rect 2614 16028 2626 16031
rect 3580 16031 3638 16037
rect 2614 16000 3096 16028
rect 2614 15997 2626 16000
rect 2568 15991 2626 15997
rect 2639 15895 2697 15901
rect 2639 15861 2651 15895
rect 2685 15892 2697 15895
rect 2866 15892 2872 15904
rect 2685 15864 2872 15892
rect 2685 15861 2697 15864
rect 2639 15855 2697 15861
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 3068 15901 3096 16000
rect 3580 15997 3592 16031
rect 3626 16028 3638 16031
rect 3626 16000 4108 16028
rect 3626 15997 3638 16000
rect 3580 15991 3638 15997
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15892 3111 15895
rect 3970 15892 3976 15904
rect 3099 15864 3976 15892
rect 3099 15861 3111 15864
rect 3053 15855 3111 15861
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 4080 15901 4108 16000
rect 4522 15988 4528 16040
rect 4580 16028 4586 16040
rect 4744 16031 4802 16037
rect 4744 16028 4756 16031
rect 4580 16000 4756 16028
rect 4580 15988 4586 16000
rect 4744 15997 4756 16000
rect 4790 16028 4802 16031
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 4790 16000 5181 16028
rect 4790 15997 4802 16000
rect 4744 15991 4802 15997
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5718 16028 5724 16040
rect 5682 16000 5724 16028
rect 5169 15991 5227 15997
rect 5718 15988 5724 16000
rect 5776 16037 5782 16040
rect 5776 16031 5830 16037
rect 5776 15997 5784 16031
rect 5818 16028 5830 16031
rect 6638 16028 6644 16040
rect 5818 16000 6644 16028
rect 5818 15997 5830 16000
rect 5776 15991 5830 15997
rect 5776 15988 5782 15991
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 7812 16031 7870 16037
rect 7812 15997 7824 16031
rect 7858 16028 7870 16031
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7858 16000 8033 16028
rect 7858 15997 7870 16000
rect 7812 15991 7870 15997
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 9861 16031 9919 16037
rect 9861 15997 9873 16031
rect 9907 16028 9919 16031
rect 10134 16028 10140 16040
rect 9907 16000 10140 16028
rect 9907 15997 9919 16000
rect 9861 15991 9919 15997
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10778 16028 10784 16040
rect 10739 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 11348 16037 11376 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 11333 16031 11391 16037
rect 11333 15997 11345 16031
rect 11379 15997 11391 16031
rect 11333 15991 11391 15997
rect 12504 16031 12562 16037
rect 12504 15997 12516 16031
rect 12550 16028 12562 16031
rect 12802 16028 12808 16040
rect 12550 16000 12808 16028
rect 12550 15997 12562 16000
rect 12504 15991 12562 15997
rect 5859 15963 5917 15969
rect 5859 15929 5871 15963
rect 5905 15960 5917 15963
rect 6822 15960 6828 15972
rect 5905 15932 6828 15960
rect 5905 15929 5917 15932
rect 5859 15923 5917 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 7653 15963 7711 15969
rect 7653 15929 7665 15963
rect 7699 15960 7711 15963
rect 8662 15960 8668 15972
rect 7699 15932 8668 15960
rect 7699 15929 7711 15932
rect 7653 15923 7711 15929
rect 8662 15920 8668 15932
rect 8720 15960 8726 15972
rect 8757 15963 8815 15969
rect 8757 15960 8769 15963
rect 8720 15932 8769 15960
rect 8720 15920 8726 15932
rect 8757 15929 8769 15932
rect 8803 15929 8815 15963
rect 9490 15960 9496 15972
rect 9451 15932 9496 15960
rect 8757 15923 8815 15929
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 10689 15963 10747 15969
rect 10689 15929 10701 15963
rect 10735 15960 10747 15963
rect 11348 15960 11376 15991
rect 12802 15988 12808 16000
rect 12860 16028 12866 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12860 16000 12909 16028
rect 12860 15988 12866 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 13446 16028 13452 16040
rect 13407 16000 13452 16028
rect 12897 15991 12955 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 14016 16037 14044 16136
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 16209 16031 16267 16037
rect 16209 15997 16221 16031
rect 16255 16028 16267 16031
rect 16298 16028 16304 16040
rect 16255 16000 16304 16028
rect 16255 15997 16267 16000
rect 16209 15991 16267 15997
rect 11422 15960 11428 15972
rect 10735 15932 11428 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 11422 15920 11428 15932
rect 11480 15920 11486 15972
rect 11517 15963 11575 15969
rect 11517 15929 11529 15963
rect 11563 15960 11575 15963
rect 11606 15960 11612 15972
rect 11563 15932 11612 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 11606 15920 11612 15932
rect 11664 15920 11670 15972
rect 12710 15960 12716 15972
rect 12084 15932 12716 15960
rect 4065 15895 4123 15901
rect 4065 15861 4077 15895
rect 4111 15892 4123 15895
rect 4338 15892 4344 15904
rect 4111 15864 4344 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6638 15892 6644 15904
rect 6599 15864 6644 15892
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 7883 15895 7941 15901
rect 7883 15861 7895 15895
rect 7929 15892 7941 15895
rect 8110 15892 8116 15904
rect 7929 15864 8116 15892
rect 7929 15861 7941 15864
rect 7883 15855 7941 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 8573 15895 8631 15901
rect 8573 15861 8585 15895
rect 8619 15892 8631 15895
rect 8846 15892 8852 15904
rect 8619 15864 8852 15892
rect 8619 15861 8631 15864
rect 8573 15855 8631 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 12084 15901 12112 15932
rect 12710 15920 12716 15932
rect 12768 15920 12774 15972
rect 14016 15904 14044 15991
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 16485 16031 16543 16037
rect 16485 15997 16497 16031
rect 16531 15997 16543 16031
rect 16485 15991 16543 15997
rect 14185 15963 14243 15969
rect 14185 15929 14197 15963
rect 14231 15960 14243 15963
rect 14274 15960 14280 15972
rect 14231 15932 14280 15960
rect 14231 15929 14243 15932
rect 14185 15923 14243 15929
rect 14274 15920 14280 15932
rect 14332 15920 14338 15972
rect 15381 15963 15439 15969
rect 15381 15929 15393 15963
rect 15427 15960 15439 15963
rect 16114 15960 16120 15972
rect 15427 15932 16120 15960
rect 15427 15929 15439 15932
rect 15381 15923 15439 15929
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 10376 15864 12081 15892
rect 10376 15852 10382 15864
rect 12069 15861 12081 15864
rect 12115 15861 12127 15895
rect 12069 15855 12127 15861
rect 12575 15895 12633 15901
rect 12575 15861 12587 15895
rect 12621 15892 12633 15895
rect 12802 15892 12808 15904
rect 12621 15864 12808 15892
rect 12621 15861 12633 15864
rect 12575 15855 12633 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 14056 15864 14473 15892
rect 14056 15852 14062 15864
rect 14461 15861 14473 15864
rect 14507 15861 14519 15895
rect 14461 15855 14519 15861
rect 15841 15895 15899 15901
rect 15841 15861 15853 15895
rect 15887 15892 15899 15895
rect 16500 15892 16528 15991
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 19188 16031 19246 16037
rect 19188 16028 19200 16031
rect 17368 16000 19200 16028
rect 17368 15988 17374 16000
rect 19188 15997 19200 16000
rect 19234 16028 19246 16031
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19234 16000 19993 16028
rect 19234 15997 19246 16000
rect 19188 15991 19246 15997
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 16666 15960 16672 15972
rect 16627 15932 16672 15960
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 19291 15963 19349 15969
rect 19291 15929 19303 15963
rect 19337 15960 19349 15963
rect 19702 15960 19708 15972
rect 19337 15932 19708 15960
rect 19337 15929 19349 15932
rect 19291 15923 19349 15929
rect 19702 15920 19708 15932
rect 19760 15920 19766 15972
rect 16942 15892 16948 15904
rect 15887 15864 16948 15892
rect 15887 15861 15899 15864
rect 15841 15855 15899 15861
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 18141 15895 18199 15901
rect 18141 15861 18153 15895
rect 18187 15892 18199 15895
rect 18874 15892 18880 15904
rect 18187 15864 18880 15892
rect 18187 15861 18199 15864
rect 18141 15855 18199 15861
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 1104 15802 20884 15824
rect 1104 15750 8315 15802
rect 8367 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 15648 15802
rect 15700 15750 15712 15802
rect 15764 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 20884 15802
rect 1104 15728 20884 15750
rect 5074 15688 5080 15700
rect 5035 15660 5080 15688
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 15427 15691 15485 15697
rect 15427 15657 15439 15691
rect 15473 15688 15485 15691
rect 18966 15688 18972 15700
rect 15473 15660 18972 15688
rect 15473 15657 15485 15660
rect 15427 15651 15485 15657
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19245 15691 19303 15697
rect 19245 15657 19257 15691
rect 19291 15688 19303 15691
rect 21542 15688 21548 15700
rect 19291 15660 21548 15688
rect 19291 15657 19303 15660
rect 19245 15651 19303 15657
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 3878 15580 3884 15632
rect 3936 15620 3942 15632
rect 7926 15620 7932 15632
rect 3936 15592 7932 15620
rect 3936 15580 3942 15592
rect 7926 15580 7932 15592
rect 7984 15620 7990 15632
rect 8021 15623 8079 15629
rect 8021 15620 8033 15623
rect 7984 15592 8033 15620
rect 7984 15580 7990 15592
rect 8021 15589 8033 15592
rect 8067 15589 8079 15623
rect 11330 15620 11336 15632
rect 8021 15583 8079 15589
rect 8312 15592 11336 15620
rect 2996 15555 3054 15561
rect 2996 15521 3008 15555
rect 3042 15521 3054 15555
rect 2996 15515 3054 15521
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15521 5135 15555
rect 5350 15552 5356 15564
rect 5311 15524 5356 15552
rect 5077 15515 5135 15521
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 3011 15416 3039 15515
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5092 15484 5120 15515
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 6512 15524 6561 15552
rect 6512 15512 6518 15524
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 6549 15515 6607 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8312 15484 8340 15592
rect 11330 15580 11336 15592
rect 11388 15580 11394 15632
rect 9766 15552 9772 15564
rect 9727 15524 9772 15552
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 11422 15552 11428 15564
rect 11383 15524 11428 15552
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 13722 15552 13728 15564
rect 13683 15524 13728 15552
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 13998 15552 14004 15564
rect 13959 15524 14004 15552
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 15356 15555 15414 15561
rect 15356 15521 15368 15555
rect 15402 15552 15414 15555
rect 15470 15552 15476 15564
rect 15402 15524 15476 15552
rect 15402 15521 15414 15524
rect 15356 15515 15414 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 16172 15524 16313 15552
rect 16172 15512 16178 15524
rect 16301 15521 16313 15524
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 16942 15552 16948 15564
rect 16899 15524 16948 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17770 15512 17776 15564
rect 17828 15552 17834 15564
rect 18084 15555 18142 15561
rect 18084 15552 18096 15555
rect 17828 15524 18096 15552
rect 17828 15512 17834 15524
rect 18084 15521 18096 15524
rect 18130 15521 18142 15555
rect 18084 15515 18142 15521
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15552 19119 15555
rect 19150 15552 19156 15564
rect 19107 15524 19156 15552
rect 19107 15521 19119 15524
rect 19061 15515 19119 15521
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 5040 15456 8340 15484
rect 5040 15444 5046 15456
rect 9030 15444 9036 15496
rect 9088 15444 9094 15496
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 3234 15416 3240 15428
rect 3011 15388 3240 15416
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 7098 15376 7104 15428
rect 7156 15416 7162 15428
rect 9048 15416 9076 15444
rect 9401 15419 9459 15425
rect 9401 15416 9413 15419
rect 7156 15388 9413 15416
rect 7156 15376 7162 15388
rect 9401 15385 9413 15388
rect 9447 15416 9459 15419
rect 9692 15416 9720 15447
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11296 15456 11345 15484
rect 11296 15444 11302 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 14182 15484 14188 15496
rect 14143 15456 14188 15484
rect 11333 15447 11391 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 17034 15484 17040 15496
rect 16995 15456 17040 15484
rect 17034 15444 17040 15456
rect 17092 15444 17098 15496
rect 9447 15388 9720 15416
rect 12437 15419 12495 15425
rect 9447 15385 9459 15388
rect 9401 15379 9459 15385
rect 12437 15385 12449 15419
rect 12483 15416 12495 15419
rect 12894 15416 12900 15428
rect 12483 15388 12900 15416
rect 12483 15385 12495 15388
rect 12437 15379 12495 15385
rect 12894 15376 12900 15388
rect 12952 15416 12958 15428
rect 13538 15416 13544 15428
rect 12952 15388 13544 15416
rect 12952 15376 12958 15388
rect 13538 15376 13544 15388
rect 13596 15416 13602 15428
rect 17402 15416 17408 15428
rect 13596 15388 17408 15416
rect 13596 15376 13602 15388
rect 17402 15376 17408 15388
rect 17460 15376 17466 15428
rect 3099 15351 3157 15357
rect 3099 15317 3111 15351
rect 3145 15348 3157 15351
rect 4246 15348 4252 15360
rect 3145 15320 4252 15348
rect 3145 15317 3157 15320
rect 3099 15311 3157 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 6963 15320 9137 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 9125 15317 9137 15320
rect 9171 15348 9183 15351
rect 9306 15348 9312 15360
rect 9171 15320 9312 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 14458 15348 14464 15360
rect 14419 15320 14464 15348
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 16025 15351 16083 15357
rect 16025 15317 16037 15351
rect 16071 15348 16083 15351
rect 16298 15348 16304 15360
rect 16071 15320 16304 15348
rect 16071 15317 16083 15320
rect 16025 15311 16083 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18187 15351 18245 15357
rect 18187 15348 18199 15351
rect 18012 15320 18199 15348
rect 18012 15308 18018 15320
rect 18187 15317 18199 15320
rect 18233 15317 18245 15351
rect 18187 15311 18245 15317
rect 1104 15258 20884 15280
rect 1104 15206 4648 15258
rect 4700 15206 4712 15258
rect 4764 15206 4776 15258
rect 4828 15206 4840 15258
rect 4892 15206 11982 15258
rect 12034 15206 12046 15258
rect 12098 15206 12110 15258
rect 12162 15206 12174 15258
rect 12226 15206 19315 15258
rect 19367 15206 19379 15258
rect 19431 15206 19443 15258
rect 19495 15206 19507 15258
rect 19559 15206 20884 15258
rect 1104 15184 20884 15206
rect 2041 15147 2099 15153
rect 2041 15113 2053 15147
rect 2087 15144 2099 15147
rect 2314 15144 2320 15156
rect 2087 15116 2320 15144
rect 2087 15113 2099 15116
rect 2041 15107 2099 15113
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1854 14940 1860 14952
rect 1443 14912 1860 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1854 14900 1860 14912
rect 1912 14940 1918 14952
rect 2056 14940 2084 15107
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 2593 15147 2651 15153
rect 2593 15113 2605 15147
rect 2639 15144 2651 15147
rect 3234 15144 3240 15156
rect 2639 15116 3240 15144
rect 2639 15113 2651 15116
rect 2593 15107 2651 15113
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 7892 15116 8125 15144
rect 7892 15104 7898 15116
rect 8113 15113 8125 15116
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9766 15144 9772 15156
rect 9456 15116 9772 15144
rect 9456 15104 9462 15116
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 14090 15144 14096 15156
rect 13786 15116 14096 15144
rect 2332 15076 2360 15104
rect 13786 15088 13814 15116
rect 14090 15104 14096 15116
rect 14148 15144 14154 15156
rect 14185 15147 14243 15153
rect 14185 15144 14197 15147
rect 14148 15116 14197 15144
rect 14148 15104 14154 15116
rect 14185 15113 14197 15116
rect 14231 15113 14243 15147
rect 17402 15144 17408 15156
rect 17363 15116 17408 15144
rect 14185 15107 14243 15113
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 17770 15144 17776 15156
rect 17731 15116 17776 15144
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 19150 15144 19156 15156
rect 19111 15116 19156 15144
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 4522 15076 4528 15088
rect 2332 15048 4528 15076
rect 4522 15036 4528 15048
rect 4580 15036 4586 15088
rect 10778 15076 10784 15088
rect 8772 15048 10784 15076
rect 4430 14968 4436 15020
rect 4488 15008 4494 15020
rect 6454 15008 6460 15020
rect 4488 14980 6460 15008
rect 4488 14968 4494 14980
rect 6454 14968 6460 14980
rect 6512 14968 6518 15020
rect 8772 15008 8800 15048
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 13722 15036 13728 15088
rect 13780 15048 13814 15088
rect 13909 15079 13967 15085
rect 13780 15036 13786 15048
rect 13909 15045 13921 15079
rect 13955 15076 13967 15079
rect 13998 15076 14004 15088
rect 13955 15048 14004 15076
rect 13955 15045 13967 15048
rect 13909 15039 13967 15045
rect 13998 15036 14004 15048
rect 14056 15076 14062 15088
rect 18322 15076 18328 15088
rect 14056 15048 18328 15076
rect 14056 15036 14062 15048
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 8938 15008 8944 15020
rect 8680 14980 8800 15008
rect 8899 14980 8944 15008
rect 2958 14940 2964 14952
rect 1912 14912 2084 14940
rect 2871 14912 2964 14940
rect 1912 14900 1918 14912
rect 2958 14900 2964 14912
rect 3016 14940 3022 14952
rect 3145 14943 3203 14949
rect 3145 14940 3157 14943
rect 3016 14912 3157 14940
rect 3016 14900 3022 14912
rect 3145 14909 3157 14912
rect 3191 14909 3203 14943
rect 3145 14903 3203 14909
rect 3602 14900 3608 14952
rect 3660 14940 3666 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3660 14912 4077 14940
rect 3660 14900 3666 14912
rect 4065 14909 4077 14912
rect 4111 14940 4123 14943
rect 5258 14940 5264 14952
rect 4111 14912 5264 14940
rect 4111 14909 4123 14912
rect 4065 14903 4123 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14909 5503 14943
rect 5445 14903 5503 14909
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 7190 14940 7196 14952
rect 7147 14912 7196 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 3050 14872 3056 14884
rect 3011 14844 3056 14872
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 5350 14872 5356 14884
rect 4816 14844 5356 14872
rect 106 14764 112 14816
rect 164 14804 170 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 164 14776 1593 14804
rect 164 14764 170 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 4522 14804 4528 14816
rect 4483 14776 4528 14804
rect 1581 14767 1639 14773
rect 4522 14764 4528 14776
rect 4580 14804 4586 14816
rect 4816 14813 4844 14844
rect 5350 14832 5356 14844
rect 5408 14872 5414 14884
rect 5460 14872 5488 14903
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 6089 14875 6147 14881
rect 6089 14872 6101 14875
rect 5408 14844 6101 14872
rect 5408 14832 5414 14844
rect 6089 14841 6101 14844
rect 6135 14872 6147 14875
rect 7300 14872 7328 14903
rect 7926 14900 7932 14952
rect 7984 14940 7990 14952
rect 8680 14949 8708 14980
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 9490 15008 9496 15020
rect 9364 14980 9496 15008
rect 9364 14968 9370 14980
rect 9490 14968 9496 14980
rect 9548 15008 9554 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 9548 14980 10977 15008
rect 9548 14968 9554 14980
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 7984 14912 8677 14940
rect 7984 14900 7990 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8846 14940 8852 14952
rect 8807 14912 8852 14940
rect 8665 14903 8723 14909
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 10152 14949 10180 14980
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 14458 15008 14464 15020
rect 10965 14971 11023 14977
rect 13786 14980 14464 15008
rect 13786 14952 13814 14980
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 14700 14980 15884 15008
rect 14700 14968 14706 14980
rect 10137 14943 10195 14949
rect 10137 14909 10149 14943
rect 10183 14909 10195 14943
rect 10502 14940 10508 14952
rect 10463 14912 10508 14940
rect 10137 14903 10195 14909
rect 10502 14900 10508 14912
rect 10560 14900 10566 14952
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 11330 14940 11336 14952
rect 10836 14912 11336 14940
rect 10836 14900 10842 14912
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 13786 14940 13820 14952
rect 13587 14912 13820 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 15856 14949 15884 14980
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 17828 14980 19691 15008
rect 17828 14968 17834 14980
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15841 14943 15899 14949
rect 15151 14912 15516 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 12894 14872 12900 14884
rect 6135 14844 7328 14872
rect 12855 14844 12900 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 12894 14832 12900 14844
rect 12952 14832 12958 14884
rect 12989 14875 13047 14881
rect 12989 14841 13001 14875
rect 13035 14841 13047 14875
rect 12989 14835 13047 14841
rect 14553 14875 14611 14881
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 14642 14872 14648 14884
rect 14599 14844 14648 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 4801 14807 4859 14813
rect 4801 14804 4813 14807
rect 4580 14776 4813 14804
rect 4580 14764 4586 14776
rect 4801 14773 4813 14776
rect 4847 14773 4859 14807
rect 4801 14767 4859 14773
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5166 14804 5172 14816
rect 5123 14776 5172 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 6917 14807 6975 14813
rect 6917 14773 6929 14807
rect 6963 14804 6975 14807
rect 7006 14804 7012 14816
rect 6963 14776 7012 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 9088 14776 10057 14804
rect 9088 14764 9094 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 10045 14767 10103 14773
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 11333 14807 11391 14813
rect 11333 14804 11345 14807
rect 10468 14776 11345 14804
rect 10468 14764 10474 14776
rect 11333 14773 11345 14776
rect 11379 14804 11391 14807
rect 11422 14804 11428 14816
rect 11379 14776 11428 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12713 14807 12771 14813
rect 12713 14773 12725 14807
rect 12759 14804 12771 14807
rect 13004 14804 13032 14835
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 15488 14816 15516 14912
rect 15841 14909 15853 14943
rect 15887 14940 15899 14943
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15887 14912 16037 14940
rect 15887 14909 15899 14912
rect 15841 14903 15899 14909
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 17402 14900 17408 14952
rect 17460 14940 17466 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17460 14912 18061 14940
rect 17460 14900 17466 14912
rect 18049 14909 18061 14912
rect 18095 14940 18107 14943
rect 18230 14940 18236 14952
rect 18095 14912 18236 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 19663 14949 19691 14980
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18380 14912 18521 14940
rect 18380 14900 18386 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 19648 14943 19706 14949
rect 19648 14909 19660 14943
rect 19694 14940 19706 14943
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 19694 14912 20085 14940
rect 19694 14909 19706 14912
rect 19648 14903 19706 14909
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 20073 14903 20131 14909
rect 15930 14872 15936 14884
rect 15891 14844 15936 14872
rect 15930 14832 15936 14844
rect 15988 14832 15994 14884
rect 18782 14832 18788 14884
rect 18840 14872 18846 14884
rect 19751 14875 19809 14881
rect 19751 14872 19763 14875
rect 18840 14844 19763 14872
rect 18840 14832 18846 14844
rect 19751 14841 19763 14844
rect 19797 14841 19809 14875
rect 19751 14835 19809 14841
rect 13538 14804 13544 14816
rect 12759 14776 13544 14804
rect 12759 14773 12771 14776
rect 12713 14767 12771 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 15470 14804 15476 14816
rect 15431 14776 15476 14804
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17037 14807 17095 14813
rect 17037 14804 17049 14807
rect 17000 14776 17049 14804
rect 17000 14764 17006 14776
rect 17037 14773 17049 14776
rect 17083 14804 17095 14807
rect 17402 14804 17408 14816
rect 17083 14776 17408 14804
rect 17083 14773 17095 14776
rect 17037 14767 17095 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 18138 14804 18144 14816
rect 18099 14776 18144 14804
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 1104 14714 20884 14736
rect 1104 14662 8315 14714
rect 8367 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 15648 14714
rect 15700 14662 15712 14714
rect 15764 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 20884 14714
rect 1104 14640 20884 14662
rect 1670 14600 1676 14612
rect 1583 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14600 1734 14612
rect 5718 14600 5724 14612
rect 1728 14572 5724 14600
rect 1728 14560 1734 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6638 14600 6644 14612
rect 6595 14572 6644 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 11330 14600 11336 14612
rect 8987 14572 10548 14600
rect 11291 14572 11336 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 10520 14544 10548 14572
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 12894 14600 12900 14612
rect 12855 14572 12900 14600
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14642 14600 14648 14612
rect 14507 14572 14648 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 15930 14600 15936 14612
rect 15488 14572 15936 14600
rect 4522 14492 4528 14544
rect 4580 14532 4586 14544
rect 7466 14532 7472 14544
rect 4580 14504 5396 14532
rect 4580 14492 4586 14504
rect 2222 14464 2228 14476
rect 2183 14436 2228 14464
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 2740 14436 4813 14464
rect 2740 14424 2746 14436
rect 4801 14433 4813 14436
rect 4847 14464 4859 14467
rect 4982 14464 4988 14476
rect 4847 14436 4988 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5368 14473 5396 14504
rect 6748 14504 7472 14532
rect 6748 14473 6776 14504
rect 7466 14492 7472 14504
rect 7524 14532 7530 14544
rect 9306 14532 9312 14544
rect 7524 14504 9312 14532
rect 7524 14492 7530 14504
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 9490 14492 9496 14544
rect 9548 14532 9554 14544
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9548 14504 9873 14532
rect 9548 14492 9554 14504
rect 9861 14501 9873 14504
rect 9907 14501 9919 14535
rect 9861 14495 9919 14501
rect 10502 14492 10508 14544
rect 10560 14532 10566 14544
rect 10560 14504 10732 14532
rect 10560 14492 10566 14504
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14433 6975 14467
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 6917 14427 6975 14433
rect 5184 14328 5212 14427
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5316 14368 5457 14396
rect 5316 14356 5322 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 6932 14396 6960 14427
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 8619 14436 8708 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 7190 14396 7196 14408
rect 6512 14368 7196 14396
rect 6512 14356 6518 14368
rect 7190 14356 7196 14368
rect 7248 14396 7254 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7248 14368 7481 14396
rect 7248 14356 7254 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 8680 14340 8708 14436
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 9306 14396 9312 14408
rect 8803 14368 9312 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 10008 14368 10057 14396
rect 10008 14356 10014 14368
rect 10045 14365 10057 14368
rect 10091 14396 10103 14399
rect 10502 14396 10508 14408
rect 10091 14368 10508 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 5350 14328 5356 14340
rect 5184 14300 5356 14328
rect 5350 14288 5356 14300
rect 5408 14328 5414 14340
rect 5408 14300 7671 14328
rect 5408 14288 5414 14300
rect 2590 14260 2596 14272
rect 2551 14232 2596 14260
rect 2590 14220 2596 14232
rect 2648 14220 2654 14272
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3145 14263 3203 14269
rect 3145 14260 3157 14263
rect 2832 14232 3157 14260
rect 2832 14220 2838 14232
rect 3145 14229 3157 14232
rect 3191 14229 3203 14263
rect 7643 14260 7671 14300
rect 8662 14288 8668 14340
rect 8720 14328 8726 14340
rect 8846 14328 8852 14340
rect 8720 14300 8852 14328
rect 8720 14288 8726 14300
rect 8846 14288 8852 14300
rect 8904 14328 8910 14340
rect 10704 14337 10732 14504
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 12342 14532 12348 14544
rect 11848 14504 12348 14532
rect 11848 14492 11854 14504
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 13170 14532 13176 14544
rect 13131 14504 13176 14532
rect 13170 14492 13176 14504
rect 13228 14492 13234 14544
rect 13725 14535 13783 14541
rect 13725 14501 13737 14535
rect 13771 14532 13783 14535
rect 13814 14532 13820 14544
rect 13771 14504 13820 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 15102 14492 15108 14544
rect 15160 14532 15166 14544
rect 15488 14541 15516 14572
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 16942 14600 16948 14612
rect 16903 14572 16948 14600
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 17920 14572 18521 14600
rect 17920 14560 17926 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 15473 14535 15531 14541
rect 15473 14532 15485 14535
rect 15160 14504 15485 14532
rect 15160 14492 15166 14504
rect 15473 14501 15485 14504
rect 15519 14501 15531 14535
rect 15473 14495 15531 14501
rect 18141 14535 18199 14541
rect 18141 14501 18153 14535
rect 18187 14532 18199 14535
rect 18322 14532 18328 14544
rect 18187 14504 18328 14532
rect 18187 14501 18199 14504
rect 18141 14495 18199 14501
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 10778 14424 10784 14476
rect 10836 14464 10842 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 10836 14436 11253 14464
rect 10836 14424 10842 14436
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 11480 14436 11713 14464
rect 11480 14424 11486 14436
rect 11701 14433 11713 14436
rect 11747 14433 11759 14467
rect 11701 14427 11759 14433
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 16758 14464 16764 14476
rect 16540 14436 16764 14464
rect 16540 14424 16546 14436
rect 16758 14424 16764 14436
rect 16816 14464 16822 14476
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16816 14436 16865 14464
rect 16816 14424 16822 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 17402 14464 17408 14476
rect 17363 14436 17408 14464
rect 16853 14427 16911 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18288 14436 18429 14464
rect 18288 14424 18294 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18966 14464 18972 14476
rect 18927 14436 18972 14464
rect 18417 14427 18475 14433
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12618 14396 12624 14408
rect 11848 14368 12624 14396
rect 11848 14356 11854 14368
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 13081 14399 13139 14405
rect 13081 14396 13093 14399
rect 12860 14368 13093 14396
rect 12860 14356 12866 14368
rect 13081 14365 13093 14368
rect 13127 14365 13139 14399
rect 15378 14396 15384 14408
rect 15339 14368 15384 14396
rect 13081 14359 13139 14365
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15528 14368 15669 14396
rect 15528 14356 15534 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 9033 14331 9091 14337
rect 9033 14328 9045 14331
rect 8904 14300 9045 14328
rect 8904 14288 8910 14300
rect 9033 14297 9045 14300
rect 9079 14297 9091 14331
rect 9033 14291 9091 14297
rect 10689 14331 10747 14337
rect 10689 14297 10701 14331
rect 10735 14328 10747 14331
rect 13722 14328 13728 14340
rect 10735 14300 13728 14328
rect 10735 14297 10747 14300
rect 10689 14291 10747 14297
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 14090 14288 14096 14340
rect 14148 14328 14154 14340
rect 16114 14328 16120 14340
rect 14148 14300 16120 14328
rect 14148 14288 14154 14300
rect 16114 14288 16120 14300
rect 16172 14328 16178 14340
rect 16301 14331 16359 14337
rect 16301 14328 16313 14331
rect 16172 14300 16313 14328
rect 16172 14288 16178 14300
rect 16301 14297 16313 14300
rect 16347 14297 16359 14331
rect 16301 14291 16359 14297
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 7643 14232 8953 14260
rect 3145 14223 3203 14229
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10836 14232 11161 14260
rect 10836 14220 10842 14232
rect 11149 14229 11161 14232
rect 11195 14260 11207 14263
rect 12710 14260 12716 14272
rect 11195 14232 12716 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 18322 14260 18328 14272
rect 13504 14232 18328 14260
rect 13504 14220 13510 14232
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 1104 14170 20884 14192
rect 1104 14118 4648 14170
rect 4700 14118 4712 14170
rect 4764 14118 4776 14170
rect 4828 14118 4840 14170
rect 4892 14118 11982 14170
rect 12034 14118 12046 14170
rect 12098 14118 12110 14170
rect 12162 14118 12174 14170
rect 12226 14118 19315 14170
rect 19367 14118 19379 14170
rect 19431 14118 19443 14170
rect 19495 14118 19507 14170
rect 19559 14118 20884 14170
rect 1104 14096 20884 14118
rect 3789 14059 3847 14065
rect 3789 14056 3801 14059
rect 2884 14028 3801 14056
rect 2590 13948 2596 14000
rect 2648 13988 2654 14000
rect 2884 13997 2912 14028
rect 3789 14025 3801 14028
rect 3835 14025 3847 14059
rect 3789 14019 3847 14025
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 8294 14056 8300 14068
rect 7708 14028 8300 14056
rect 7708 14016 7714 14028
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 8352 14028 9720 14056
rect 8352 14016 8358 14028
rect 2869 13991 2927 13997
rect 2869 13988 2881 13991
rect 2648 13960 2881 13988
rect 2648 13948 2654 13960
rect 2869 13957 2881 13960
rect 2915 13957 2927 13991
rect 2869 13951 2927 13957
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 5718 13988 5724 14000
rect 3568 13960 5724 13988
rect 3568 13948 3574 13960
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 8113 13991 8171 13997
rect 8113 13957 8125 13991
rect 8159 13988 8171 13991
rect 8662 13988 8668 14000
rect 8159 13960 8668 13988
rect 8159 13957 8171 13960
rect 8113 13951 8171 13957
rect 8662 13948 8668 13960
rect 8720 13948 8726 14000
rect 8754 13948 8760 14000
rect 8812 13988 8818 14000
rect 9582 13988 9588 14000
rect 8812 13960 9588 13988
rect 8812 13948 8818 13960
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 9692 13988 9720 14028
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 9824 14028 10149 14056
rect 9824 14016 9830 14028
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 10137 14019 10195 14025
rect 12575 14059 12633 14065
rect 12575 14025 12587 14059
rect 12621 14056 12633 14059
rect 12894 14056 12900 14068
rect 12621 14028 12900 14056
rect 12621 14025 12633 14028
rect 12575 14019 12633 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 12989 14059 13047 14065
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 13081 14059 13139 14065
rect 13081 14056 13093 14059
rect 13035 14028 13093 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13081 14025 13093 14028
rect 13127 14056 13139 14059
rect 13354 14056 13360 14068
rect 13127 14028 13360 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14642 14056 14648 14068
rect 14415 14028 14648 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15102 14056 15108 14068
rect 15063 14028 15108 14056
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 16577 14059 16635 14065
rect 16577 14056 16589 14059
rect 16540 14028 16589 14056
rect 16540 14016 16546 14028
rect 16577 14025 16589 14028
rect 16623 14025 16635 14059
rect 16577 14019 16635 14025
rect 9858 13988 9864 14000
rect 9692 13960 9864 13988
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 10318 13988 10324 14000
rect 10203 13960 10324 13988
rect 3234 13880 3240 13932
rect 3292 13920 3298 13932
rect 5350 13920 5356 13932
rect 3292 13892 3924 13920
rect 3292 13880 3298 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 2774 13852 2780 13864
rect 2188 13824 2780 13852
rect 2188 13812 2194 13824
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 3053 13855 3111 13861
rect 3053 13852 3065 13855
rect 3016 13824 3065 13852
rect 3016 13812 3022 13824
rect 3053 13821 3065 13824
rect 3099 13821 3111 13855
rect 3510 13852 3516 13864
rect 3471 13824 3516 13852
rect 3053 13815 3111 13821
rect 2222 13784 2228 13796
rect 2183 13756 2228 13784
rect 2222 13744 2228 13756
rect 2280 13744 2286 13796
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 2593 13719 2651 13725
rect 2593 13716 2605 13719
rect 2556 13688 2605 13716
rect 2556 13676 2562 13688
rect 2593 13685 2605 13688
rect 2639 13716 2651 13719
rect 3068 13716 3096 13815
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3896 13852 3924 13892
rect 5276 13892 5356 13920
rect 4341 13855 4399 13861
rect 4341 13852 4353 13855
rect 3896 13824 4353 13852
rect 4341 13821 4353 13824
rect 4387 13852 4399 13855
rect 4982 13852 4988 13864
rect 4387 13824 4988 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 4982 13812 4988 13824
rect 5040 13852 5046 13864
rect 5276 13861 5304 13892
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 7466 13920 7472 13932
rect 7300 13892 7472 13920
rect 7300 13861 7328 13892
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13920 8539 13923
rect 8846 13920 8852 13932
rect 8527 13892 8852 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 10203 13920 10231 13960
rect 10318 13948 10324 13960
rect 10376 13948 10382 14000
rect 10502 13948 10508 14000
rect 10560 13988 10566 14000
rect 10965 13991 11023 13997
rect 10965 13988 10977 13991
rect 10560 13960 10977 13988
rect 10560 13948 10566 13960
rect 10965 13957 10977 13960
rect 11011 13957 11023 13991
rect 10965 13951 11023 13957
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 12802 13988 12808 14000
rect 12299 13960 12808 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 14737 13991 14795 13997
rect 14737 13957 14749 13991
rect 14783 13988 14795 13991
rect 15378 13988 15384 14000
rect 14783 13960 15384 13988
rect 14783 13957 14795 13960
rect 14737 13951 14795 13957
rect 15378 13948 15384 13960
rect 15436 13948 15442 14000
rect 16758 13948 16764 14000
rect 16816 13988 16822 14000
rect 16899 13991 16957 13997
rect 16816 13948 16850 13988
rect 16899 13957 16911 13991
rect 16945 13988 16957 13991
rect 20622 13988 20628 14000
rect 16945 13960 20628 13988
rect 16945 13957 16957 13960
rect 16899 13951 16957 13957
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 9824 13892 10231 13920
rect 10413 13923 10471 13929
rect 9824 13880 9830 13892
rect 10413 13889 10425 13923
rect 10459 13920 10471 13923
rect 10778 13920 10784 13932
rect 10459 13892 10784 13920
rect 10459 13889 10471 13892
rect 10413 13883 10471 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11422 13920 11428 13932
rect 11335 13892 11428 13920
rect 11422 13880 11428 13892
rect 11480 13920 11486 13932
rect 13262 13920 13268 13932
rect 11480 13892 13268 13920
rect 11480 13880 11486 13892
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13786 13892 15884 13920
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5040 13824 5273 13852
rect 5040 13812 5046 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5261 13815 5319 13821
rect 5362 13824 5641 13852
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 5077 13787 5135 13793
rect 5077 13784 5089 13787
rect 3476 13756 5089 13784
rect 3476 13744 3482 13756
rect 5077 13753 5089 13756
rect 5123 13784 5135 13787
rect 5362 13784 5390 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 5629 13815 5687 13821
rect 6472 13824 7297 13852
rect 5123 13756 5390 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 2639 13688 3096 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4617 13719 4675 13725
rect 4617 13716 4629 13719
rect 4580 13688 4629 13716
rect 4580 13676 4586 13688
rect 4617 13685 4629 13688
rect 4663 13685 4675 13719
rect 5442 13716 5448 13728
rect 5403 13688 5448 13716
rect 4617 13679 4675 13685
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 6086 13676 6092 13728
rect 6144 13716 6150 13728
rect 6472 13725 6500 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13852 7619 13855
rect 7650 13852 7656 13864
rect 7607 13824 7656 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13852 8631 13855
rect 8754 13852 8760 13864
rect 8619 13824 8760 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 12504 13855 12562 13861
rect 12504 13821 12516 13855
rect 12550 13852 12562 13855
rect 12894 13852 12900 13864
rect 12550 13824 12900 13852
rect 12550 13821 12562 13824
rect 12504 13815 12562 13821
rect 12894 13812 12900 13824
rect 12952 13852 12958 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12952 13824 13093 13852
rect 12952 13812 12958 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13446 13852 13452 13864
rect 13407 13824 13452 13852
rect 13081 13815 13139 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 13786 13852 13814 13892
rect 15856 13861 15884 13892
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16482 13920 16488 13932
rect 16172 13892 16488 13920
rect 16172 13880 16178 13892
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16822 13861 16850 13948
rect 18322 13920 18328 13932
rect 18064 13892 18328 13920
rect 13596 13824 13814 13852
rect 15841 13855 15899 13861
rect 13596 13812 13602 13824
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15887 13824 16221 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16807 13855 16865 13861
rect 16807 13821 16819 13855
rect 16853 13821 16865 13855
rect 16807 13815 16865 13821
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 18064 13861 18092 13892
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18049 13855 18107 13861
rect 17460 13824 17632 13852
rect 17460 13812 17466 13824
rect 7742 13784 7748 13796
rect 7703 13756 7748 13784
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 10505 13787 10563 13793
rect 10505 13753 10517 13787
rect 10551 13753 10563 13787
rect 13770 13787 13828 13793
rect 13770 13784 13782 13787
rect 10505 13747 10563 13753
rect 13280 13756 13782 13784
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 6144 13688 6469 13716
rect 6144 13676 6150 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 6457 13679 6515 13685
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8904 13688 8953 13716
rect 8904 13676 8910 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 9490 13716 9496 13728
rect 9451 13688 9496 13716
rect 8941 13679 8999 13685
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 10520 13716 10548 13747
rect 10870 13716 10876 13728
rect 10520 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11793 13719 11851 13725
rect 11793 13685 11805 13719
rect 11839 13716 11851 13719
rect 12066 13716 12072 13728
rect 11839 13688 12072 13716
rect 11839 13685 11851 13688
rect 11793 13679 11851 13685
rect 12066 13676 12072 13688
rect 12124 13676 12130 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13280 13725 13308 13756
rect 13770 13753 13782 13756
rect 13816 13753 13828 13787
rect 13770 13747 13828 13753
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 15197 13787 15255 13793
rect 15197 13784 15209 13787
rect 14700 13756 15209 13784
rect 14700 13744 14706 13756
rect 15197 13753 15209 13756
rect 15243 13753 15255 13787
rect 15197 13747 15255 13753
rect 15470 13744 15476 13796
rect 15528 13784 15534 13796
rect 17494 13784 17500 13796
rect 15528 13756 17500 13784
rect 15528 13744 15534 13756
rect 17494 13744 17500 13756
rect 17552 13744 17558 13796
rect 17604 13784 17632 13824
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 18049 13815 18107 13821
rect 18156 13824 18521 13852
rect 18156 13784 18184 13824
rect 18509 13821 18521 13824
rect 18555 13852 18567 13855
rect 18966 13852 18972 13864
rect 18555 13824 18972 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 18966 13812 18972 13824
rect 19024 13852 19030 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 19024 13824 19073 13852
rect 19024 13812 19030 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 19648 13855 19706 13861
rect 19648 13852 19660 13855
rect 19208 13824 19660 13852
rect 19208 13812 19214 13824
rect 19648 13821 19660 13824
rect 19694 13852 19706 13855
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19694 13824 20085 13852
rect 19694 13821 19706 13824
rect 19648 13815 19706 13821
rect 20073 13821 20085 13824
rect 20119 13821 20131 13855
rect 20073 13815 20131 13821
rect 17604 13756 18184 13784
rect 13265 13719 13323 13725
rect 13265 13716 13277 13719
rect 12768 13688 13277 13716
rect 12768 13676 12774 13688
rect 13265 13685 13277 13688
rect 13311 13685 13323 13719
rect 13265 13679 13323 13685
rect 16114 13676 16120 13728
rect 16172 13716 16178 13728
rect 17221 13719 17279 13725
rect 17221 13716 17233 13719
rect 16172 13688 17233 13716
rect 16172 13676 16178 13688
rect 17221 13685 17233 13688
rect 17267 13716 17279 13719
rect 17604 13716 17632 13756
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 17267 13688 17785 13716
rect 17267 13685 17279 13688
rect 17221 13679 17279 13685
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 18138 13716 18144 13728
rect 18099 13688 18144 13716
rect 17773 13679 17831 13685
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 19610 13676 19616 13728
rect 19668 13716 19674 13728
rect 19751 13719 19809 13725
rect 19751 13716 19763 13719
rect 19668 13688 19763 13716
rect 19668 13676 19674 13688
rect 19751 13685 19763 13688
rect 19797 13685 19809 13719
rect 19751 13679 19809 13685
rect 1104 13626 20884 13648
rect 1104 13574 8315 13626
rect 8367 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 15648 13626
rect 15700 13574 15712 13626
rect 15764 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 20884 13626
rect 1104 13552 20884 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 1949 13515 2007 13521
rect 1949 13512 1961 13515
rect 1820 13484 1961 13512
rect 1820 13472 1826 13484
rect 1949 13481 1961 13484
rect 1995 13512 2007 13515
rect 3510 13512 3516 13524
rect 1995 13484 3516 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3786 13472 3792 13524
rect 3844 13512 3850 13524
rect 3844 13484 4384 13512
rect 3844 13472 3850 13484
rect 1397 13447 1455 13453
rect 1397 13413 1409 13447
rect 1443 13444 1455 13447
rect 3881 13447 3939 13453
rect 1443 13416 3601 13444
rect 1443 13413 1455 13416
rect 1397 13407 1455 13413
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 2240 13348 2421 13376
rect 2240 13240 2268 13348
rect 2409 13345 2421 13348
rect 2455 13345 2467 13379
rect 2958 13376 2964 13388
rect 2919 13348 2964 13376
rect 2409 13339 2467 13345
rect 2958 13336 2964 13348
rect 3016 13376 3022 13388
rect 3418 13376 3424 13388
rect 3016 13348 3424 13376
rect 3016 13336 3022 13348
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3326 13308 3332 13320
rect 3191 13280 3332 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3573 13308 3601 13416
rect 3881 13413 3893 13447
rect 3927 13444 3939 13447
rect 3970 13444 3976 13456
rect 3927 13416 3976 13444
rect 3927 13413 3939 13416
rect 3881 13407 3939 13413
rect 3970 13404 3976 13416
rect 4028 13444 4034 13456
rect 4249 13447 4307 13453
rect 4249 13444 4261 13447
rect 4028 13416 4261 13444
rect 4028 13404 4034 13416
rect 4249 13413 4261 13416
rect 4295 13413 4307 13447
rect 4356 13444 4384 13484
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 5040 13484 5181 13512
rect 5040 13472 5046 13484
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 5721 13515 5779 13521
rect 5721 13512 5733 13515
rect 5684 13484 5733 13512
rect 5684 13472 5690 13484
rect 5721 13481 5733 13484
rect 5767 13481 5779 13515
rect 9490 13512 9496 13524
rect 9451 13484 9496 13512
rect 5721 13475 5779 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 11422 13512 11428 13524
rect 9692 13484 11428 13512
rect 5534 13444 5540 13456
rect 4356 13416 5540 13444
rect 4249 13407 4307 13413
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 8754 13444 8760 13456
rect 8667 13416 8760 13444
rect 8754 13404 8760 13416
rect 8812 13444 8818 13456
rect 9033 13447 9091 13453
rect 9033 13444 9045 13447
rect 8812 13416 9045 13444
rect 8812 13404 8818 13416
rect 9033 13413 9045 13416
rect 9079 13413 9091 13447
rect 9033 13407 9091 13413
rect 5718 13376 5724 13388
rect 5679 13348 5724 13376
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 6086 13376 6092 13388
rect 6047 13348 6092 13376
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6454 13336 6460 13388
rect 6512 13336 6518 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 8662 13376 8668 13388
rect 8619 13348 8668 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 8662 13336 8668 13348
rect 8720 13376 8726 13388
rect 9692 13376 9720 13484
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13538 13512 13544 13524
rect 12943 13484 13544 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 14323 13515 14381 13521
rect 14323 13481 14335 13515
rect 14369 13512 14381 13515
rect 16574 13512 16580 13524
rect 14369 13484 16580 13512
rect 14369 13481 14381 13484
rect 14323 13475 14381 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 18288 13484 18613 13512
rect 18288 13472 18294 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 18601 13475 18659 13481
rect 9950 13444 9956 13456
rect 9911 13416 9956 13444
rect 9950 13404 9956 13416
rect 10008 13444 10014 13456
rect 12298 13447 12356 13453
rect 12298 13444 12310 13447
rect 10008 13416 12310 13444
rect 10008 13404 10014 13416
rect 12298 13413 12310 13416
rect 12344 13444 12356 13447
rect 12710 13444 12716 13456
rect 12344 13416 12716 13444
rect 12344 13413 12356 13416
rect 12298 13407 12356 13413
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 13170 13444 13176 13456
rect 13131 13416 13176 13444
rect 13170 13404 13176 13416
rect 13228 13444 13234 13456
rect 14642 13444 14648 13456
rect 13228 13416 14648 13444
rect 13228 13404 13234 13416
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 15105 13447 15163 13453
rect 15105 13413 15117 13447
rect 15151 13444 15163 13447
rect 15194 13444 15200 13456
rect 15151 13416 15200 13444
rect 15151 13413 15163 13416
rect 15105 13407 15163 13413
rect 15194 13404 15200 13416
rect 15252 13444 15258 13456
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 15252 13416 15485 13444
rect 15252 13404 15258 13416
rect 15473 13413 15485 13416
rect 15519 13413 15531 13447
rect 15473 13407 15531 13413
rect 17399 13447 17457 13453
rect 17399 13413 17411 13447
rect 17445 13444 17457 13447
rect 17678 13444 17684 13456
rect 17445 13416 17684 13444
rect 17445 13413 17457 13416
rect 17399 13407 17457 13413
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 18969 13447 19027 13453
rect 18969 13444 18981 13447
rect 18708 13416 18981 13444
rect 18708 13388 18736 13416
rect 18969 13413 18981 13416
rect 19015 13413 19027 13447
rect 18969 13407 19027 13413
rect 8720 13348 9720 13376
rect 8720 13336 8726 13348
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 14220 13379 14278 13385
rect 14220 13376 14232 13379
rect 14056 13348 14232 13376
rect 14056 13336 14062 13348
rect 14220 13345 14232 13348
rect 14266 13345 14278 13379
rect 14220 13339 14278 13345
rect 17957 13379 18015 13385
rect 17957 13345 17969 13379
rect 18003 13376 18015 13379
rect 18690 13376 18696 13388
rect 18003 13348 18696 13376
rect 18003 13345 18015 13348
rect 17957 13339 18015 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 4154 13308 4160 13320
rect 3573 13280 4160 13308
rect 4154 13268 4160 13280
rect 4212 13308 4218 13320
rect 4212 13280 4257 13308
rect 4212 13268 4218 13280
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4433 13311 4491 13317
rect 4433 13308 4445 13311
rect 4396 13280 4445 13308
rect 4396 13268 4402 13280
rect 4433 13277 4445 13280
rect 4479 13277 4491 13311
rect 6472 13308 6500 13336
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 4433 13271 4491 13277
rect 6104 13280 6653 13308
rect 6104 13240 6132 13280
rect 6641 13277 6653 13280
rect 6687 13308 6699 13311
rect 8018 13308 8024 13320
rect 6687 13280 8024 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 9674 13308 9680 13320
rect 9364 13280 9680 13308
rect 9364 13268 9370 13280
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11480 13280 11989 13308
rect 11480 13268 11486 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 15102 13268 15108 13320
rect 15160 13308 15166 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15160 13280 15393 13308
rect 15160 13268 15166 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 15381 13271 15439 13277
rect 16022 13268 16028 13280
rect 16080 13308 16086 13320
rect 16758 13308 16764 13320
rect 16080 13280 16764 13308
rect 16080 13268 16086 13280
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 17000 13280 17049 13308
rect 17000 13268 17006 13280
rect 17037 13277 17049 13280
rect 17083 13308 17095 13311
rect 17494 13308 17500 13320
rect 17083 13280 17500 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 18874 13308 18880 13320
rect 18835 13280 18880 13308
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19153 13311 19211 13317
rect 19153 13308 19165 13311
rect 19116 13280 19165 13308
rect 19116 13268 19122 13280
rect 19153 13277 19165 13280
rect 19199 13277 19211 13311
rect 19153 13271 19211 13277
rect 2240 13212 6132 13240
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 2240 13181 2268 13212
rect 6454 13200 6460 13252
rect 6512 13240 6518 13252
rect 7377 13243 7435 13249
rect 7377 13240 7389 13243
rect 6512 13212 7389 13240
rect 6512 13200 6518 13212
rect 7377 13209 7389 13212
rect 7423 13240 7435 13243
rect 7650 13240 7656 13252
rect 7423 13212 7656 13240
rect 7423 13209 7435 13212
rect 7377 13203 7435 13209
rect 7650 13200 7656 13212
rect 7708 13200 7714 13252
rect 9490 13200 9496 13252
rect 9548 13240 9554 13252
rect 10612 13240 10640 13268
rect 9548 13212 10640 13240
rect 9548 13200 9554 13212
rect 12066 13200 12072 13252
rect 12124 13240 12130 13252
rect 12124 13212 16344 13240
rect 12124 13200 12130 13212
rect 16316 13184 16344 13212
rect 2225 13175 2283 13181
rect 2225 13172 2237 13175
rect 1728 13144 2237 13172
rect 1728 13132 1734 13144
rect 2225 13141 2237 13144
rect 2271 13141 2283 13175
rect 3418 13172 3424 13184
rect 3379 13144 3424 13172
rect 2225 13135 2283 13141
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 5994 13172 6000 13184
rect 5408 13144 6000 13172
rect 5408 13132 5414 13144
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 6144 13144 7021 13172
rect 6144 13132 6150 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 7009 13135 7067 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10870 13172 10876 13184
rect 10831 13144 10876 13172
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 13538 13172 13544 13184
rect 13499 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 16942 13172 16948 13184
rect 16356 13144 16948 13172
rect 16356 13132 16362 13144
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 18230 13172 18236 13184
rect 18191 13144 18236 13172
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 1104 13082 20884 13104
rect 1104 13030 4648 13082
rect 4700 13030 4712 13082
rect 4764 13030 4776 13082
rect 4828 13030 4840 13082
rect 4892 13030 11982 13082
rect 12034 13030 12046 13082
rect 12098 13030 12110 13082
rect 12162 13030 12174 13082
rect 12226 13030 19315 13082
rect 19367 13030 19379 13082
rect 19431 13030 19443 13082
rect 19495 13030 19507 13082
rect 19559 13030 20884 13082
rect 1104 13008 20884 13030
rect 3970 12968 3976 12980
rect 3931 12940 3976 12968
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 4212 12940 4261 12968
rect 4212 12928 4218 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 4249 12931 4307 12937
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5810 12968 5816 12980
rect 5224 12940 5816 12968
rect 5224 12928 5230 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5951 12940 6009 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 5997 12937 6009 12940
rect 6043 12968 6055 12971
rect 8294 12968 8300 12980
rect 6043 12940 8300 12968
rect 6043 12937 6055 12940
rect 5997 12931 6055 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 9398 12968 9404 12980
rect 8812 12940 9404 12968
rect 8812 12928 8818 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10137 12971 10195 12977
rect 10137 12937 10149 12971
rect 10183 12968 10195 12971
rect 10870 12968 10876 12980
rect 10183 12940 10876 12968
rect 10183 12937 10195 12940
rect 10137 12931 10195 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 13906 12968 13912 12980
rect 13867 12940 13912 12968
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 15289 12971 15347 12977
rect 15289 12968 15301 12971
rect 15252 12940 15301 12968
rect 15252 12928 15258 12940
rect 15289 12937 15301 12940
rect 15335 12937 15347 12971
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 15289 12931 15347 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 18932 12940 19625 12968
rect 18932 12928 18938 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 19613 12931 19671 12937
rect 6638 12860 6644 12912
rect 6696 12900 6702 12912
rect 7098 12900 7104 12912
rect 6696 12872 7104 12900
rect 6696 12860 6702 12872
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 10781 12903 10839 12909
rect 10781 12900 10793 12903
rect 9732 12872 10793 12900
rect 9732 12860 9738 12872
rect 10781 12869 10793 12872
rect 10827 12869 10839 12903
rect 10781 12863 10839 12869
rect 11241 12903 11299 12909
rect 11241 12869 11253 12903
rect 11287 12900 11299 12903
rect 11422 12900 11428 12912
rect 11287 12872 11428 12900
rect 11287 12869 11299 12872
rect 11241 12863 11299 12869
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 13354 12900 13360 12912
rect 11664 12872 13360 12900
rect 11664 12860 11670 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2958 12832 2964 12844
rect 2639 12804 2964 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3418 12832 3424 12844
rect 3099 12804 3424 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 4396 12804 5181 12832
rect 4396 12792 4402 12804
rect 5169 12801 5181 12804
rect 5215 12832 5227 12835
rect 5350 12832 5356 12844
rect 5215 12804 5356 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5776 12804 6009 12832
rect 5776 12792 5782 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6788 12804 6929 12832
rect 6788 12792 6794 12804
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 8352 12804 8493 12832
rect 8352 12792 8358 12804
rect 8481 12801 8493 12804
rect 8527 12832 8539 12835
rect 9490 12832 9496 12844
rect 8527 12804 9496 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 12400 12804 12541 12832
rect 12400 12792 12406 12804
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 12802 12832 12808 12844
rect 12763 12804 12808 12832
rect 12529 12795 12587 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13228 12804 13461 12832
rect 13228 12792 13234 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13924 12832 13952 12928
rect 15841 12903 15899 12909
rect 15841 12869 15853 12903
rect 15887 12900 15899 12903
rect 16114 12900 16120 12912
rect 15887 12872 16120 12900
rect 15887 12869 15899 12872
rect 15841 12863 15899 12869
rect 16114 12860 16120 12872
rect 16172 12900 16178 12912
rect 16574 12900 16580 12912
rect 16172 12872 16580 12900
rect 16172 12860 16178 12872
rect 16574 12860 16580 12872
rect 16632 12860 16638 12912
rect 18598 12860 18604 12912
rect 18656 12900 18662 12912
rect 19981 12903 20039 12909
rect 19981 12900 19993 12903
rect 18656 12872 19993 12900
rect 18656 12860 18662 12872
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13924 12804 14381 12832
rect 13449 12795 13507 12801
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2038 12764 2044 12776
rect 1999 12736 2044 12764
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 9214 12764 9220 12776
rect 9175 12736 9220 12764
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 11400 12767 11458 12773
rect 11400 12733 11412 12767
rect 11446 12733 11458 12767
rect 11400 12727 11458 12733
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 3142 12696 3148 12708
rect 3007 12668 3148 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 3142 12656 3148 12668
rect 3200 12696 3206 12708
rect 3374 12699 3432 12705
rect 3374 12696 3386 12699
rect 3200 12668 3386 12696
rect 3200 12656 3206 12668
rect 3374 12665 3386 12668
rect 3420 12665 3432 12699
rect 4890 12696 4896 12708
rect 4851 12668 4896 12696
rect 3374 12659 3432 12665
rect 4890 12656 4896 12668
rect 4948 12656 4954 12708
rect 4985 12699 5043 12705
rect 4985 12665 4997 12699
rect 5031 12665 5043 12699
rect 4985 12659 5043 12665
rect 7009 12699 7067 12705
rect 7009 12665 7021 12699
rect 7055 12665 7067 12699
rect 7009 12659 7067 12665
rect 7561 12699 7619 12705
rect 7561 12665 7573 12699
rect 7607 12696 7619 12699
rect 7834 12696 7840 12708
rect 7607 12668 7840 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 1302 12588 1308 12640
rect 1360 12628 1366 12640
rect 1581 12631 1639 12637
rect 1581 12628 1593 12631
rect 1360 12600 1593 12628
rect 1360 12588 1366 12600
rect 1581 12597 1593 12600
rect 1627 12597 1639 12631
rect 1581 12591 1639 12597
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 4212 12600 4629 12628
rect 4212 12588 4218 12600
rect 4617 12597 4629 12600
rect 4663 12628 4675 12631
rect 5000 12628 5028 12659
rect 4663 12600 5028 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6270 12628 6276 12640
rect 6144 12600 6276 12628
rect 6144 12588 6150 12600
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12628 6702 12640
rect 7024 12628 7052 12659
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 9538 12699 9596 12705
rect 9538 12665 9550 12699
rect 9584 12665 9596 12699
rect 11415 12696 11443 12727
rect 11885 12699 11943 12705
rect 11885 12696 11897 12699
rect 11415 12668 11897 12696
rect 9538 12659 9596 12665
rect 11885 12665 11897 12668
rect 11931 12696 11943 12699
rect 11931 12668 12296 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 6696 12600 7052 12628
rect 8113 12631 8171 12637
rect 6696 12588 6702 12600
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8662 12628 8668 12640
rect 8159 12600 8668 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 9033 12631 9091 12637
rect 9033 12628 9045 12631
rect 8904 12600 9045 12628
rect 8904 12588 8910 12600
rect 9033 12597 9045 12600
rect 9079 12628 9091 12631
rect 9553 12628 9581 12659
rect 9950 12628 9956 12640
rect 9079 12600 9956 12628
rect 9079 12597 9091 12600
rect 9033 12591 9091 12597
rect 9950 12588 9956 12600
rect 10008 12628 10014 12640
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 10008 12600 10425 12628
rect 10008 12588 10014 12600
rect 10413 12597 10425 12600
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 11471 12631 11529 12637
rect 11471 12597 11483 12631
rect 11517 12628 11529 12631
rect 11606 12628 11612 12640
rect 11517 12600 11612 12628
rect 11517 12597 11529 12600
rect 11471 12591 11529 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 12158 12628 12164 12640
rect 12119 12600 12164 12628
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12268 12628 12296 12668
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 12676 12668 12721 12696
rect 12676 12656 12682 12668
rect 12710 12628 12716 12640
rect 12268 12600 12716 12628
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13464 12628 13492 12795
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 16850 12832 16856 12844
rect 16264 12804 16856 12832
rect 16264 12792 16270 12804
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17494 12832 17500 12844
rect 17368 12804 17500 12832
rect 17368 12792 17374 12804
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 18708 12841 18736 12872
rect 19981 12869 19993 12872
rect 20027 12869 20039 12903
rect 19981 12863 20039 12869
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12801 18751 12835
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18693 12795 18751 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 13872 12736 15577 12764
rect 13872 12724 13878 12736
rect 15565 12733 15577 12736
rect 15611 12764 15623 12767
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 15611 12736 16129 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 16117 12733 16129 12736
rect 16163 12733 16175 12767
rect 16574 12764 16580 12776
rect 16535 12736 16580 12764
rect 16117 12727 16175 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 13998 12696 14004 12708
rect 13786 12668 14004 12696
rect 13786 12628 13814 12668
rect 13998 12656 14004 12668
rect 14056 12656 14062 12708
rect 14690 12699 14748 12705
rect 14690 12696 14702 12699
rect 14200 12668 14702 12696
rect 13464 12600 13814 12628
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 14200 12637 14228 12668
rect 14690 12665 14702 12668
rect 14736 12696 14748 12699
rect 16850 12696 16856 12708
rect 14736 12668 16068 12696
rect 16811 12668 16856 12696
rect 14736 12665 14748 12668
rect 14690 12659 14748 12665
rect 14185 12631 14243 12637
rect 14185 12628 14197 12631
rect 14148 12600 14197 12628
rect 14148 12588 14154 12600
rect 14185 12597 14197 12600
rect 14231 12597 14243 12631
rect 14185 12591 14243 12597
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 15841 12631 15899 12637
rect 15841 12628 15853 12631
rect 15436 12600 15853 12628
rect 15436 12588 15442 12600
rect 15841 12597 15853 12600
rect 15887 12628 15899 12631
rect 15933 12631 15991 12637
rect 15933 12628 15945 12631
rect 15887 12600 15945 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 15933 12597 15945 12600
rect 15979 12597 15991 12631
rect 16040 12628 16068 12668
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 18785 12699 18843 12705
rect 18785 12665 18797 12699
rect 18831 12665 18843 12699
rect 18785 12659 18843 12665
rect 17129 12631 17187 12637
rect 17129 12628 17141 12631
rect 16040 12600 17141 12628
rect 15933 12591 15991 12597
rect 17129 12597 17141 12600
rect 17175 12628 17187 12631
rect 17310 12628 17316 12640
rect 17175 12600 17316 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 18509 12631 18567 12637
rect 18509 12628 18521 12631
rect 18104 12600 18521 12628
rect 18104 12588 18110 12600
rect 18509 12597 18521 12600
rect 18555 12628 18567 12631
rect 18800 12628 18828 12659
rect 18555 12600 18828 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 1104 12538 20884 12560
rect 1104 12486 8315 12538
rect 8367 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 15648 12538
rect 15700 12486 15712 12538
rect 15764 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 20884 12538
rect 1104 12464 20884 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 2225 12427 2283 12433
rect 2225 12424 2237 12427
rect 1820 12396 2237 12424
rect 1820 12384 1826 12396
rect 2225 12393 2237 12396
rect 2271 12393 2283 12427
rect 2225 12387 2283 12393
rect 1949 12359 2007 12365
rect 1949 12325 1961 12359
rect 1995 12356 2007 12359
rect 2038 12356 2044 12368
rect 1995 12328 2044 12356
rect 1995 12325 2007 12328
rect 1949 12319 2007 12325
rect 2038 12316 2044 12328
rect 2096 12316 2102 12368
rect 1464 12291 1522 12297
rect 1464 12257 1476 12291
rect 1510 12288 1522 12291
rect 1578 12288 1584 12300
rect 1510 12260 1584 12288
rect 1510 12257 1522 12260
rect 1464 12251 1522 12257
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 2056 12220 2084 12316
rect 2240 12288 2268 12387
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3384 12396 3801 12424
rect 3384 12384 3390 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 3789 12387 3847 12393
rect 4126 12396 4445 12424
rect 3145 12359 3203 12365
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 3418 12356 3424 12368
rect 3191 12328 3424 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 2240 12260 2421 12288
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2958 12288 2964 12300
rect 2919 12260 2964 12288
rect 2409 12251 2467 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 3804 12288 3832 12387
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 4126 12356 4154 12396
rect 4433 12393 4445 12396
rect 4479 12393 4491 12427
rect 4433 12387 4491 12393
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 5629 12427 5687 12433
rect 5629 12424 5641 12427
rect 5500 12396 5641 12424
rect 5500 12384 5506 12396
rect 5629 12393 5641 12396
rect 5675 12393 5687 12427
rect 5629 12387 5687 12393
rect 4028 12328 4154 12356
rect 4028 12316 4034 12328
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3804 12260 4077 12288
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 5644 12288 5672 12387
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 6144 12396 6193 12424
rect 6144 12384 6150 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 6181 12387 6239 12393
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 6696 12396 6745 12424
rect 6696 12384 6702 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 6733 12387 6791 12393
rect 10410 12384 10416 12436
rect 10468 12424 10474 12436
rect 11238 12424 11244 12436
rect 10468 12396 11244 12424
rect 10468 12384 10474 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12400 12396 12909 12424
rect 12400 12384 12406 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 14274 12424 14280 12436
rect 14235 12396 14280 12424
rect 12897 12387 12955 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 15102 12424 15108 12436
rect 15063 12396 15108 12424
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 17092 12396 17141 12424
rect 17092 12384 17098 12396
rect 17129 12393 17141 12396
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 9214 12356 9220 12368
rect 8803 12328 9220 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 9306 12316 9312 12368
rect 9364 12356 9370 12368
rect 9953 12359 10011 12365
rect 9953 12356 9965 12359
rect 9364 12328 9965 12356
rect 9364 12316 9370 12328
rect 9953 12325 9965 12328
rect 9999 12356 10011 12359
rect 10594 12356 10600 12368
rect 9999 12328 10600 12356
rect 9999 12325 10011 12328
rect 9953 12319 10011 12325
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 11695 12359 11753 12365
rect 11695 12325 11707 12359
rect 11741 12325 11753 12359
rect 13722 12356 13728 12368
rect 11695 12319 11753 12325
rect 13188 12328 13728 12356
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5644 12260 5825 12288
rect 4065 12251 4123 12257
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6788 12260 7021 12288
rect 6788 12248 6794 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 7009 12251 7067 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8570 12288 8576 12300
rect 8531 12260 8576 12288
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 10502 12248 10508 12300
rect 10560 12288 10566 12300
rect 11710 12288 11738 12319
rect 12158 12288 12164 12300
rect 10560 12260 10605 12288
rect 11710 12260 12164 12288
rect 10560 12248 10566 12260
rect 12158 12248 12164 12260
rect 12216 12288 12222 12300
rect 12342 12288 12348 12300
rect 12216 12260 12348 12288
rect 12216 12248 12222 12260
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 13188 12297 13216 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 15068 12328 15485 12356
rect 15068 12316 15074 12328
rect 15473 12325 15485 12328
rect 15519 12325 15531 12359
rect 15473 12319 15531 12325
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12257 13231 12291
rect 13173 12251 13231 12257
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 13320 12260 13645 12288
rect 13320 12248 13326 12260
rect 13633 12257 13645 12260
rect 13679 12257 13691 12291
rect 17144 12288 17172 12387
rect 17310 12384 17316 12436
rect 17368 12424 17374 12436
rect 18233 12427 18291 12433
rect 17368 12396 17493 12424
rect 17368 12384 17374 12396
rect 17465 12356 17493 12396
rect 18233 12393 18245 12427
rect 18279 12424 18291 12427
rect 19150 12424 19156 12436
rect 18279 12396 19156 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 19150 12384 19156 12396
rect 19208 12424 19214 12436
rect 19208 12396 19288 12424
rect 19208 12384 19214 12396
rect 17678 12365 17684 12368
rect 17635 12359 17684 12365
rect 17635 12356 17647 12359
rect 17465 12328 17647 12356
rect 17635 12325 17647 12328
rect 17681 12325 17684 12359
rect 17635 12319 17684 12325
rect 17678 12316 17684 12319
rect 17736 12356 17742 12368
rect 17736 12328 17783 12356
rect 17736 12316 17742 12328
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19260 12365 19288 12396
rect 18785 12359 18843 12365
rect 18785 12356 18797 12359
rect 18748 12328 18797 12356
rect 18748 12316 18754 12328
rect 18785 12325 18797 12328
rect 18831 12325 18843 12359
rect 18785 12319 18843 12325
rect 19245 12359 19303 12365
rect 19245 12325 19257 12359
rect 19291 12325 19303 12359
rect 19245 12319 19303 12325
rect 17313 12291 17371 12297
rect 17313 12288 17325 12291
rect 17144 12260 17325 12288
rect 13633 12251 13691 12257
rect 17313 12257 17325 12260
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 2774 12220 2780 12232
rect 2056 12192 2780 12220
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 1535 12155 1593 12161
rect 1535 12121 1547 12155
rect 1581 12152 1593 12155
rect 4522 12152 4528 12164
rect 1581 12124 4528 12152
rect 1581 12121 1593 12124
rect 1535 12115 1593 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 4890 12112 4896 12164
rect 4948 12152 4954 12164
rect 9876 12152 9904 12183
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11296 12192 11345 12220
rect 11296 12180 11302 12192
rect 11333 12189 11345 12192
rect 11379 12220 11391 12223
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 11379 12192 13553 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14700 12192 15393 12220
rect 14700 12180 14706 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 16022 12220 16028 12232
rect 15983 12192 16028 12220
rect 15381 12183 15439 12189
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 18966 12180 18972 12232
rect 19024 12220 19030 12232
rect 19153 12223 19211 12229
rect 19153 12220 19165 12223
rect 19024 12192 19165 12220
rect 19024 12180 19030 12192
rect 19153 12189 19165 12192
rect 19199 12189 19211 12223
rect 19153 12183 19211 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 10502 12152 10508 12164
rect 4948 12124 5212 12152
rect 9876 12124 10508 12152
rect 4948 12112 4954 12124
rect 5184 12096 5212 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 19058 12112 19064 12164
rect 19116 12152 19122 12164
rect 19444 12152 19472 12183
rect 19116 12124 19472 12152
rect 19116 12112 19122 12124
rect 3418 12084 3424 12096
rect 3379 12056 3424 12084
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 4982 12084 4988 12096
rect 4943 12056 4988 12084
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5261 12087 5319 12093
rect 5261 12084 5273 12087
rect 5224 12056 5273 12084
rect 5224 12044 5230 12056
rect 5261 12053 5273 12056
rect 5307 12053 5319 12087
rect 5261 12047 5319 12053
rect 12253 12087 12311 12093
rect 12253 12053 12265 12087
rect 12299 12084 12311 12087
rect 12618 12084 12624 12096
rect 12299 12056 12624 12084
rect 12299 12053 12311 12056
rect 12253 12047 12311 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 1104 11994 20884 12016
rect 1104 11942 4648 11994
rect 4700 11942 4712 11994
rect 4764 11942 4776 11994
rect 4828 11942 4840 11994
rect 4892 11942 11982 11994
rect 12034 11942 12046 11994
rect 12098 11942 12110 11994
rect 12162 11942 12174 11994
rect 12226 11942 19315 11994
rect 19367 11942 19379 11994
rect 19431 11942 19443 11994
rect 19495 11942 19507 11994
rect 19559 11942 20884 11994
rect 1104 11920 20884 11942
rect 3142 11880 3148 11892
rect 3103 11852 3148 11880
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4893 11883 4951 11889
rect 4212 11852 4257 11880
rect 4212 11840 4218 11852
rect 4893 11849 4905 11883
rect 4939 11880 4951 11883
rect 4982 11880 4988 11892
rect 4939 11852 4988 11880
rect 4939 11849 4951 11852
rect 4893 11843 4951 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8076 11852 8861 11880
rect 8076 11840 8082 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 8849 11843 8907 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 11238 11880 11244 11892
rect 11199 11852 11244 11880
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13320 11852 13461 11880
rect 13320 11840 13326 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 17310 11880 17316 11892
rect 17271 11852 17316 11880
rect 13449 11843 13507 11849
rect 17310 11840 17316 11852
rect 17368 11880 17374 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17368 11852 17785 11880
rect 17368 11840 17374 11852
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 17773 11843 17831 11849
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 19245 11883 19303 11889
rect 19245 11880 19257 11883
rect 19208 11852 19257 11880
rect 19208 11840 19214 11852
rect 19245 11849 19257 11852
rect 19291 11849 19303 11883
rect 19245 11843 19303 11849
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 4525 11815 4583 11821
rect 4525 11812 4537 11815
rect 4028 11784 4537 11812
rect 4028 11772 4034 11784
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 2455 11716 3249 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 3237 11713 3249 11716
rect 3283 11744 3295 11747
rect 3418 11744 3424 11756
rect 3283 11716 3424 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 1946 11676 1952 11688
rect 1907 11648 1952 11676
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2271 11648 2360 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2332 11552 2360 11648
rect 3142 11568 3148 11620
rect 3200 11608 3206 11620
rect 3558 11611 3616 11617
rect 3558 11608 3570 11611
rect 3200 11580 3570 11608
rect 3200 11568 3206 11580
rect 3558 11577 3570 11580
rect 3604 11608 3616 11611
rect 4126 11608 4154 11784
rect 4525 11781 4537 11784
rect 4571 11812 4583 11815
rect 6086 11812 6092 11824
rect 4571 11784 6092 11812
rect 4571 11781 4583 11784
rect 4525 11775 4583 11781
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 16298 11772 16304 11824
rect 16356 11812 16362 11824
rect 18598 11812 18604 11824
rect 16356 11784 18604 11812
rect 16356 11772 16362 11784
rect 18598 11772 18604 11784
rect 18656 11772 18662 11824
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 5074 11744 5080 11756
rect 4396 11716 5080 11744
rect 4396 11704 4402 11716
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5350 11744 5356 11756
rect 5311 11716 5356 11744
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 6914 11744 6920 11756
rect 6875 11716 6920 11744
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11744 9919 11747
rect 10042 11744 10048 11756
rect 9907 11716 10048 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10594 11704 10600 11756
rect 10652 11744 10658 11756
rect 10873 11747 10931 11753
rect 10652 11716 10732 11744
rect 10652 11704 10658 11716
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8570 11676 8576 11688
rect 8159 11648 8576 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8570 11636 8576 11648
rect 8628 11676 8634 11688
rect 9306 11676 9312 11688
rect 8628 11648 9312 11676
rect 8628 11636 8634 11648
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 10704 11676 10732 11716
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 11606 11744 11612 11756
rect 10919 11716 11612 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 11606 11704 11612 11716
rect 11664 11744 11670 11756
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 11664 11716 12541 11744
rect 11664 11704 11670 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14274 11744 14280 11756
rect 14231 11716 14280 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 16942 11744 16948 11756
rect 15703 11716 16948 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 11146 11676 11152 11688
rect 10704 11648 11152 11676
rect 11146 11636 11152 11648
rect 11204 11676 11210 11688
rect 16408 11685 16436 11716
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11744 18107 11747
rect 18138 11744 18144 11756
rect 18095 11716 18144 11744
rect 18095 11713 18107 11716
rect 18049 11707 18107 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 11368 11679 11426 11685
rect 11368 11676 11380 11679
rect 11204 11648 11380 11676
rect 11204 11636 11210 11648
rect 11368 11645 11380 11648
rect 11414 11676 11426 11679
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11414 11648 11805 11676
rect 11414 11645 11426 11648
rect 11368 11639 11426 11645
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16577 11679 16635 11685
rect 16577 11645 16589 11679
rect 16623 11645 16635 11679
rect 16577 11639 16635 11645
rect 5074 11608 5080 11620
rect 3604 11580 4154 11608
rect 5035 11580 5080 11608
rect 3604 11577 3616 11580
rect 3558 11571 3616 11577
rect 5074 11568 5080 11580
rect 5132 11568 5138 11620
rect 5169 11611 5227 11617
rect 5169 11577 5181 11611
rect 5215 11577 5227 11611
rect 5169 11571 5227 11577
rect 7009 11611 7067 11617
rect 7009 11577 7021 11611
rect 7055 11577 7067 11611
rect 7558 11608 7564 11620
rect 7519 11580 7564 11608
rect 7009 11571 7067 11577
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2685 11543 2743 11549
rect 2685 11540 2697 11543
rect 2372 11512 2697 11540
rect 2372 11500 2378 11512
rect 2685 11509 2697 11512
rect 2731 11540 2743 11543
rect 2958 11540 2964 11552
rect 2731 11512 2964 11540
rect 2731 11509 2743 11512
rect 2685 11503 2743 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 4982 11500 4988 11552
rect 5040 11540 5046 11552
rect 5184 11540 5212 11571
rect 6086 11540 6092 11552
rect 5040 11512 5212 11540
rect 6047 11512 6092 11540
rect 5040 11500 5046 11512
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7024 11540 7052 11571
rect 7558 11568 7564 11580
rect 7616 11568 7622 11620
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 9858 11608 9864 11620
rect 9723 11580 9864 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 9858 11568 9864 11580
rect 9916 11608 9922 11620
rect 9953 11611 10011 11617
rect 9953 11608 9965 11611
rect 9916 11580 9965 11608
rect 9916 11568 9922 11580
rect 9953 11577 9965 11580
rect 9999 11577 10011 11611
rect 10502 11608 10508 11620
rect 10415 11580 10508 11608
rect 9953 11571 10011 11577
rect 10502 11568 10508 11580
rect 10560 11608 10566 11620
rect 10560 11580 12296 11608
rect 10560 11568 10566 11580
rect 6696 11512 7052 11540
rect 6696 11500 6702 11512
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8168 11512 8401 11540
rect 8168 11500 8174 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 11471 11543 11529 11549
rect 11471 11509 11483 11543
rect 11517 11540 11529 11543
rect 11606 11540 11612 11552
rect 11517 11512 11612 11540
rect 11517 11509 11529 11512
rect 11471 11503 11529 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12268 11540 12296 11580
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 13173 11611 13231 11617
rect 12676 11580 12721 11608
rect 12676 11568 12682 11580
rect 13173 11577 13185 11611
rect 13219 11608 13231 11611
rect 13262 11608 13268 11620
rect 13219 11580 13268 11608
rect 13219 11577 13231 11580
rect 13173 11571 13231 11577
rect 13188 11540 13216 11571
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 14506 11611 14564 11617
rect 14506 11577 14518 11611
rect 14552 11577 14564 11611
rect 14506 11571 14564 11577
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16298 11608 16304 11620
rect 16071 11580 16304 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 14090 11540 14096 11552
rect 12268 11512 13216 11540
rect 14051 11512 14096 11540
rect 14090 11500 14096 11512
rect 14148 11540 14154 11552
rect 14521 11540 14549 11571
rect 16298 11568 16304 11580
rect 16356 11608 16362 11620
rect 16592 11608 16620 11639
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 18966 11676 18972 11688
rect 17092 11648 18972 11676
rect 17092 11636 17098 11648
rect 18966 11636 18972 11648
rect 19024 11676 19030 11688
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19024 11648 19625 11676
rect 19024 11636 19030 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 16356 11580 16620 11608
rect 16356 11568 16362 11580
rect 16758 11568 16764 11620
rect 16816 11608 16822 11620
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 16816 11580 16865 11608
rect 16816 11568 16822 11580
rect 16853 11577 16865 11580
rect 16899 11577 16911 11611
rect 16853 11571 16911 11577
rect 17310 11568 17316 11620
rect 17368 11608 17374 11620
rect 18370 11611 18428 11617
rect 18370 11608 18382 11611
rect 17368 11580 18382 11608
rect 17368 11568 17374 11580
rect 18370 11577 18382 11580
rect 18416 11577 18428 11611
rect 18370 11571 18428 11577
rect 15102 11540 15108 11552
rect 14148 11512 14549 11540
rect 15063 11512 15108 11540
rect 14148 11500 14154 11512
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 18969 11543 19027 11549
rect 18969 11509 18981 11543
rect 19015 11540 19027 11543
rect 19058 11540 19064 11552
rect 19015 11512 19064 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 19058 11500 19064 11512
rect 19116 11500 19122 11552
rect 1104 11450 20884 11472
rect 1104 11398 8315 11450
rect 8367 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 15648 11450
rect 15700 11398 15712 11450
rect 15764 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 20884 11450
rect 1104 11376 20884 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11336 1642 11348
rect 2038 11336 2044 11348
rect 1636 11308 2044 11336
rect 1636 11296 1642 11308
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2406 11336 2412 11348
rect 2367 11308 2412 11336
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 6454 11336 6460 11348
rect 3568 11308 6460 11336
rect 3568 11296 3574 11308
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6880 11308 6929 11336
rect 6880 11296 6886 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 10042 11336 10048 11348
rect 9999 11308 10048 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 12158 11336 12164 11348
rect 11204 11308 12164 11336
rect 11204 11296 11210 11308
rect 1946 11228 1952 11280
rect 2004 11268 2010 11280
rect 3528 11268 3556 11296
rect 2004 11240 3556 11268
rect 2004 11228 2010 11240
rect 2608 11209 2636 11240
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4249 11271 4307 11277
rect 4249 11268 4261 11271
rect 4028 11240 4261 11268
rect 4028 11228 4034 11240
rect 4249 11237 4261 11240
rect 4295 11237 4307 11271
rect 4249 11231 4307 11237
rect 5970 11271 6028 11277
rect 5970 11237 5982 11271
rect 6016 11268 6028 11271
rect 6086 11268 6092 11280
rect 6016 11240 6092 11268
rect 6016 11237 6028 11240
rect 5970 11231 6028 11237
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 6696 11240 7665 11268
rect 6696 11228 6702 11240
rect 7653 11237 7665 11240
rect 7699 11237 7711 11271
rect 7653 11231 7711 11237
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11268 9551 11271
rect 10502 11268 10508 11280
rect 9539 11240 10508 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 11238 11268 11244 11280
rect 10836 11240 11244 11268
rect 10836 11228 10842 11240
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 11485 11277 11513 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12618 11336 12624 11348
rect 12575 11308 12624 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 13780 11308 13921 11336
rect 13780 11296 13786 11308
rect 13909 11305 13921 11308
rect 13955 11305 13967 11339
rect 13909 11299 13967 11305
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 14240 11308 14289 11336
rect 14240 11296 14246 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 15010 11336 15016 11348
rect 14971 11308 15016 11336
rect 14277 11299 14335 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 18196 11308 18337 11336
rect 18196 11296 18202 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 18506 11296 18512 11348
rect 18564 11336 18570 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 18564 11308 18705 11336
rect 18564 11296 18570 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 18693 11299 18751 11305
rect 11470 11271 11528 11277
rect 11470 11237 11482 11271
rect 11516 11237 11528 11271
rect 11470 11231 11528 11237
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 13081 11271 13139 11277
rect 13081 11268 13093 11271
rect 12400 11240 13093 11268
rect 12400 11228 12406 11240
rect 13081 11237 13093 11240
rect 13127 11237 13139 11271
rect 13081 11231 13139 11237
rect 15102 11228 15108 11280
rect 15160 11268 15166 11280
rect 15473 11271 15531 11277
rect 15473 11268 15485 11271
rect 15160 11240 15485 11268
rect 15160 11228 15166 11240
rect 15473 11237 15485 11240
rect 15519 11237 15531 11271
rect 16022 11268 16028 11280
rect 15983 11240 16028 11268
rect 15473 11231 15531 11237
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 17310 11228 17316 11280
rect 17368 11268 17374 11280
rect 17450 11271 17508 11277
rect 17450 11268 17462 11271
rect 17368 11240 17462 11268
rect 17368 11228 17374 11240
rect 17450 11237 17462 11240
rect 17496 11237 17508 11271
rect 19058 11268 19064 11280
rect 19019 11240 19064 11268
rect 17450 11231 17508 11237
rect 19058 11228 19064 11240
rect 19116 11228 19122 11280
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11169 2651 11203
rect 2774 11200 2780 11212
rect 2735 11172 2780 11200
rect 2593 11163 2651 11169
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6972 11172 7297 11200
rect 6972 11160 6978 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 10042 11200 10048 11212
rect 9272 11172 10048 11200
rect 9272 11160 9278 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11330 11200 11336 11212
rect 11195 11172 11336 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17862 11200 17868 11212
rect 17175 11172 17868 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 4154 11132 4160 11144
rect 2924 11104 4160 11132
rect 2924 11092 2930 11104
rect 4154 11092 4160 11104
rect 4212 11132 4218 11144
rect 4801 11135 4859 11141
rect 4212 11104 4257 11132
rect 4212 11092 4218 11104
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 5718 11132 5724 11144
rect 5679 11104 5724 11132
rect 4801 11095 4859 11101
rect 2222 11024 2228 11076
rect 2280 11064 2286 11076
rect 3602 11064 3608 11076
rect 2280 11036 3608 11064
rect 2280 11024 2286 11036
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 4816 11064 4844 11095
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7432 11104 7573 11132
rect 7432 11092 7438 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7834 11132 7840 11144
rect 7795 11104 7840 11132
rect 7561 11095 7619 11101
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 8076 11104 10701 11132
rect 8076 11092 8082 11104
rect 10689 11101 10701 11104
rect 10735 11132 10747 11135
rect 10778 11132 10784 11144
rect 10735 11104 10784 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 12710 11132 12716 11144
rect 11756 11104 12716 11132
rect 11756 11092 11762 11104
rect 12710 11092 12716 11104
rect 12768 11132 12774 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12768 11104 13001 11132
rect 12768 11092 12774 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 12989 11095 13047 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 15252 11104 15393 11132
rect 15252 11092 15258 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17310 11132 17316 11144
rect 17000 11104 17316 11132
rect 17000 11092 17006 11104
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 18969 11135 19027 11141
rect 18969 11101 18981 11135
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 5074 11064 5080 11076
rect 4816 11036 5080 11064
rect 5074 11024 5080 11036
rect 5132 11064 5138 11076
rect 5169 11067 5227 11073
rect 5169 11064 5181 11067
rect 5132 11036 5181 11064
rect 5132 11024 5138 11036
rect 5169 11033 5181 11036
rect 5215 11064 5227 11067
rect 7852 11064 7880 11092
rect 12894 11064 12900 11076
rect 5215 11036 7880 11064
rect 11716 11036 12900 11064
rect 5215 11033 5227 11036
rect 5169 11027 5227 11033
rect 11716 11008 11744 11036
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 18874 11024 18880 11076
rect 18932 11064 18938 11076
rect 18984 11064 19012 11095
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 19208 11104 19257 11132
rect 19208 11092 19214 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 18932 11036 19012 11064
rect 18932 11024 18938 11036
rect 2041 10999 2099 11005
rect 2041 10965 2053 10999
rect 2087 10996 2099 10999
rect 2314 10996 2320 11008
rect 2087 10968 2320 10996
rect 2087 10965 2099 10968
rect 2041 10959 2099 10965
rect 2314 10956 2320 10968
rect 2372 10956 2378 11008
rect 3421 10999 3479 11005
rect 3421 10965 3433 10999
rect 3467 10996 3479 10999
rect 3510 10996 3516 11008
rect 3467 10968 3516 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3694 10996 3700 11008
rect 3655 10968 3700 10996
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 5442 10996 5448 11008
rect 5403 10968 5448 10996
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 6638 10996 6644 11008
rect 6599 10968 6644 10996
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 10275 10999 10333 11005
rect 10275 10965 10287 10999
rect 10321 10996 10333 10999
rect 10594 10996 10600 11008
rect 10321 10968 10600 10996
rect 10321 10965 10333 10968
rect 10275 10959 10333 10965
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 11698 10956 11704 11008
rect 11756 10956 11762 11008
rect 12069 10999 12127 11005
rect 12069 10965 12081 10999
rect 12115 10996 12127 10999
rect 12342 10996 12348 11008
rect 12115 10968 12348 10996
rect 12115 10965 12127 10968
rect 12069 10959 12127 10965
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 14642 10996 14648 11008
rect 14603 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 1104 10906 20884 10928
rect 1104 10854 4648 10906
rect 4700 10854 4712 10906
rect 4764 10854 4776 10906
rect 4828 10854 4840 10906
rect 4892 10854 11982 10906
rect 12034 10854 12046 10906
rect 12098 10854 12110 10906
rect 12162 10854 12174 10906
rect 12226 10854 19315 10906
rect 19367 10854 19379 10906
rect 19431 10854 19443 10906
rect 19495 10854 19507 10906
rect 19559 10854 20884 10906
rect 1104 10832 20884 10854
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10792 2651 10795
rect 2774 10792 2780 10804
rect 2639 10764 2780 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 2961 10795 3019 10801
rect 2961 10761 2973 10795
rect 3007 10792 3019 10795
rect 3142 10792 3148 10804
rect 3007 10764 3148 10792
rect 3007 10761 3019 10764
rect 2961 10755 3019 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4212 10764 4629 10792
rect 4212 10752 4218 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 4617 10755 4675 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 8110 10792 8116 10804
rect 6748 10764 8116 10792
rect 1946 10684 1952 10736
rect 2004 10724 2010 10736
rect 3878 10724 3884 10736
rect 2004 10696 3884 10724
rect 2004 10684 2010 10696
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 5902 10724 5908 10736
rect 5859 10696 5908 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3142 10656 3148 10668
rect 3099 10628 3148 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3694 10656 3700 10668
rect 3200 10628 3700 10656
rect 3200 10616 3206 10628
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 5123 10628 5273 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5261 10625 5273 10628
rect 5307 10656 5319 10659
rect 6748 10656 6776 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9858 10792 9864 10804
rect 9819 10764 9864 10792
rect 9858 10752 9864 10764
rect 9916 10792 9922 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 9916 10764 10517 10792
rect 9916 10752 9922 10764
rect 10505 10761 10517 10764
rect 10551 10792 10563 10795
rect 10870 10792 10876 10804
rect 10551 10764 10876 10792
rect 10551 10761 10563 10764
rect 10505 10755 10563 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12802 10752 12808 10804
rect 12860 10752 12866 10804
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 15381 10795 15439 10801
rect 15381 10792 15393 10795
rect 15160 10764 15393 10792
rect 15160 10752 15166 10764
rect 15381 10761 15393 10764
rect 15427 10761 15439 10795
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 15381 10755 15439 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 18104 10764 18337 10792
rect 18104 10752 18110 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 6822 10684 6828 10736
rect 6880 10724 6886 10736
rect 6880 10696 6960 10724
rect 6880 10684 6886 10696
rect 6932 10665 6960 10696
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7432 10696 8217 10724
rect 7432 10684 7438 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 11333 10727 11391 10733
rect 11333 10693 11345 10727
rect 11379 10724 11391 10727
rect 12820 10724 12848 10752
rect 13081 10727 13139 10733
rect 13081 10724 13093 10727
rect 11379 10696 13093 10724
rect 11379 10693 11391 10696
rect 11333 10687 11391 10693
rect 13081 10693 13093 10696
rect 13127 10693 13139 10727
rect 17034 10724 17040 10736
rect 16995 10696 17040 10724
rect 13081 10687 13139 10693
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 5307 10628 6776 10656
rect 6917 10659 6975 10665
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 6917 10619 6975 10625
rect 7282 10616 7288 10628
rect 7340 10656 7346 10668
rect 7558 10656 7564 10668
rect 7340 10628 7564 10656
rect 7340 10616 7346 10628
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8938 10656 8944 10668
rect 8899 10628 8944 10656
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 10778 10656 10784 10668
rect 10739 10628 10784 10656
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 11940 10628 12541 10656
rect 11940 10616 11946 10628
rect 12529 10625 12541 10628
rect 12575 10656 12587 10659
rect 12802 10656 12808 10668
rect 12575 10628 12808 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 14182 10656 14188 10668
rect 14143 10628 14188 10656
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16574 10656 16580 10668
rect 16531 10628 16580 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16574 10616 16580 10628
rect 16632 10656 16638 10668
rect 17218 10656 17224 10668
rect 16632 10628 17224 10656
rect 16632 10616 16638 10628
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2314 10588 2320 10600
rect 2087 10560 2320 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 6086 10548 6092 10600
rect 6144 10588 6150 10600
rect 6273 10591 6331 10597
rect 6273 10588 6285 10591
rect 6144 10560 6285 10588
rect 6144 10548 6150 10560
rect 6273 10557 6285 10560
rect 6319 10588 6331 10591
rect 6730 10588 6736 10600
rect 6319 10560 6736 10588
rect 6319 10557 6331 10560
rect 6273 10551 6331 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 15068 10560 15117 10588
rect 15068 10548 15074 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 2222 10520 2228 10532
rect 2183 10492 2228 10520
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 3374 10523 3432 10529
rect 3374 10520 3386 10523
rect 3292 10492 3386 10520
rect 3292 10480 3298 10492
rect 3374 10489 3386 10492
rect 3420 10489 3432 10523
rect 3374 10483 3432 10489
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5408 10492 5453 10520
rect 5408 10480 5414 10492
rect 6638 10480 6644 10532
rect 6696 10520 6702 10532
rect 7009 10523 7067 10529
rect 7009 10520 7021 10523
rect 6696 10492 7021 10520
rect 6696 10480 6702 10492
rect 7009 10489 7021 10492
rect 7055 10489 7067 10523
rect 9262 10523 9320 10529
rect 9262 10520 9274 10523
rect 7009 10483 7067 10489
rect 8864 10492 9274 10520
rect 3970 10452 3976 10464
rect 3883 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10452 4034 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 4028 10424 4261 10452
rect 4028 10412 4034 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6822 10452 6828 10464
rect 6328 10424 6828 10452
rect 6328 10412 6334 10424
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7024 10452 7052 10483
rect 8864 10464 8892 10492
rect 9262 10489 9274 10492
rect 9308 10489 9320 10523
rect 9262 10483 9320 10489
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 12621 10523 12679 10529
rect 10928 10492 10973 10520
rect 10928 10480 10934 10492
rect 12621 10489 12633 10523
rect 12667 10489 12679 10523
rect 12621 10483 12679 10489
rect 14506 10523 14564 10529
rect 14506 10489 14518 10523
rect 14552 10489 14564 10523
rect 14506 10483 14564 10489
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 16577 10523 16635 10529
rect 16577 10520 16589 10523
rect 16347 10492 16589 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 16577 10489 16589 10492
rect 16623 10520 16635 10523
rect 16942 10520 16948 10532
rect 16623 10492 16948 10520
rect 16623 10489 16635 10492
rect 16577 10483 16635 10489
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7024 10424 7849 10452
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8846 10452 8852 10464
rect 8807 10424 8852 10452
rect 7837 10415 7895 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 10042 10452 10048 10464
rect 9732 10424 10048 10452
rect 9732 10412 9738 10424
rect 10042 10412 10048 10424
rect 10100 10452 10106 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 10100 10424 10149 10452
rect 10100 10412 10106 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 10137 10415 10195 10421
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11146 10452 11152 10464
rect 10560 10424 11152 10452
rect 10560 10412 10566 10424
rect 11146 10412 11152 10424
rect 11204 10452 11210 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11204 10424 11713 10452
rect 11204 10412 11210 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12636 10452 12664 10483
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 12400 10424 13461 10452
rect 12400 10412 12406 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 14090 10452 14096 10464
rect 14051 10424 14096 10452
rect 13449 10415 13507 10421
rect 14090 10412 14096 10424
rect 14148 10452 14154 10464
rect 14521 10452 14549 10483
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 18340 10520 18368 10755
rect 19058 10752 19064 10804
rect 19116 10792 19122 10804
rect 19521 10795 19579 10801
rect 19521 10792 19533 10795
rect 19116 10764 19533 10792
rect 19116 10752 19122 10764
rect 19521 10761 19533 10764
rect 19567 10761 19579 10795
rect 19521 10755 19579 10761
rect 18506 10684 18512 10736
rect 18564 10724 18570 10736
rect 18564 10696 18644 10724
rect 18564 10684 18570 10696
rect 18616 10665 18644 10696
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18874 10656 18880 10668
rect 18835 10628 18880 10656
rect 18601 10619 18659 10625
rect 18874 10616 18880 10628
rect 18932 10656 18938 10668
rect 19889 10659 19947 10665
rect 19889 10656 19901 10659
rect 18932 10628 19901 10656
rect 18932 10616 18938 10628
rect 19889 10625 19901 10628
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 18693 10523 18751 10529
rect 18693 10520 18705 10523
rect 18340 10492 18705 10520
rect 18693 10489 18705 10492
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 14148 10424 14549 10452
rect 14148 10412 14154 10424
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 15749 10455 15807 10461
rect 15749 10452 15761 10455
rect 15252 10424 15761 10452
rect 15252 10412 15258 10424
rect 15749 10421 15761 10424
rect 15795 10421 15807 10455
rect 15749 10415 15807 10421
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17368 10424 17417 10452
rect 17368 10412 17374 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 1104 10362 20884 10384
rect 1104 10310 8315 10362
rect 8367 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 15648 10362
rect 15700 10310 15712 10362
rect 15764 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 20884 10362
rect 1104 10288 20884 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1673 10251 1731 10257
rect 1673 10248 1685 10251
rect 1544 10220 1685 10248
rect 1544 10208 1550 10220
rect 1673 10217 1685 10220
rect 1719 10217 1731 10251
rect 1673 10211 1731 10217
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 5718 10248 5724 10260
rect 2280 10220 5724 10248
rect 2280 10208 2286 10220
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 7282 10248 7288 10260
rect 6288 10220 7288 10248
rect 1949 10183 2007 10189
rect 1949 10149 1961 10183
rect 1995 10180 2007 10183
rect 2314 10180 2320 10192
rect 1995 10152 2320 10180
rect 1995 10149 2007 10152
rect 1949 10143 2007 10149
rect 2314 10140 2320 10152
rect 2372 10180 2378 10192
rect 3142 10180 3148 10192
rect 2372 10152 3004 10180
rect 3103 10152 3148 10180
rect 2372 10140 2378 10152
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 1670 10112 1676 10124
rect 1510 10084 1676 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2976 10121 3004 10152
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 3418 10180 3424 10192
rect 3379 10152 3424 10180
rect 3418 10140 3424 10152
rect 3476 10180 3482 10192
rect 3694 10180 3700 10192
rect 3476 10152 3700 10180
rect 3476 10140 3482 10152
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 4028 10152 4261 10180
rect 4028 10140 4034 10152
rect 4249 10149 4261 10152
rect 4295 10149 4307 10183
rect 4249 10143 4307 10149
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 5074 10180 5080 10192
rect 4847 10152 5080 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 5074 10140 5080 10152
rect 5132 10180 5138 10192
rect 6288 10180 6316 10220
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 11330 10248 11336 10260
rect 11287 10220 11336 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 12526 10248 12532 10260
rect 12487 10220 12532 10248
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 12802 10248 12808 10260
rect 12763 10220 12808 10248
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 16390 10248 16396 10260
rect 15611 10220 16396 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16574 10248 16580 10260
rect 16531 10220 16580 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 21450 10248 21456 10260
rect 19760 10220 21456 10248
rect 19760 10208 19766 10220
rect 21450 10208 21456 10220
rect 21508 10208 21514 10260
rect 6454 10180 6460 10192
rect 5132 10152 6316 10180
rect 6415 10152 6460 10180
rect 5132 10140 5138 10152
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 8018 10180 8024 10192
rect 7979 10152 8024 10180
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 9398 10140 9404 10192
rect 9456 10180 9462 10192
rect 9858 10180 9864 10192
rect 9456 10152 9864 10180
rect 9456 10140 9462 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 9953 10183 10011 10189
rect 9953 10149 9965 10183
rect 9999 10180 10011 10183
rect 11146 10180 11152 10192
rect 9999 10152 11152 10180
rect 9999 10149 10011 10152
rect 9953 10143 10011 10149
rect 11146 10140 11152 10152
rect 11204 10180 11210 10192
rect 11517 10183 11575 10189
rect 11517 10180 11529 10183
rect 11204 10152 11529 10180
rect 11204 10140 11210 10152
rect 11517 10149 11529 10152
rect 11563 10149 11575 10183
rect 11517 10143 11575 10149
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 12768 10152 13185 10180
rect 12768 10140 12774 10152
rect 13173 10149 13185 10152
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 13811 10183 13869 10189
rect 13811 10149 13823 10183
rect 13857 10180 13869 10183
rect 14090 10180 14096 10192
rect 13857 10152 14096 10180
rect 13857 10149 13869 10152
rect 13811 10143 13869 10149
rect 14090 10140 14096 10152
rect 14148 10180 14154 10192
rect 17082 10183 17140 10189
rect 17082 10180 17094 10183
rect 14148 10152 17094 10180
rect 14148 10140 14154 10152
rect 17082 10149 17094 10152
rect 17128 10180 17140 10183
rect 17310 10180 17316 10192
rect 17128 10152 17316 10180
rect 17128 10149 17140 10152
rect 17082 10143 17140 10149
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 18693 10183 18751 10189
rect 18693 10180 18705 10183
rect 17696 10152 18705 10180
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3234 10112 3240 10124
rect 3007 10084 3240 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13446 10112 13452 10124
rect 12952 10084 13452 10112
rect 12952 10072 12958 10084
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 3510 10044 3516 10056
rect 2363 10016 3516 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4246 10044 4252 10056
rect 4203 10016 4252 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4246 10004 4252 10016
rect 4304 10044 4310 10056
rect 5534 10044 5540 10056
rect 4304 10016 5540 10044
rect 4304 10004 4310 10016
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10013 6699 10047
rect 7926 10044 7932 10056
rect 7887 10016 7932 10044
rect 6641 10007 6699 10013
rect 1762 9936 1768 9988
rect 1820 9976 1826 9988
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 1820 9948 3801 9976
rect 1820 9936 1826 9948
rect 3789 9945 3801 9948
rect 3835 9945 3847 9979
rect 3789 9939 3847 9945
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 6656 9976 6684 10007
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 8205 10007 8263 10013
rect 8220 9976 8248 10007
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11112 10016 11437 10044
rect 11112 10004 11118 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10013 11759 10047
rect 15672 10044 15700 10075
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 16761 10115 16819 10121
rect 16761 10112 16773 10115
rect 16724 10084 16773 10112
rect 16724 10072 16730 10084
rect 16761 10081 16773 10084
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 17696 10121 17724 10152
rect 18693 10149 18705 10152
rect 18739 10180 18751 10183
rect 19058 10180 19064 10192
rect 18739 10152 19064 10180
rect 18739 10149 18751 10152
rect 18693 10143 18751 10149
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 17000 10084 17693 10112
rect 17000 10072 17006 10084
rect 17681 10081 17693 10084
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 15746 10044 15752 10056
rect 15659 10016 15752 10044
rect 11701 10007 11759 10013
rect 5960 9948 8248 9976
rect 5960 9936 5966 9948
rect 5258 9908 5264 9920
rect 5219 9880 5264 9908
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 6086 9908 6092 9920
rect 6047 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 11716 9908 11744 10007
rect 15746 10004 15752 10016
rect 15804 10044 15810 10056
rect 17770 10044 17776 10056
rect 15804 10016 17776 10044
rect 15804 10004 15810 10016
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 18414 10004 18420 10056
rect 18472 10044 18478 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18472 10016 18613 10044
rect 18472 10004 18478 10016
rect 18601 10013 18613 10016
rect 18647 10013 18659 10047
rect 18874 10044 18880 10056
rect 18835 10016 18880 10044
rect 18601 10007 18659 10013
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 13814 9976 13820 9988
rect 13786 9936 13820 9976
rect 13872 9936 13878 9988
rect 15841 9979 15899 9985
rect 15841 9945 15853 9979
rect 15887 9976 15899 9979
rect 16114 9976 16120 9988
rect 15887 9948 16120 9976
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 13786 9920 13814 9936
rect 7984 9880 11744 9908
rect 7984 9868 7990 9880
rect 13722 9868 13728 9920
rect 13780 9880 13814 9920
rect 14369 9911 14427 9917
rect 13780 9868 13786 9880
rect 14369 9877 14381 9911
rect 14415 9908 14427 9911
rect 14458 9908 14464 9920
rect 14415 9880 14464 9908
rect 14415 9877 14427 9880
rect 14369 9871 14427 9877
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 1104 9818 20884 9840
rect 1104 9766 4648 9818
rect 4700 9766 4712 9818
rect 4764 9766 4776 9818
rect 4828 9766 4840 9818
rect 4892 9766 11982 9818
rect 12034 9766 12046 9818
rect 12098 9766 12110 9818
rect 12162 9766 12174 9818
rect 12226 9766 19315 9818
rect 19367 9766 19379 9818
rect 19431 9766 19443 9818
rect 19495 9766 19507 9818
rect 19559 9766 20884 9818
rect 1104 9744 20884 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 4028 9676 4445 9704
rect 4028 9664 4034 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4433 9667 4491 9673
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5316 9676 5917 9704
rect 5316 9664 5322 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 9030 9704 9036 9716
rect 8991 9676 9036 9704
rect 5905 9667 5963 9673
rect 9030 9664 9036 9676
rect 9088 9704 9094 9716
rect 9088 9676 9536 9704
rect 9088 9664 9094 9676
rect 1486 9596 1492 9648
rect 1544 9636 1550 9648
rect 2130 9636 2136 9648
rect 1544 9608 2136 9636
rect 1544 9596 1550 9608
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 5350 9636 5356 9648
rect 4580 9608 5356 9636
rect 4580 9596 4586 9608
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 6365 9639 6423 9645
rect 6365 9605 6377 9639
rect 6411 9636 6423 9639
rect 6454 9636 6460 9648
rect 6411 9608 6460 9636
rect 6411 9605 6423 9608
rect 6365 9599 6423 9605
rect 6454 9596 6460 9608
rect 6512 9636 6518 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 6512 9608 8585 9636
rect 6512 9596 6518 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 8573 9599 8631 9605
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5074 9568 5080 9580
rect 5031 9540 5080 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5074 9528 5080 9540
rect 5132 9568 5138 9580
rect 5626 9568 5632 9580
rect 5132 9540 5632 9568
rect 5132 9528 5138 9540
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 8018 9568 8024 9580
rect 7239 9540 8024 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 9508 9577 9536 9676
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 10008 9676 10425 9704
rect 10008 9664 10014 9676
rect 10413 9673 10425 9676
rect 10459 9704 10471 9707
rect 11146 9704 11152 9716
rect 10459 9676 11152 9704
rect 10459 9673 10471 9676
rect 10413 9667 10471 9673
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 15746 9704 15752 9716
rect 15707 9676 15752 9704
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16301 9707 16359 9713
rect 16301 9673 16313 9707
rect 16347 9704 16359 9707
rect 16666 9704 16672 9716
rect 16347 9676 16672 9704
rect 16347 9673 16359 9676
rect 16301 9667 16359 9673
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 19058 9704 19064 9716
rect 19019 9676 19064 9704
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11054 9636 11060 9648
rect 10827 9608 11060 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11425 9639 11483 9645
rect 11425 9605 11437 9639
rect 11471 9636 11483 9639
rect 11471 9608 12756 9636
rect 11471 9605 11483 9608
rect 11425 9599 11483 9605
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 9493 9531 9551 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12728 9568 12756 9608
rect 13446 9596 13452 9648
rect 13504 9636 13510 9648
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13504 9608 13829 9636
rect 13504 9596 13510 9608
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 15470 9636 15476 9648
rect 13817 9599 13875 9605
rect 13924 9608 15476 9636
rect 13924 9568 13952 9608
rect 15470 9596 15476 9608
rect 15528 9596 15534 9648
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 17034 9636 17040 9648
rect 16448 9608 16528 9636
rect 16995 9608 17040 9636
rect 16448 9596 16454 9608
rect 12728 9540 13952 9568
rect 14553 9571 14611 9577
rect 14553 9537 14565 9571
rect 14599 9568 14611 9571
rect 14734 9568 14740 9580
rect 14599 9540 14740 9568
rect 14599 9537 14611 9540
rect 14553 9531 14611 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 16114 9568 16120 9580
rect 15436 9540 16120 9568
rect 15436 9528 15442 9540
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 16500 9577 16528 9608
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 18414 9596 18420 9648
rect 18472 9636 18478 9648
rect 19429 9639 19487 9645
rect 19429 9636 19441 9639
rect 18472 9608 19441 9636
rect 18472 9596 18478 9608
rect 19429 9605 19441 9608
rect 19475 9605 19487 9639
rect 19429 9599 19487 9605
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18138 9568 18144 9580
rect 17644 9540 18144 9568
rect 17644 9528 17650 9540
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 18874 9568 18880 9580
rect 18831 9540 18880 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 1596 9500 1624 9528
rect 2130 9500 2136 9512
rect 1596 9472 2136 9500
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 2866 9500 2872 9512
rect 2455 9472 2872 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 2424 9432 2452 9463
rect 2866 9460 2872 9472
rect 2924 9500 2930 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 2924 9472 3249 9500
rect 2924 9460 2930 9472
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 1811 9404 2452 9432
rect 2593 9435 2651 9441
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2774 9432 2780 9444
rect 2639 9404 2780 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2774 9392 2780 9404
rect 2832 9392 2838 9444
rect 3252 9432 3280 9463
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3384 9472 3433 9500
rect 3384 9460 3390 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 7742 9500 7748 9512
rect 7699 9472 7748 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 3896 9432 3924 9463
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 11146 9460 11152 9512
rect 11204 9500 11210 9512
rect 11241 9503 11299 9509
rect 11241 9500 11253 9503
rect 11204 9472 11253 9500
rect 11204 9460 11210 9472
rect 11241 9469 11253 9472
rect 11287 9500 11299 9503
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11287 9472 11805 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 11793 9463 11851 9469
rect 19680 9503 19738 9509
rect 19680 9469 19692 9503
rect 19726 9500 19738 9503
rect 20070 9500 20076 9512
rect 19726 9472 20076 9500
rect 19726 9469 19738 9472
rect 19680 9463 19738 9469
rect 20070 9460 20076 9472
rect 20128 9500 20134 9512
rect 21542 9500 21548 9512
rect 20128 9472 21548 9500
rect 20128 9460 20134 9472
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 3252 9404 3924 9432
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 4522 9432 4528 9444
rect 4203 9404 4528 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4522 9392 4528 9404
rect 4580 9392 4586 9444
rect 4893 9435 4951 9441
rect 4893 9401 4905 9435
rect 4939 9432 4951 9435
rect 5347 9435 5405 9441
rect 5347 9432 5359 9435
rect 4939 9404 5359 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 5347 9401 5359 9404
rect 5393 9432 5405 9435
rect 6914 9432 6920 9444
rect 5393 9404 6920 9432
rect 5393 9401 5405 9404
rect 5347 9395 5405 9401
rect 6914 9392 6920 9404
rect 6972 9432 6978 9444
rect 7558 9432 7564 9444
rect 6972 9404 7564 9432
rect 6972 9392 6978 9404
rect 7558 9392 7564 9404
rect 7616 9432 7622 9444
rect 8015 9435 8073 9441
rect 8015 9432 8027 9435
rect 7616 9404 8027 9432
rect 7616 9392 7622 9404
rect 8015 9401 8027 9404
rect 8061 9432 8073 9435
rect 8846 9432 8852 9444
rect 8061 9404 8852 9432
rect 8061 9401 8073 9404
rect 8015 9395 8073 9401
rect 8846 9392 8852 9404
rect 8904 9432 8910 9444
rect 9401 9435 9459 9441
rect 9401 9432 9413 9435
rect 8904 9404 9413 9432
rect 8904 9392 8910 9404
rect 9401 9401 9413 9404
rect 9447 9432 9459 9435
rect 9855 9435 9913 9441
rect 9855 9432 9867 9435
rect 9447 9404 9867 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 9855 9401 9867 9404
rect 9901 9432 9913 9435
rect 10502 9432 10508 9444
rect 9901 9404 10508 9432
rect 9901 9401 9913 9404
rect 9855 9395 9913 9401
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12621 9435 12679 9441
rect 12621 9432 12633 9435
rect 12299 9404 12633 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12621 9401 12633 9404
rect 12667 9432 12679 9435
rect 12894 9432 12900 9444
rect 12667 9404 12900 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 14645 9435 14703 9441
rect 14645 9401 14657 9435
rect 14691 9401 14703 9435
rect 15194 9432 15200 9444
rect 15155 9404 15200 9432
rect 14645 9395 14703 9401
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3142 9364 3148 9376
rect 3007 9336 3148 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10686 9364 10692 9376
rect 10284 9336 10692 9364
rect 10284 9324 10290 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9364 13510 9376
rect 14090 9364 14096 9376
rect 13504 9336 14096 9364
rect 13504 9324 13510 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 14458 9364 14464 9376
rect 14415 9336 14464 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 14458 9324 14464 9336
rect 14516 9364 14522 9376
rect 14660 9364 14688 9395
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 18233 9435 18291 9441
rect 16632 9404 16677 9432
rect 16632 9392 16638 9404
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 15378 9364 15384 9376
rect 14516 9336 15384 9364
rect 14516 9324 14522 9336
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17368 9336 17417 9364
rect 17368 9324 17374 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17405 9327 17463 9333
rect 17770 9324 17776 9336
rect 17828 9364 17834 9376
rect 18248 9364 18276 9395
rect 17828 9336 18276 9364
rect 17828 9324 17834 9336
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 19751 9367 19809 9373
rect 19751 9364 19763 9367
rect 19576 9336 19763 9364
rect 19576 9324 19582 9336
rect 19751 9333 19763 9336
rect 19797 9333 19809 9367
rect 19751 9327 19809 9333
rect 1104 9274 20884 9296
rect 1104 9222 8315 9274
rect 8367 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 15648 9274
rect 15700 9222 15712 9274
rect 15764 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 20884 9274
rect 1104 9200 20884 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1762 9160 1768 9172
rect 1452 9132 1532 9160
rect 1452 9120 1458 9132
rect 1504 9101 1532 9132
rect 1596 9132 1768 9160
rect 1596 9101 1624 9132
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 3384 9132 3433 9160
rect 3384 9120 3390 9132
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 3421 9123 3479 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8018 9160 8024 9172
rect 7975 9132 8024 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 11606 9160 11612 9172
rect 10612 9132 11612 9160
rect 1489 9095 1547 9101
rect 1489 9061 1501 9095
rect 1535 9061 1547 9095
rect 1489 9055 1547 9061
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9061 1639 9095
rect 1581 9055 1639 9061
rect 1670 9052 1676 9104
rect 1728 9092 1734 9104
rect 2133 9095 2191 9101
rect 2133 9092 2145 9095
rect 1728 9064 2145 9092
rect 1728 9052 1734 9064
rect 2133 9061 2145 9064
rect 2179 9092 2191 9095
rect 3878 9092 3884 9104
rect 2179 9064 3884 9092
rect 2179 9061 2191 9064
rect 2133 9055 2191 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4246 9092 4252 9104
rect 4207 9064 4252 9092
rect 4246 9052 4252 9064
rect 4304 9052 4310 9104
rect 4801 9095 4859 9101
rect 4801 9061 4813 9095
rect 4847 9092 4859 9095
rect 5442 9092 5448 9104
rect 4847 9064 5448 9092
rect 4847 9061 4859 9064
rect 4801 9055 4859 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 7098 9092 7104 9104
rect 7024 9064 7104 9092
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 5626 9024 5632 9036
rect 5587 8996 5632 9024
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 7024 9033 7052 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 7371 9095 7429 9101
rect 7371 9061 7383 9095
rect 7417 9092 7429 9095
rect 7558 9092 7564 9104
rect 7417 9064 7564 9092
rect 7417 9061 7429 9064
rect 7371 9055 7429 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 10612 9101 10640 9132
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13630 9160 13636 9172
rect 13587 9132 13636 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13630 9120 13636 9132
rect 13688 9160 13694 9172
rect 14734 9160 14740 9172
rect 13688 9132 13768 9160
rect 14695 9132 14740 9160
rect 13688 9120 13694 9132
rect 10229 9095 10287 9101
rect 10229 9092 10241 9095
rect 9916 9064 10241 9092
rect 9916 9052 9922 9064
rect 10229 9061 10241 9064
rect 10275 9061 10287 9095
rect 10229 9055 10287 9061
rect 10597 9095 10655 9101
rect 10597 9061 10609 9095
rect 10643 9061 10655 9095
rect 10597 9055 10655 9061
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 10744 9064 10789 9092
rect 10744 9052 10750 9064
rect 11882 9052 11888 9104
rect 11940 9092 11946 9104
rect 12253 9095 12311 9101
rect 12253 9092 12265 9095
rect 11940 9064 12265 9092
rect 11940 9052 11946 9064
rect 12253 9061 12265 9064
rect 12299 9061 12311 9095
rect 12253 9055 12311 9061
rect 12805 9095 12863 9101
rect 12805 9061 12817 9095
rect 12851 9092 12863 9095
rect 13170 9092 13176 9104
rect 12851 9064 13176 9092
rect 12851 9061 12863 9064
rect 12805 9055 12863 9061
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 13740 9101 13768 9132
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 16485 9163 16543 9169
rect 16485 9129 16497 9163
rect 16531 9160 16543 9163
rect 16574 9160 16580 9172
rect 16531 9132 16580 9160
rect 16531 9129 16543 9132
rect 16485 9123 16543 9129
rect 16574 9120 16580 9132
rect 16632 9160 16638 9172
rect 17770 9160 17776 9172
rect 16632 9132 17776 9160
rect 16632 9120 16638 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18138 9160 18144 9172
rect 18099 9132 18144 9160
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 13725 9095 13783 9101
rect 13725 9061 13737 9095
rect 13771 9061 13783 9095
rect 13725 9055 13783 9061
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 13872 9064 13917 9092
rect 13872 9052 13878 9064
rect 14550 9052 14556 9104
rect 14608 9092 14614 9104
rect 15010 9092 15016 9104
rect 14608 9064 15016 9092
rect 14608 9052 14614 9064
rect 15010 9052 15016 9064
rect 15068 9052 15074 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15473 9095 15531 9101
rect 15473 9092 15485 9095
rect 15436 9064 15485 9092
rect 15436 9052 15442 9064
rect 15473 9061 15485 9064
rect 15519 9061 15531 9095
rect 15473 9055 15531 9061
rect 17215 9095 17273 9101
rect 17215 9061 17227 9095
rect 17261 9092 17273 9095
rect 17310 9092 17316 9104
rect 17261 9064 17316 9092
rect 17261 9061 17273 9064
rect 17215 9055 17273 9061
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 18782 9092 18788 9104
rect 18743 9064 18788 9092
rect 18782 9052 18788 9064
rect 18840 9052 18846 9104
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6696 8996 7021 9024
rect 6696 8984 6702 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 7984 8996 8217 9024
rect 7984 8984 7990 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 16850 9024 16856 9036
rect 16811 8996 16856 9024
rect 8205 8987 8263 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2682 8956 2688 8968
rect 2280 8928 2688 8956
rect 2280 8916 2286 8928
rect 2682 8916 2688 8928
rect 2740 8956 2746 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 2740 8928 3801 8956
rect 2740 8916 2746 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 3789 8919 3847 8925
rect 3988 8928 4169 8956
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 3326 8888 3332 8900
rect 2915 8860 3332 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 2130 8780 2136 8832
rect 2188 8820 2194 8832
rect 2409 8823 2467 8829
rect 2409 8820 2421 8823
rect 2188 8792 2421 8820
rect 2188 8780 2194 8792
rect 2409 8789 2421 8792
rect 2455 8789 2467 8823
rect 2409 8783 2467 8789
rect 3099 8823 3157 8829
rect 3099 8789 3111 8823
rect 3145 8820 3157 8823
rect 3234 8820 3240 8832
rect 3145 8792 3240 8820
rect 3145 8789 3157 8792
rect 3099 8783 3157 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 3988 8820 4016 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 5644 8956 5672 8984
rect 7834 8956 7840 8968
rect 5644 8928 7840 8956
rect 4157 8919 4215 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 10652 8928 11897 8956
rect 10652 8916 10658 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 6641 8891 6699 8897
rect 6641 8888 6653 8891
rect 5368 8860 6653 8888
rect 5368 8820 5396 8860
rect 6641 8857 6653 8860
rect 6687 8888 6699 8891
rect 6914 8888 6920 8900
rect 6687 8860 6920 8888
rect 6687 8857 6699 8860
rect 6641 8851 6699 8857
rect 6914 8848 6920 8860
rect 6972 8848 6978 8900
rect 11146 8888 11152 8900
rect 11107 8860 11152 8888
rect 11146 8848 11152 8860
rect 11204 8888 11210 8900
rect 12176 8888 12204 8919
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15160 8928 15393 8956
rect 15160 8916 15166 8928
rect 15381 8925 15393 8928
rect 15427 8956 15439 8959
rect 15838 8956 15844 8968
rect 15427 8928 15844 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 17920 8928 18705 8956
rect 17920 8916 17926 8928
rect 18693 8925 18705 8928
rect 18739 8956 18751 8959
rect 19518 8956 19524 8968
rect 18739 8928 19524 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 12618 8888 12624 8900
rect 11204 8860 12624 8888
rect 11204 8848 11210 8860
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 14277 8891 14335 8897
rect 14277 8857 14289 8891
rect 14323 8888 14335 8891
rect 14642 8888 14648 8900
rect 14323 8860 14648 8888
rect 14323 8857 14335 8860
rect 14277 8851 14335 8857
rect 14642 8848 14648 8860
rect 14700 8888 14706 8900
rect 16040 8888 16068 8916
rect 14700 8860 16068 8888
rect 14700 8848 14706 8860
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 19245 8891 19303 8897
rect 19245 8888 19257 8891
rect 19116 8860 19257 8888
rect 19116 8848 19122 8860
rect 19245 8857 19257 8860
rect 19291 8857 19303 8891
rect 19245 8851 19303 8857
rect 3936 8792 5396 8820
rect 5767 8823 5825 8829
rect 3936 8780 3942 8792
rect 5767 8789 5779 8823
rect 5813 8820 5825 8823
rect 5994 8820 6000 8832
rect 5813 8792 6000 8820
rect 5813 8789 5825 8792
rect 5767 8783 5825 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6362 8820 6368 8832
rect 6323 8792 6368 8820
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12710 8820 12716 8832
rect 11848 8792 12716 8820
rect 11848 8780 11854 8792
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 1104 8730 20884 8752
rect 1104 8678 4648 8730
rect 4700 8678 4712 8730
rect 4764 8678 4776 8730
rect 4828 8678 4840 8730
rect 4892 8678 11982 8730
rect 12034 8678 12046 8730
rect 12098 8678 12110 8730
rect 12162 8678 12174 8730
rect 12226 8678 19315 8730
rect 19367 8678 19379 8730
rect 19431 8678 19443 8730
rect 19495 8678 19507 8730
rect 19559 8678 20884 8730
rect 1104 8656 20884 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2096 8588 2697 8616
rect 2096 8576 2102 8588
rect 2685 8585 2697 8588
rect 2731 8616 2743 8619
rect 2958 8616 2964 8628
rect 2731 8588 2964 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 3743 8588 4169 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 4157 8585 4169 8588
rect 4203 8616 4215 8619
rect 4246 8616 4252 8628
rect 4203 8588 4252 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 6270 8616 6276 8628
rect 4540 8588 6276 8616
rect 4540 8548 4568 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6638 8616 6644 8628
rect 6599 8588 6644 8616
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 10226 8616 10232 8628
rect 10187 8588 10232 8616
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10468 8588 10609 8616
rect 10468 8576 10474 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 10597 8579 10655 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12986 8616 12992 8628
rect 12947 8588 12992 8616
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 16908 8588 17233 8616
rect 16908 8576 16914 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17221 8579 17279 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18414 8616 18420 8628
rect 18327 8588 18420 8616
rect 18414 8576 18420 8588
rect 18472 8616 18478 8628
rect 18782 8616 18788 8628
rect 18472 8588 18788 8616
rect 18472 8576 18478 8588
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 19610 8616 19616 8628
rect 19571 8588 19616 8616
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 6086 8548 6092 8560
rect 2602 8520 4568 8548
rect 4632 8520 6092 8548
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 2602 8480 2630 8520
rect 2774 8480 2780 8492
rect 1636 8452 2630 8480
rect 2735 8452 2780 8480
rect 1636 8440 1642 8452
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 4632 8489 4660 8520
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 6362 8508 6368 8560
rect 6420 8548 6426 8560
rect 8297 8551 8355 8557
rect 8297 8548 8309 8551
rect 6420 8520 8309 8548
rect 6420 8508 6426 8520
rect 8297 8517 8309 8520
rect 8343 8548 8355 8551
rect 8343 8520 9996 8548
rect 8343 8517 8355 8520
rect 8297 8511 8355 8517
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5442 8480 5448 8492
rect 5307 8452 5448 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7524 8452 7757 8480
rect 7524 8440 7530 8452
rect 7745 8449 7757 8452
rect 7791 8480 7803 8483
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 7791 8452 8677 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9968 8489 9996 8520
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 9180 8452 9321 8480
rect 9180 8440 9186 8452
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10134 8480 10140 8492
rect 9999 8452 10140 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10594 8440 10600 8492
rect 10652 8480 10658 8492
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10652 8452 10885 8480
rect 10652 8440 10658 8452
rect 10873 8449 10885 8452
rect 10919 8449 10931 8483
rect 11146 8480 11152 8492
rect 11107 8452 11152 8480
rect 10873 8443 10931 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13320 8452 13814 8480
rect 13320 8440 13326 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 5626 8412 5632 8424
rect 1443 8384 2084 8412
rect 5587 8384 5632 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2056 8285 2084 8384
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12584 8384 12817 8412
rect 12584 8372 12590 8384
rect 12805 8381 12817 8384
rect 12851 8412 12863 8415
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 12851 8384 13369 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 13357 8381 13369 8384
rect 13403 8381 13415 8415
rect 13786 8412 13814 8452
rect 15010 8440 15016 8492
rect 15068 8480 15074 8492
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15068 8452 15761 8480
rect 15068 8440 15074 8452
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 16022 8480 16028 8492
rect 15983 8452 16028 8480
rect 15749 8443 15807 8449
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 19628 8480 19656 8576
rect 18647 8452 19656 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 13906 8412 13912 8424
rect 13786 8384 13912 8412
rect 13357 8375 13415 8381
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 3139 8347 3197 8353
rect 3139 8313 3151 8347
rect 3185 8344 3197 8347
rect 3326 8344 3332 8356
rect 3185 8316 3332 8344
rect 3185 8313 3197 8316
rect 3139 8307 3197 8313
rect 3326 8304 3332 8316
rect 3384 8344 3390 8356
rect 3384 8316 4568 8344
rect 3384 8304 3390 8316
rect 2041 8279 2099 8285
rect 2041 8245 2053 8279
rect 2087 8276 2099 8279
rect 4062 8276 4068 8288
rect 2087 8248 4068 8276
rect 2087 8245 2099 8248
rect 2041 8239 2099 8245
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4540 8276 4568 8316
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 7101 8347 7159 8353
rect 4764 8316 4809 8344
rect 4764 8304 4770 8316
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7558 8344 7564 8356
rect 7147 8316 7564 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8313 9459 8347
rect 9401 8307 9459 8313
rect 5074 8276 5080 8288
rect 4540 8248 5080 8276
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5994 8276 6000 8288
rect 5955 8248 6000 8276
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 7466 8276 7472 8288
rect 7427 8248 7472 8276
rect 7466 8236 7472 8248
rect 7524 8276 7530 8288
rect 7852 8276 7880 8307
rect 9030 8276 9036 8288
rect 7524 8248 7880 8276
rect 8991 8248 9036 8276
rect 7524 8236 7530 8248
rect 9030 8236 9036 8248
rect 9088 8276 9094 8288
rect 9416 8276 9444 8307
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10965 8347 11023 8353
rect 10965 8344 10977 8347
rect 10468 8316 10977 8344
rect 10468 8304 10474 8316
rect 10965 8313 10977 8316
rect 11011 8313 11023 8347
rect 14230 8347 14288 8353
rect 14230 8344 14242 8347
rect 10965 8307 11023 8313
rect 13740 8316 14242 8344
rect 9088 8248 9444 8276
rect 9088 8236 9094 8248
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 10134 8276 10140 8288
rect 9824 8248 10140 8276
rect 9824 8236 9830 8248
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11940 8248 12081 8276
rect 11940 8236 11946 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 13630 8276 13636 8288
rect 13504 8248 13636 8276
rect 13504 8236 13510 8248
rect 13630 8236 13636 8248
rect 13688 8276 13694 8288
rect 13740 8285 13768 8316
rect 14230 8313 14242 8316
rect 14276 8313 14288 8347
rect 14230 8307 14288 8313
rect 15841 8347 15899 8353
rect 15841 8313 15853 8347
rect 15887 8313 15899 8347
rect 15841 8307 15899 8313
rect 18693 8347 18751 8353
rect 18693 8313 18705 8347
rect 18739 8313 18751 8347
rect 18693 8307 18751 8313
rect 13725 8279 13783 8285
rect 13725 8276 13737 8279
rect 13688 8248 13737 8276
rect 13688 8236 13694 8248
rect 13725 8245 13737 8248
rect 13771 8245 13783 8279
rect 13725 8239 13783 8245
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14829 8279 14887 8285
rect 14829 8276 14841 8279
rect 13872 8248 14841 8276
rect 13872 8236 13878 8248
rect 14829 8245 14841 8248
rect 14875 8245 14887 8279
rect 14829 8239 14887 8245
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 15856 8276 15884 8307
rect 15528 8248 15884 8276
rect 16945 8279 17003 8285
rect 15528 8236 15534 8248
rect 16945 8245 16957 8279
rect 16991 8276 17003 8279
rect 17310 8276 17316 8288
rect 16991 8248 17316 8276
rect 16991 8245 17003 8248
rect 16945 8239 17003 8245
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 18708 8276 18736 8307
rect 19058 8304 19064 8356
rect 19116 8344 19122 8356
rect 19245 8347 19303 8353
rect 19245 8344 19257 8347
rect 19116 8316 19257 8344
rect 19116 8304 19122 8316
rect 19245 8313 19257 8316
rect 19291 8313 19303 8347
rect 19245 8307 19303 8313
rect 18564 8248 18736 8276
rect 18564 8236 18570 8248
rect 1104 8186 20884 8208
rect 1104 8134 8315 8186
rect 8367 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 15648 8186
rect 15700 8134 15712 8186
rect 15764 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 20884 8186
rect 1104 8112 20884 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1452 8044 1961 8072
rect 1452 8032 1458 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2832 8044 3433 8072
rect 2832 8032 2838 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 3421 8035 3479 8041
rect 4126 8044 4629 8072
rect 1670 8004 1676 8016
rect 1583 7976 1676 8004
rect 1670 7964 1676 7976
rect 1728 8004 1734 8016
rect 2587 8007 2645 8013
rect 2587 8004 2599 8007
rect 1728 7976 2599 8004
rect 1728 7964 1734 7976
rect 2587 7973 2599 7976
rect 2633 8004 2645 8007
rect 3326 8004 3332 8016
rect 2633 7976 3332 8004
rect 2633 7973 2645 7976
rect 2587 7967 2645 7973
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2406 7936 2412 7948
rect 2271 7908 2412 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 4126 7936 4154 8044
rect 4617 8041 4629 8044
rect 4663 8072 4675 8075
rect 4706 8072 4712 8084
rect 4663 8044 4712 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 5132 8044 5181 8072
rect 5132 8032 5138 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 8846 8072 8852 8084
rect 6328 8044 8852 8072
rect 6328 8032 6334 8044
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 9180 8044 9229 8072
rect 9180 8032 9186 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 9364 8044 10057 8072
rect 9364 8032 9370 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 10045 8035 10103 8041
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 10284 8044 12081 8072
rect 10284 8032 10290 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 13964 8044 14657 8072
rect 13964 8032 13970 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 14645 8035 14703 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16482 8072 16488 8084
rect 16439 8044 16488 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17494 8072 17500 8084
rect 17000 8044 17500 8072
rect 17000 8032 17006 8044
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 7463 8007 7521 8013
rect 7463 7973 7475 8007
rect 7509 8004 7521 8007
rect 7558 8004 7564 8016
rect 7509 7976 7564 8004
rect 7509 7973 7521 7976
rect 7463 7967 7521 7973
rect 7558 7964 7564 7976
rect 7616 7964 7622 8016
rect 11511 8007 11569 8013
rect 11511 7973 11523 8007
rect 11557 8004 11569 8007
rect 11790 8004 11796 8016
rect 11557 7976 11796 8004
rect 11557 7973 11569 7976
rect 11511 7967 11569 7973
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 13541 8007 13599 8013
rect 13541 7973 13553 8007
rect 13587 8004 13599 8007
rect 13814 8004 13820 8016
rect 13587 7976 13820 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13814 7964 13820 7976
rect 13872 8004 13878 8016
rect 15470 8004 15476 8016
rect 13872 7976 13917 8004
rect 15431 7976 15476 8004
rect 13872 7964 13878 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 17194 8007 17252 8013
rect 17194 7973 17206 8007
rect 17240 8004 17252 8007
rect 17310 8004 17316 8016
rect 17240 7976 17316 8004
rect 17240 7973 17252 7976
rect 17194 7967 17252 7973
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 18506 7964 18512 8016
rect 18564 8004 18570 8016
rect 18877 8007 18935 8013
rect 18877 8004 18889 8007
rect 18564 7976 18889 8004
rect 18564 7964 18570 7976
rect 18877 7973 18889 7976
rect 18923 7973 18935 8007
rect 18877 7967 18935 7973
rect 3191 7908 4154 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4580 7908 4813 7936
rect 4580 7896 4586 7908
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 9766 7936 9772 7948
rect 9727 7908 9772 7936
rect 4801 7899 4859 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7936 10011 7939
rect 10689 7939 10747 7945
rect 10689 7936 10701 7939
rect 9999 7908 10701 7936
rect 9999 7905 10011 7908
rect 9953 7899 10011 7905
rect 10689 7905 10701 7908
rect 10735 7936 10747 7939
rect 12618 7936 12624 7948
rect 10735 7908 12624 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 2424 7868 2452 7896
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 2424 7840 3801 7868
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 6270 7828 6276 7880
rect 6328 7868 6334 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 6328 7840 7113 7868
rect 6328 7828 6334 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9582 7868 9588 7880
rect 9180 7840 9588 7868
rect 9180 7828 9186 7840
rect 9582 7828 9588 7840
rect 9640 7868 9646 7880
rect 9968 7868 9996 7899
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 16945 7939 17003 7945
rect 16945 7936 16957 7939
rect 16816 7908 16957 7936
rect 16816 7896 16822 7908
rect 16945 7905 16957 7908
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7936 17923 7939
rect 18414 7936 18420 7948
rect 17911 7908 18420 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 9640 7840 9996 7868
rect 11072 7840 11161 7868
rect 9640 7828 9646 7840
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 4126 7772 6009 7800
rect 1302 7692 1308 7744
rect 1360 7732 1366 7744
rect 4126 7732 4154 7772
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 5997 7763 6055 7769
rect 6098 7772 6960 7800
rect 1360 7704 4154 7732
rect 1360 7692 1366 7704
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 5721 7735 5779 7741
rect 5721 7732 5733 7735
rect 5408 7704 5733 7732
rect 5408 7692 5414 7704
rect 5721 7701 5733 7704
rect 5767 7732 5779 7735
rect 6098 7732 6126 7772
rect 6362 7732 6368 7744
rect 5767 7704 6126 7732
rect 6323 7704 6368 7732
rect 5767 7701 5779 7704
rect 5721 7695 5779 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 6932 7741 6960 7772
rect 11072 7744 11100 7840
rect 11149 7837 11161 7840
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7868 13231 7871
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13219 7840 13737 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 13725 7837 13737 7840
rect 13771 7868 13783 7871
rect 14826 7868 14832 7880
rect 13771 7840 14832 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 15378 7868 15384 7880
rect 15339 7840 15384 7868
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 14277 7803 14335 7809
rect 14277 7769 14289 7803
rect 14323 7800 14335 7803
rect 15194 7800 15200 7812
rect 14323 7772 15200 7800
rect 14323 7769 14335 7772
rect 14277 7763 14335 7769
rect 15194 7760 15200 7772
rect 15252 7800 15258 7812
rect 15672 7800 15700 7831
rect 17954 7828 17960 7880
rect 18012 7868 18018 7880
rect 18782 7868 18788 7880
rect 18012 7840 18788 7868
rect 18012 7828 18018 7840
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 19061 7871 19119 7877
rect 19061 7868 19073 7871
rect 18932 7840 19073 7868
rect 18932 7828 18938 7840
rect 19061 7837 19073 7840
rect 19107 7837 19119 7871
rect 19061 7831 19119 7837
rect 15252 7772 15700 7800
rect 15252 7760 15258 7772
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7006 7732 7012 7744
rect 6963 7704 7012 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7524 7704 8033 7732
rect 7524 7692 7530 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8570 7732 8576 7744
rect 8531 7704 8576 7732
rect 8021 7695 8079 7701
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 11054 7732 11060 7744
rect 11015 7704 11060 7732
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 12342 7732 12348 7744
rect 12303 7704 12348 7732
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 18506 7732 18512 7744
rect 18467 7704 18512 7732
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 1104 7642 20884 7664
rect 1104 7590 4648 7642
rect 4700 7590 4712 7642
rect 4764 7590 4776 7642
rect 4828 7590 4840 7642
rect 4892 7590 11982 7642
rect 12034 7590 12046 7642
rect 12098 7590 12110 7642
rect 12162 7590 12174 7642
rect 12226 7590 19315 7642
rect 19367 7590 19379 7642
rect 19431 7590 19443 7642
rect 19495 7590 19507 7642
rect 19559 7590 20884 7642
rect 1104 7568 20884 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 1820 7500 2329 7528
rect 1820 7488 1826 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2685 7531 2743 7537
rect 2685 7497 2697 7531
rect 2731 7528 2743 7531
rect 3326 7528 3332 7540
rect 2731 7500 3332 7528
rect 2731 7497 2743 7500
rect 2685 7491 2743 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 4580 7500 6193 7528
rect 4580 7488 4586 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 6181 7491 6239 7497
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 10100 7500 12449 7528
rect 10100 7488 10106 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12802 7528 12808 7540
rect 12763 7500 12808 7528
rect 12437 7491 12495 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 14829 7531 14887 7537
rect 14829 7497 14841 7531
rect 14875 7528 14887 7531
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 14875 7500 15393 7528
rect 14875 7497 14887 7500
rect 14829 7491 14887 7497
rect 15381 7497 15393 7500
rect 15427 7528 15439 7531
rect 15470 7528 15476 7540
rect 15427 7500 15476 7528
rect 15427 7497 15439 7500
rect 15381 7491 15439 7497
rect 15470 7488 15476 7500
rect 15528 7528 15534 7540
rect 15657 7531 15715 7537
rect 15657 7528 15669 7531
rect 15528 7500 15669 7528
rect 15528 7488 15534 7500
rect 15657 7497 15669 7500
rect 15703 7497 15715 7531
rect 15657 7491 15715 7497
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 16298 7528 16304 7540
rect 16255 7500 16304 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 16816 7500 17693 7528
rect 16816 7488 16822 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 18414 7528 18420 7540
rect 18375 7500 18420 7528
rect 17681 7491 17739 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 18506 7488 18512 7540
rect 18564 7528 18570 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 18564 7500 19533 7528
rect 18564 7488 18570 7500
rect 19521 7497 19533 7500
rect 19567 7497 19579 7531
rect 19521 7491 19579 7497
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 5184 7432 5825 7460
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 1360 7364 1409 7392
rect 1360 7352 1366 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 5184 7392 5212 7432
rect 5813 7429 5825 7432
rect 5859 7460 5871 7463
rect 6086 7460 6092 7472
rect 5859 7432 6092 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 11517 7463 11575 7469
rect 11517 7429 11529 7463
rect 11563 7460 11575 7463
rect 11882 7460 11888 7472
rect 11563 7432 11888 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 11882 7420 11888 7432
rect 11940 7460 11946 7472
rect 13446 7460 13452 7472
rect 11940 7432 13452 7460
rect 11940 7420 11946 7432
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 3927 7364 5212 7392
rect 5261 7395 5319 7401
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5994 7392 6000 7404
rect 5307 7364 6000 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6972 7364 7205 7392
rect 6972 7352 6978 7364
rect 7193 7361 7205 7364
rect 7239 7392 7251 7395
rect 7282 7392 7288 7404
rect 7239 7364 7288 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 11146 7392 11152 7404
rect 10643 7364 11152 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 11146 7352 11152 7364
rect 11204 7392 11210 7404
rect 12342 7392 12348 7404
rect 11204 7364 12348 7392
rect 11204 7352 11210 7364
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 16316 7392 16344 7488
rect 18782 7420 18788 7472
rect 18840 7460 18846 7472
rect 19889 7463 19947 7469
rect 19889 7460 19901 7463
rect 18840 7432 19901 7460
rect 18840 7420 18846 7432
rect 19889 7429 19901 7432
rect 19935 7429 19947 7463
rect 19889 7423 19947 7429
rect 18601 7395 18659 7401
rect 16316 7364 16804 7392
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8570 7324 8576 7336
rect 8527 7296 8576 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8570 7284 8576 7296
rect 8628 7324 8634 7336
rect 12437 7327 12495 7333
rect 8628 7296 11514 7324
rect 8628 7284 8634 7296
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3237 7259 3295 7265
rect 3237 7256 3249 7259
rect 3016 7228 3249 7256
rect 3016 7216 3022 7228
rect 3237 7225 3249 7228
rect 3283 7225 3295 7259
rect 3237 7219 3295 7225
rect 3326 7216 3332 7268
rect 3384 7256 3390 7268
rect 4525 7259 4583 7265
rect 3384 7228 3429 7256
rect 3384 7216 3390 7228
rect 4525 7225 4537 7259
rect 4571 7256 4583 7259
rect 5350 7256 5356 7268
rect 4571 7228 5356 7256
rect 4571 7225 4583 7228
rect 4525 7219 4583 7225
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 6914 7256 6920 7268
rect 5460 7228 6684 7256
rect 6875 7228 6920 7256
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 1765 7191 1823 7197
rect 1765 7188 1777 7191
rect 1728 7160 1777 7188
rect 1728 7148 1734 7160
rect 1765 7157 1777 7160
rect 1811 7157 1823 7191
rect 1765 7151 1823 7157
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3344 7188 3372 7216
rect 3099 7160 3372 7188
rect 4893 7191 4951 7197
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 5074 7188 5080 7200
rect 4939 7160 5080 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 5074 7148 5080 7160
rect 5132 7188 5138 7200
rect 5460 7188 5488 7228
rect 5132 7160 5488 7188
rect 5132 7148 5138 7160
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6328 7160 6561 7188
rect 6328 7148 6334 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 6656 7188 6684 7228
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7064 7228 7109 7256
rect 7064 7216 7070 7228
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7616 7228 7941 7256
rect 7616 7216 7622 7228
rect 7929 7225 7941 7228
rect 7975 7256 7987 7259
rect 8389 7259 8447 7265
rect 8389 7256 8401 7259
rect 7975 7228 8401 7256
rect 7975 7225 7987 7228
rect 7929 7219 7987 7225
rect 8389 7225 8401 7228
rect 8435 7256 8447 7259
rect 8843 7259 8901 7265
rect 8843 7256 8855 7259
rect 8435 7228 8855 7256
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 8843 7225 8855 7228
rect 8889 7256 8901 7259
rect 10502 7256 10508 7268
rect 8889 7228 10508 7256
rect 8889 7225 8901 7228
rect 8843 7219 8901 7225
rect 10502 7216 10508 7228
rect 10560 7256 10566 7268
rect 10959 7259 11017 7265
rect 10959 7256 10971 7259
rect 10560 7228 10971 7256
rect 10560 7216 10566 7228
rect 10959 7225 10971 7228
rect 11005 7225 11017 7259
rect 11486 7256 11514 7296
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12483 7296 12725 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12713 7293 12725 7296
rect 12759 7324 12771 7327
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 12759 7296 13369 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 13357 7293 13369 7296
rect 13403 7324 13415 7327
rect 13909 7327 13967 7333
rect 13403 7296 13814 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 12342 7256 12348 7268
rect 11486 7228 12348 7256
rect 10959 7219 11017 7225
rect 7576 7188 7604 7216
rect 6656 7160 7604 7188
rect 6549 7151 6607 7157
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 9088 7160 9413 7188
rect 9088 7148 9094 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9401 7151 9459 7157
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10980 7188 11008 7219
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 12529 7259 12587 7265
rect 12529 7225 12541 7259
rect 12575 7225 12587 7259
rect 13786 7256 13814 7296
rect 13909 7293 13921 7327
rect 13955 7324 13967 7327
rect 13998 7324 14004 7336
rect 13955 7296 14004 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 16482 7324 16488 7336
rect 16443 7296 16488 7324
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 16776 7333 16804 7364
rect 18601 7361 18613 7395
rect 18647 7392 18659 7395
rect 18690 7392 18696 7404
rect 18647 7364 18696 7392
rect 18647 7361 18659 7364
rect 18601 7355 18659 7361
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 18874 7392 18880 7404
rect 18835 7364 18880 7392
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 14458 7256 14464 7268
rect 13786 7228 14464 7256
rect 12529 7219 12587 7225
rect 11882 7188 11888 7200
rect 10980 7160 11888 7188
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12544 7188 12572 7219
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 17037 7259 17095 7265
rect 17037 7225 17049 7259
rect 17083 7256 17095 7259
rect 18138 7256 18144 7268
rect 17083 7228 18144 7256
rect 17083 7225 17095 7228
rect 17037 7219 17095 7225
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18693 7259 18751 7265
rect 18693 7225 18705 7259
rect 18739 7225 18751 7259
rect 18693 7219 18751 7225
rect 13262 7188 13268 7200
rect 12299 7160 13268 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 13688 7160 13737 7188
rect 13688 7148 13694 7160
rect 13725 7157 13737 7160
rect 13771 7188 13783 7191
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 13771 7160 14289 7188
rect 13771 7157 13783 7160
rect 13725 7151 13783 7157
rect 14277 7157 14289 7160
rect 14323 7157 14335 7191
rect 17310 7188 17316 7200
rect 17271 7160 17316 7188
rect 14277 7151 14335 7157
rect 17310 7148 17316 7160
rect 17368 7148 17374 7200
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 18708 7188 18736 7219
rect 18472 7160 18736 7188
rect 18472 7148 18478 7160
rect 1104 7098 20884 7120
rect 1104 7046 8315 7098
rect 8367 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 15648 7098
rect 15700 7046 15712 7098
rect 15764 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 20884 7098
rect 1104 7024 20884 7046
rect 1535 6987 1593 6993
rect 1535 6953 1547 6987
rect 1581 6984 1593 6987
rect 6733 6987 6791 6993
rect 6733 6984 6745 6987
rect 1581 6956 6745 6984
rect 1581 6953 1593 6956
rect 1535 6947 1593 6953
rect 6733 6953 6745 6956
rect 6779 6984 6791 6987
rect 6914 6984 6920 6996
rect 6779 6956 6920 6984
rect 6779 6953 6791 6956
rect 6733 6947 6791 6953
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 8938 6984 8944 6996
rect 7708 6956 8944 6984
rect 7708 6944 7714 6956
rect 8938 6944 8944 6956
rect 8996 6984 9002 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8996 6956 9045 6984
rect 8996 6944 9002 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 11054 6984 11060 6996
rect 11015 6956 11060 6984
rect 9033 6947 9091 6953
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 11882 6944 11888 6996
rect 11940 6984 11946 6996
rect 13630 6984 13636 6996
rect 11940 6956 13636 6984
rect 11940 6944 11946 6956
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 13872 6956 13921 6984
rect 13872 6944 13878 6956
rect 13909 6953 13921 6956
rect 13955 6953 13967 6987
rect 13909 6947 13967 6953
rect 13998 6944 14004 6996
rect 14056 6984 14062 6996
rect 14369 6987 14427 6993
rect 14369 6984 14381 6987
rect 14056 6956 14381 6984
rect 14056 6944 14062 6956
rect 14369 6953 14381 6956
rect 14415 6984 14427 6987
rect 17402 6984 17408 6996
rect 14415 6956 17408 6984
rect 14415 6953 14427 6956
rect 14369 6947 14427 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 17865 6987 17923 6993
rect 17865 6953 17877 6987
rect 17911 6984 17923 6987
rect 18506 6984 18512 6996
rect 17911 6956 18512 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 18601 6987 18659 6993
rect 18601 6953 18613 6987
rect 18647 6984 18659 6987
rect 18690 6984 18696 6996
rect 18647 6956 18696 6984
rect 18647 6953 18659 6956
rect 18601 6947 18659 6953
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 1946 6916 1952 6928
rect 1907 6888 1952 6916
rect 1946 6876 1952 6888
rect 2004 6876 2010 6928
rect 2222 6916 2228 6928
rect 2183 6888 2228 6916
rect 2222 6876 2228 6888
rect 2280 6876 2286 6928
rect 2593 6919 2651 6925
rect 2593 6885 2605 6919
rect 2639 6916 2651 6919
rect 3326 6916 3332 6928
rect 2639 6888 3332 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 3786 6876 3792 6928
rect 3844 6916 3850 6928
rect 4709 6919 4767 6925
rect 3844 6888 4108 6916
rect 3844 6876 3850 6888
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 1578 6848 1584 6860
rect 1510 6820 1584 6848
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3878 6848 3884 6860
rect 3191 6820 3884 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 4080 6857 4108 6888
rect 4709 6885 4721 6919
rect 4755 6916 4767 6919
rect 5074 6916 5080 6928
rect 4755 6888 5080 6916
rect 4755 6885 4767 6888
rect 4709 6879 4767 6885
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 5537 6919 5595 6925
rect 5537 6885 5549 6919
rect 5583 6916 5595 6919
rect 6638 6916 6644 6928
rect 5583 6888 6644 6916
rect 5583 6885 5595 6888
rect 5537 6879 5595 6885
rect 6638 6876 6644 6888
rect 6696 6916 6702 6928
rect 7101 6919 7159 6925
rect 7101 6916 7113 6919
rect 6696 6888 7113 6916
rect 6696 6876 6702 6888
rect 7101 6885 7113 6888
rect 7147 6885 7159 6919
rect 12894 6916 12900 6928
rect 12855 6888 12900 6916
rect 7101 6879 7159 6885
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 17307 6919 17365 6925
rect 17307 6885 17319 6919
rect 17353 6885 17365 6919
rect 17307 6879 17365 6885
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4154 6848 4160 6860
rect 4111 6820 4160 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 8481 6851 8539 6857
rect 6144 6820 6189 6848
rect 6144 6808 6150 6820
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8662 6848 8668 6860
rect 8527 6820 8668 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 8904 6820 9873 6848
rect 8904 6808 8910 6820
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10928 6820 10977 6848
rect 10928 6808 10934 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 11790 6848 11796 6860
rect 11751 6820 11796 6848
rect 10965 6811 11023 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 15286 6808 15292 6860
rect 15344 6848 15350 6860
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15344 6820 15393 6848
rect 15344 6808 15350 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15930 6848 15936 6860
rect 15843 6820 15936 6848
rect 15381 6811 15439 6817
rect 15930 6808 15936 6820
rect 15988 6848 15994 6860
rect 16298 6848 16304 6860
rect 15988 6820 16304 6848
rect 15988 6808 15994 6820
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 17322 6848 17350 6879
rect 18782 6876 18788 6928
rect 18840 6916 18846 6928
rect 18877 6919 18935 6925
rect 18877 6916 18889 6919
rect 18840 6888 18889 6916
rect 18840 6876 18846 6888
rect 18877 6885 18889 6888
rect 18923 6885 18935 6919
rect 18877 6879 18935 6885
rect 17402 6848 17408 6860
rect 17322 6820 17408 6848
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1728 6752 2513 6780
rect 1728 6740 1734 6752
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5810 6780 5816 6792
rect 5491 6752 5816 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5810 6740 5816 6752
rect 5868 6780 5874 6792
rect 6362 6780 6368 6792
rect 5868 6752 6368 6780
rect 5868 6740 5874 6752
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7282 6780 7288 6792
rect 7243 6752 7288 6780
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10686 6780 10692 6792
rect 10551 6752 10692 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10686 6740 10692 6752
rect 10744 6780 10750 6792
rect 11698 6780 11704 6792
rect 10744 6752 11704 6780
rect 10744 6740 10750 6752
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16163 6752 16957 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16945 6749 16957 6752
rect 16991 6780 17003 6783
rect 17770 6780 17776 6792
rect 16991 6752 17776 6780
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 3016 6684 5206 6712
rect 3016 6672 3022 6684
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 3384 6616 3433 6644
rect 3384 6604 3390 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3421 6607 3479 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4246 6644 4252 6656
rect 4207 6616 4252 6644
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4982 6644 4988 6656
rect 4943 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5178 6644 5206 6684
rect 6178 6672 6184 6724
rect 6236 6712 6242 6724
rect 7190 6712 7196 6724
rect 6236 6684 7196 6712
rect 6236 6672 6242 6684
rect 7190 6672 7196 6684
rect 7248 6712 7254 6724
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7248 6684 7941 6712
rect 7248 6672 7254 6684
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 7929 6675 7987 6681
rect 8665 6715 8723 6721
rect 8665 6681 8677 6715
rect 8711 6712 8723 6715
rect 11054 6712 11060 6724
rect 8711 6684 11060 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 15378 6712 15384 6724
rect 14240 6684 15384 6712
rect 14240 6672 14246 6684
rect 15378 6672 15384 6684
rect 15436 6712 15442 6724
rect 16393 6715 16451 6721
rect 16393 6712 16405 6715
rect 15436 6684 16405 6712
rect 15436 6672 15442 6684
rect 16393 6681 16405 6684
rect 16439 6681 16451 6715
rect 18800 6712 18828 6743
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 19061 6783 19119 6789
rect 19061 6780 19073 6783
rect 18932 6752 19073 6780
rect 18932 6740 18938 6752
rect 19061 6749 19073 6752
rect 19107 6749 19119 6783
rect 19061 6743 19119 6749
rect 19610 6712 19616 6724
rect 18800 6684 19616 6712
rect 16393 6675 16451 6681
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 5178 6616 6377 6644
rect 6365 6613 6377 6616
rect 6411 6613 6423 6647
rect 10042 6644 10048 6656
rect 10003 6616 10048 6644
rect 6365 6607 6423 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 10652 6616 10793 6644
rect 10652 6604 10658 6616
rect 10781 6613 10793 6616
rect 10827 6613 10839 6647
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 10781 6607 10839 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 16761 6647 16819 6653
rect 16761 6644 16773 6647
rect 16540 6616 16773 6644
rect 16540 6604 16546 6616
rect 16761 6613 16773 6616
rect 16807 6613 16819 6647
rect 16761 6607 16819 6613
rect 1104 6554 20884 6576
rect 1104 6502 4648 6554
rect 4700 6502 4712 6554
rect 4764 6502 4776 6554
rect 4828 6502 4840 6554
rect 4892 6502 11982 6554
rect 12034 6502 12046 6554
rect 12098 6502 12110 6554
rect 12162 6502 12174 6554
rect 12226 6502 19315 6554
rect 19367 6502 19379 6554
rect 19431 6502 19443 6554
rect 19495 6502 19507 6554
rect 19559 6502 20884 6554
rect 1104 6480 20884 6502
rect 1535 6443 1593 6449
rect 1535 6409 1547 6443
rect 1581 6440 1593 6443
rect 2958 6440 2964 6452
rect 1581 6412 2964 6440
rect 1581 6409 1593 6412
rect 1535 6403 1593 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3326 6440 3332 6452
rect 3287 6412 3332 6440
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 5445 6443 5503 6449
rect 5445 6409 5457 6443
rect 5491 6440 5503 6443
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5491 6412 5825 6440
rect 5491 6409 5503 6412
rect 5445 6403 5503 6409
rect 5813 6409 5825 6412
rect 5859 6440 5871 6443
rect 6638 6440 6644 6452
rect 5859 6412 6644 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 8573 6443 8631 6449
rect 8573 6409 8585 6443
rect 8619 6440 8631 6443
rect 8662 6440 8668 6452
rect 8619 6412 8668 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 8904 6412 9873 6440
rect 8904 6400 8910 6412
rect 9861 6409 9873 6412
rect 9907 6409 9919 6443
rect 13446 6440 13452 6452
rect 13407 6412 13452 6440
rect 9861 6403 9919 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15344 6412 16221 6440
rect 15344 6400 15350 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 16209 6403 16267 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18509 6443 18567 6449
rect 18509 6440 18521 6443
rect 18012 6412 18521 6440
rect 18012 6400 18018 6412
rect 18509 6409 18521 6412
rect 18555 6440 18567 6443
rect 18782 6440 18788 6452
rect 18555 6412 18788 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18782 6400 18788 6412
rect 18840 6400 18846 6452
rect 3234 6332 3240 6384
rect 3292 6372 3298 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 3292 6344 6193 6372
rect 3292 6332 3298 6344
rect 6181 6341 6193 6344
rect 6227 6372 6239 6375
rect 7006 6372 7012 6384
rect 6227 6344 7012 6372
rect 6227 6341 6239 6344
rect 6181 6335 6239 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 7926 6372 7932 6384
rect 7887 6344 7932 6372
rect 7926 6332 7932 6344
rect 7984 6372 7990 6384
rect 11146 6372 11152 6384
rect 7984 6344 9260 6372
rect 11107 6344 11152 6372
rect 7984 6332 7990 6344
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1479 6276 2329 6304
rect 1479 6245 1507 6276
rect 2317 6273 2329 6276
rect 2363 6304 2375 6307
rect 4154 6304 4160 6316
rect 2363 6276 4160 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6304 4583 6307
rect 4982 6304 4988 6316
rect 4571 6276 4988 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7248 6276 7389 6304
rect 7248 6264 7254 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 8938 6304 8944 6316
rect 8899 6276 8944 6304
rect 7377 6267 7435 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9232 6313 9260 6344
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 13354 6332 13360 6384
rect 13412 6372 13418 6384
rect 13817 6375 13875 6381
rect 13817 6372 13829 6375
rect 13412 6344 13829 6372
rect 13412 6332 13418 6344
rect 13817 6341 13829 6344
rect 13863 6341 13875 6375
rect 15930 6372 15936 6384
rect 15891 6344 15936 6372
rect 13817 6335 13875 6341
rect 15930 6332 15936 6344
rect 15988 6332 15994 6384
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 14783 6276 15424 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 1464 6239 1522 6245
rect 1464 6205 1476 6239
rect 1510 6205 1522 6239
rect 2406 6236 2412 6248
rect 2367 6208 2412 6236
rect 1464 6199 1522 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 10413 6239 10471 6245
rect 3743 6208 4154 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1636 6072 1869 6100
rect 1636 6060 1642 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 3712 6100 3740 6199
rect 4126 6168 4154 6208
rect 10413 6205 10425 6239
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 4887 6171 4945 6177
rect 4887 6168 4899 6171
rect 4126 6140 4899 6168
rect 4887 6137 4899 6140
rect 4933 6168 4945 6171
rect 5074 6168 5080 6180
rect 4933 6140 5080 6168
rect 4933 6137 4945 6140
rect 4887 6131 4945 6137
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 6822 6168 6828 6180
rect 5684 6140 6828 6168
rect 5684 6128 5690 6140
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 7466 6128 7472 6180
rect 7524 6168 7530 6180
rect 7524 6140 7617 6168
rect 7524 6128 7530 6140
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9766 6168 9772 6180
rect 9088 6140 9133 6168
rect 9553 6140 9772 6168
rect 9088 6128 9094 6140
rect 4154 6100 4160 6112
rect 2823 6072 3740 6100
rect 4067 6072 4160 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 4154 6060 4160 6072
rect 4212 6100 4218 6112
rect 5994 6100 6000 6112
rect 4212 6072 6000 6100
rect 4212 6060 4218 6072
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 7193 6103 7251 6109
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7484 6100 7512 6128
rect 7239 6072 7512 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9553 6100 9581 6140
rect 9766 6128 9772 6140
rect 9824 6168 9830 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 9824 6140 10241 6168
rect 9824 6128 9830 6140
rect 10229 6137 10241 6140
rect 10275 6168 10287 6171
rect 10428 6168 10456 6199
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 11241 6239 11299 6245
rect 11241 6236 11253 6239
rect 10652 6208 11253 6236
rect 10652 6196 10658 6208
rect 11241 6205 11253 6208
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 11425 6239 11483 6245
rect 11425 6205 11437 6239
rect 11471 6236 11483 6239
rect 11698 6236 11704 6248
rect 11471 6208 11704 6236
rect 11471 6205 11483 6208
rect 11425 6199 11483 6205
rect 10870 6168 10876 6180
rect 10275 6140 10876 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 11256 6168 11284 6199
rect 11698 6196 11704 6208
rect 11756 6236 11762 6248
rect 12526 6236 12532 6248
rect 11756 6208 12296 6236
rect 12487 6208 12532 6236
rect 11756 6196 11762 6208
rect 12066 6168 12072 6180
rect 11256 6140 12072 6168
rect 12066 6128 12072 6140
rect 12124 6128 12130 6180
rect 12268 6112 12296 6208
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12860 6208 13001 6236
rect 12860 6196 12866 6208
rect 12989 6205 13001 6208
rect 13035 6236 13047 6239
rect 13722 6236 13728 6248
rect 13035 6208 13728 6236
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 13722 6196 13728 6208
rect 13780 6236 13786 6248
rect 14826 6236 14832 6248
rect 13780 6208 14832 6236
rect 13780 6196 13786 6208
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 15396 6245 15424 6276
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 15470 6236 15476 6248
rect 15427 6208 15476 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 15470 6196 15476 6208
rect 15528 6236 15534 6248
rect 15948 6236 15976 6332
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6304 17187 6307
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17175 6276 18705 6304
rect 17175 6273 17187 6276
rect 17129 6267 17187 6273
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 19058 6304 19064 6316
rect 18739 6276 19064 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 19058 6264 19064 6276
rect 19116 6304 19122 6316
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19116 6276 19993 6304
rect 19116 6264 19122 6276
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 19981 6267 20039 6273
rect 15528 6208 15976 6236
rect 15528 6196 15534 6208
rect 15565 6171 15623 6177
rect 15565 6137 15577 6171
rect 15611 6168 15623 6171
rect 16298 6168 16304 6180
rect 15611 6140 16304 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 16298 6128 16304 6140
rect 16356 6128 16362 6180
rect 16482 6168 16488 6180
rect 16443 6140 16488 6168
rect 16482 6128 16488 6140
rect 16540 6128 16546 6180
rect 16586 6171 16644 6177
rect 16586 6137 16598 6171
rect 16632 6168 16644 6171
rect 16758 6168 16764 6180
rect 16632 6140 16764 6168
rect 16632 6137 16644 6140
rect 16586 6131 16644 6137
rect 16758 6128 16764 6140
rect 16816 6168 16822 6180
rect 17954 6168 17960 6180
rect 16816 6140 17960 6168
rect 16816 6128 16822 6140
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 18785 6171 18843 6177
rect 18785 6137 18797 6171
rect 18831 6168 18843 6171
rect 18966 6168 18972 6180
rect 18831 6140 18972 6168
rect 18831 6137 18843 6140
rect 18785 6131 18843 6137
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 19334 6168 19340 6180
rect 19295 6140 19340 6168
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 8996 6072 9581 6100
rect 8996 6060 9002 6072
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11756 6072 11805 6100
rect 11756 6060 11762 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 11793 6063 11851 6069
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 12400 6072 12541 6100
rect 12400 6060 12406 6072
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 12529 6063 12587 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 19610 6100 19616 6112
rect 19571 6072 19616 6100
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 1104 6010 20884 6032
rect 1104 5958 8315 6010
rect 8367 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 15648 6010
rect 15700 5958 15712 6010
rect 15764 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 20884 6010
rect 1104 5936 20884 5958
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3108 5868 3433 5896
rect 3108 5856 3114 5868
rect 3421 5865 3433 5868
rect 3467 5896 3479 5899
rect 3694 5896 3700 5908
rect 3467 5868 3700 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3694 5856 3700 5868
rect 3752 5856 3758 5908
rect 3878 5896 3884 5908
rect 3839 5868 3884 5896
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 5500 5868 6101 5896
rect 5500 5856 5506 5868
rect 6089 5865 6101 5868
rect 6135 5896 6147 5899
rect 6178 5896 6184 5908
rect 6135 5868 6184 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 6546 5856 6552 5868
rect 6604 5896 6610 5908
rect 6604 5868 6776 5896
rect 6604 5856 6610 5868
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 2961 5831 3019 5837
rect 2961 5828 2973 5831
rect 2464 5800 2973 5828
rect 2464 5788 2470 5800
rect 2961 5797 2973 5800
rect 3007 5828 3019 5831
rect 3786 5828 3792 5840
rect 3007 5800 3792 5828
rect 3007 5797 3019 5800
rect 2961 5791 3019 5797
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 2222 5760 2228 5772
rect 2183 5732 2228 5760
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 2774 5760 2780 5772
rect 2735 5732 2780 5760
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 3896 5760 3924 5856
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 4982 5828 4988 5840
rect 4847 5800 4988 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 6748 5837 6776 5868
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 8260 5868 8493 5896
rect 8260 5856 8266 5868
rect 8481 5865 8493 5868
rect 8527 5896 8539 5899
rect 8846 5896 8852 5908
rect 8527 5868 8852 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9030 5896 9036 5908
rect 8991 5868 9036 5896
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 9769 5899 9827 5905
rect 9769 5896 9781 5899
rect 9364 5868 9781 5896
rect 9364 5856 9370 5868
rect 9769 5865 9781 5868
rect 9815 5865 9827 5899
rect 9769 5859 9827 5865
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 10965 5899 11023 5905
rect 10965 5896 10977 5899
rect 10928 5868 10977 5896
rect 10928 5856 10934 5868
rect 10965 5865 10977 5868
rect 11011 5865 11023 5899
rect 11422 5896 11428 5908
rect 11383 5868 11428 5896
rect 10965 5859 11023 5865
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13538 5896 13544 5908
rect 13499 5868 13544 5896
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14918 5856 14924 5908
rect 14976 5896 14982 5908
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14976 5868 15025 5896
rect 14976 5856 14982 5868
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 15013 5859 15071 5865
rect 15933 5899 15991 5905
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 16114 5896 16120 5908
rect 15979 5868 16120 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 16853 5899 16911 5905
rect 16853 5896 16865 5899
rect 16356 5868 16865 5896
rect 16356 5856 16362 5868
rect 16853 5865 16865 5868
rect 16899 5896 16911 5899
rect 17954 5896 17960 5908
rect 16899 5868 17080 5896
rect 17915 5868 17960 5896
rect 16899 5865 16911 5868
rect 16853 5859 16911 5865
rect 6733 5831 6791 5837
rect 6733 5797 6745 5831
rect 6779 5797 6791 5831
rect 6733 5791 6791 5797
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 6880 5800 6925 5828
rect 8220 5800 11376 5828
rect 6880 5788 6886 5800
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3896 5732 4077 5760
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4246 5760 4252 5772
rect 4111 5732 4252 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4522 5760 4528 5772
rect 4483 5732 4528 5760
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 5696 5763 5754 5769
rect 5696 5729 5708 5763
rect 5742 5760 5754 5763
rect 5742 5732 6040 5760
rect 5742 5729 5754 5732
rect 5696 5723 5754 5729
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 3786 5692 3792 5704
rect 3660 5664 3792 5692
rect 3660 5652 3666 5664
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 5810 5692 5816 5704
rect 5782 5652 5816 5692
rect 5868 5652 5874 5704
rect 6012 5692 6040 5732
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8220 5769 8248 5800
rect 11348 5772 11376 5800
rect 12066 5788 12072 5840
rect 12124 5828 12130 5840
rect 13081 5831 13139 5837
rect 13081 5828 13093 5831
rect 12124 5800 13093 5828
rect 12124 5788 12130 5800
rect 13081 5797 13093 5800
rect 13127 5828 13139 5831
rect 13127 5800 13814 5828
rect 13127 5797 13139 5800
rect 13081 5791 13139 5797
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7800 5732 8217 5760
rect 7800 5720 7806 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8352 5732 8401 5760
rect 8352 5720 8358 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 9122 5760 9128 5772
rect 8435 5732 9128 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9548 5732 9689 5760
rect 9548 5720 9554 5732
rect 9677 5729 9689 5732
rect 9723 5760 9735 5763
rect 9766 5760 9772 5772
rect 9723 5732 9772 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 11330 5760 11336 5772
rect 11243 5732 11336 5760
rect 10137 5723 10195 5729
rect 6086 5692 6092 5704
rect 5999 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5692 6150 5704
rect 6730 5692 6736 5704
rect 6144 5664 6736 5692
rect 6144 5652 6150 5664
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 6972 5664 8033 5692
rect 6972 5652 6978 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 10152 5692 10180 5723
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 11606 5760 11612 5772
rect 11480 5732 11612 5760
rect 11480 5720 11486 5732
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 11756 5732 12173 5760
rect 11756 5720 11762 5732
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 13262 5760 13268 5772
rect 13223 5732 13268 5760
rect 12161 5723 12219 5729
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 13786 5760 13814 5800
rect 14458 5788 14464 5840
rect 14516 5828 14522 5840
rect 15289 5831 15347 5837
rect 15289 5828 15301 5831
rect 14516 5800 15301 5828
rect 14516 5788 14522 5800
rect 15289 5797 15301 5800
rect 15335 5797 15347 5831
rect 15289 5791 15347 5797
rect 16485 5831 16543 5837
rect 16485 5797 16497 5831
rect 16531 5828 16543 5831
rect 16758 5828 16764 5840
rect 16531 5800 16764 5828
rect 16531 5797 16543 5800
rect 16485 5791 16543 5797
rect 16758 5788 16764 5800
rect 16816 5788 16822 5840
rect 17052 5769 17080 5868
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18233 5899 18291 5905
rect 18233 5896 18245 5899
rect 18196 5868 18245 5896
rect 18196 5856 18202 5868
rect 18233 5865 18245 5868
rect 18279 5865 18291 5899
rect 18233 5859 18291 5865
rect 17402 5837 17408 5840
rect 17399 5828 17408 5837
rect 17315 5800 17408 5828
rect 17399 5791 17408 5800
rect 17460 5828 17466 5840
rect 17862 5828 17868 5840
rect 17460 5800 17868 5828
rect 17402 5788 17408 5791
rect 17460 5788 17466 5800
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 18969 5831 19027 5837
rect 18969 5797 18981 5831
rect 19015 5828 19027 5831
rect 19150 5828 19156 5840
rect 19015 5800 19156 5828
rect 19015 5797 19027 5800
rect 18969 5791 19027 5797
rect 19150 5788 19156 5800
rect 19208 5788 19214 5840
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 13786 5732 14105 5760
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 12250 5692 12256 5704
rect 8904 5664 10180 5692
rect 12163 5664 12256 5692
rect 8904 5652 8910 5664
rect 12250 5652 12256 5664
rect 12308 5692 12314 5704
rect 13998 5692 14004 5704
rect 12308 5664 14004 5692
rect 12308 5652 12314 5664
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15252 5664 15669 5692
rect 15252 5652 15258 5664
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 18874 5692 18880 5704
rect 18835 5664 18880 5692
rect 15657 5655 15715 5661
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 19058 5652 19064 5704
rect 19116 5692 19122 5704
rect 19334 5692 19340 5704
rect 19116 5664 19340 5692
rect 19116 5652 19122 5664
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 1670 5584 1676 5636
rect 1728 5624 1734 5636
rect 5445 5627 5503 5633
rect 5445 5624 5457 5627
rect 1728 5596 5457 5624
rect 1728 5584 1734 5596
rect 5445 5593 5457 5596
rect 5491 5593 5503 5627
rect 5445 5587 5503 5593
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2314 5556 2320 5568
rect 1995 5528 2320 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2314 5516 2320 5528
rect 2372 5516 2378 5568
rect 5782 5565 5810 5652
rect 7282 5624 7288 5636
rect 7243 5596 7288 5624
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 11606 5624 11612 5636
rect 7386 5596 11612 5624
rect 5767 5559 5825 5565
rect 5767 5525 5779 5559
rect 5813 5525 5825 5559
rect 5767 5519 5825 5525
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 7386 5556 7414 5596
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 14826 5584 14832 5636
rect 14884 5624 14890 5636
rect 15565 5627 15623 5633
rect 15565 5624 15577 5627
rect 14884 5596 15577 5624
rect 14884 5584 14890 5596
rect 15565 5593 15577 5596
rect 15611 5593 15623 5627
rect 15565 5587 15623 5593
rect 7650 5556 7656 5568
rect 6052 5528 7414 5556
rect 7611 5528 7656 5556
rect 6052 5516 6058 5528
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15454 5559 15512 5565
rect 15454 5525 15466 5559
rect 15500 5556 15512 5559
rect 16022 5556 16028 5568
rect 15500 5528 16028 5556
rect 15500 5525 15512 5528
rect 15454 5519 15512 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5556 18751 5559
rect 18966 5556 18972 5568
rect 18739 5528 18972 5556
rect 18739 5525 18751 5528
rect 18693 5519 18751 5525
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 1104 5466 20884 5488
rect 1104 5414 4648 5466
rect 4700 5414 4712 5466
rect 4764 5414 4776 5466
rect 4828 5414 4840 5466
rect 4892 5414 11982 5466
rect 12034 5414 12046 5466
rect 12098 5414 12110 5466
rect 12162 5414 12174 5466
rect 12226 5414 19315 5466
rect 19367 5414 19379 5466
rect 19431 5414 19443 5466
rect 19495 5414 19507 5466
rect 19559 5414 20884 5466
rect 1104 5392 20884 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 2961 5355 3019 5361
rect 2961 5352 2973 5355
rect 2832 5324 2973 5352
rect 2832 5312 2838 5324
rect 2961 5321 2973 5324
rect 3007 5352 3019 5355
rect 4522 5352 4528 5364
rect 3007 5324 4528 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5352 4951 5355
rect 5074 5352 5080 5364
rect 4939 5324 5080 5352
rect 4939 5321 4951 5324
rect 4893 5315 4951 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 8938 5352 8944 5364
rect 6472 5324 8944 5352
rect 1946 5284 1952 5296
rect 1872 5256 1952 5284
rect 1872 5157 1900 5256
rect 1946 5244 1952 5256
rect 2004 5244 2010 5296
rect 6472 5284 6500 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9824 5324 10057 5352
rect 9824 5312 9830 5324
rect 10045 5321 10057 5324
rect 10091 5352 10103 5355
rect 10502 5352 10508 5364
rect 10091 5324 10508 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 10686 5352 10692 5364
rect 10647 5324 10692 5352
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11388 5324 12173 5352
rect 11388 5312 11394 5324
rect 12161 5321 12173 5324
rect 12207 5352 12219 5355
rect 12342 5352 12348 5364
rect 12207 5324 12348 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12575 5355 12633 5361
rect 12575 5321 12587 5355
rect 12621 5352 12633 5355
rect 14182 5352 14188 5364
rect 12621 5324 14188 5352
rect 12621 5321 12633 5324
rect 12575 5315 12633 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14458 5352 14464 5364
rect 14419 5324 14464 5352
rect 14458 5312 14464 5324
rect 14516 5352 14522 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 14516 5324 15117 5352
rect 14516 5312 14522 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 15344 5324 16865 5352
rect 15344 5312 15350 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 18966 5352 18972 5364
rect 18927 5324 18972 5352
rect 16853 5315 16911 5321
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 2608 5256 6500 5284
rect 2608 5225 2636 5256
rect 6546 5244 6552 5296
rect 6604 5284 6610 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 6604 5256 6653 5284
rect 6604 5244 6610 5256
rect 6641 5253 6653 5256
rect 6687 5284 6699 5287
rect 6822 5284 6828 5296
rect 6687 5256 6828 5284
rect 6687 5253 6699 5256
rect 6641 5247 6699 5253
rect 6822 5244 6828 5256
rect 6880 5284 6886 5296
rect 6880 5256 7604 5284
rect 6880 5244 6886 5256
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 3602 5216 3608 5228
rect 2593 5179 2651 5185
rect 3436 5188 3608 5216
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5117 2007 5151
rect 1949 5111 2007 5117
rect 2133 5151 2191 5157
rect 2133 5117 2145 5151
rect 2179 5148 2191 5151
rect 2314 5148 2320 5160
rect 2179 5120 2320 5148
rect 2179 5117 2191 5120
rect 2133 5111 2191 5117
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 1964 5080 1992 5111
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 3436 5157 3464 5188
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4522 5216 4528 5228
rect 4120 5188 4528 5216
rect 4120 5176 4126 5188
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5166 5216 5172 5228
rect 5031 5188 5172 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6914 5216 6920 5228
rect 6052 5188 6920 5216
rect 6052 5176 6058 5188
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7282 5216 7288 5228
rect 7243 5188 7288 5216
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 2464 5120 3341 5148
rect 2464 5108 2470 5120
rect 3329 5117 3341 5120
rect 3375 5148 3387 5151
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 3375 5120 3433 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3421 5117 3433 5120
rect 3467 5117 3479 5151
rect 3421 5111 3479 5117
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5117 3571 5151
rect 3694 5148 3700 5160
rect 3655 5120 3700 5148
rect 3513 5111 3571 5117
rect 2774 5080 2780 5092
rect 1811 5052 2780 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 3528 5080 3556 5111
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6730 5148 6736 5160
rect 6319 5120 6736 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 3786 5080 3792 5092
rect 3528 5052 3792 5080
rect 3786 5040 3792 5052
rect 3844 5040 3850 5092
rect 5074 5040 5080 5092
rect 5132 5080 5138 5092
rect 5306 5083 5364 5089
rect 5306 5080 5318 5083
rect 5132 5052 5318 5080
rect 5132 5040 5138 5052
rect 5306 5049 5318 5052
rect 5352 5049 5364 5083
rect 5306 5043 5364 5049
rect 7009 5083 7067 5089
rect 7009 5049 7021 5083
rect 7055 5049 7067 5083
rect 7576 5080 7604 5256
rect 8202 5244 8208 5296
rect 8260 5284 8266 5296
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8260 5256 9045 5284
rect 8260 5244 8266 5256
rect 9033 5253 9045 5256
rect 9079 5284 9091 5287
rect 9398 5284 9404 5296
rect 9079 5256 9404 5284
rect 9079 5253 9091 5256
rect 9033 5247 9091 5253
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 11425 5287 11483 5293
rect 11425 5253 11437 5287
rect 11471 5284 11483 5287
rect 11790 5284 11796 5296
rect 11471 5256 11796 5284
rect 11471 5253 11483 5256
rect 11425 5247 11483 5253
rect 11790 5244 11796 5256
rect 11848 5284 11854 5296
rect 16022 5284 16028 5296
rect 11848 5256 14228 5284
rect 15983 5256 16028 5284
rect 11848 5244 11854 5256
rect 7834 5216 7840 5228
rect 7795 5188 7840 5216
rect 7834 5176 7840 5188
rect 7892 5216 7898 5228
rect 8294 5216 8300 5228
rect 7892 5188 8300 5216
rect 7892 5176 7898 5188
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 9122 5216 9128 5228
rect 8527 5188 9128 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 10962 5216 10968 5228
rect 10919 5188 10968 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 10962 5176 10968 5188
rect 11020 5216 11026 5228
rect 12066 5216 12072 5228
rect 11020 5188 12072 5216
rect 11020 5176 11026 5188
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 13262 5216 13268 5228
rect 12400 5188 13268 5216
rect 12400 5176 12406 5188
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 13412 5188 13553 5216
rect 13412 5176 13418 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7800 5120 8217 5148
rect 7800 5108 7806 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 11606 5108 11612 5160
rect 11664 5148 11670 5160
rect 12504 5151 12562 5157
rect 12504 5148 12516 5151
rect 11664 5120 12516 5148
rect 11664 5108 11670 5120
rect 12504 5117 12516 5120
rect 12550 5148 12562 5151
rect 12550 5120 13032 5148
rect 12550 5117 12562 5120
rect 12504 5111 12562 5117
rect 8573 5083 8631 5089
rect 8573 5080 8585 5083
rect 7576 5052 8585 5080
rect 7009 5043 7067 5049
rect 8573 5049 8585 5052
rect 8619 5080 8631 5083
rect 8662 5080 8668 5092
rect 8619 5052 8668 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 3476 4984 3893 5012
rect 3476 4972 3482 4984
rect 3881 4981 3893 4984
rect 3927 4981 3939 5015
rect 3881 4975 3939 4981
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 7024 5012 7052 5043
rect 8662 5040 8668 5052
rect 8720 5040 8726 5092
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 8904 5052 9689 5080
rect 8904 5040 8910 5052
rect 9677 5049 9689 5052
rect 9723 5049 9735 5083
rect 9677 5043 9735 5049
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 11020 5052 11065 5080
rect 11020 5040 11026 5052
rect 7190 5012 7196 5024
rect 5951 4984 7196 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 7190 4972 7196 4984
rect 7248 5012 7254 5024
rect 7558 5012 7564 5024
rect 7248 4984 7564 5012
rect 7248 4972 7254 4984
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 13004 5021 13032 5120
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 14200 5089 14228 5256
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 18874 5244 18880 5296
rect 18932 5284 18938 5296
rect 19613 5287 19671 5293
rect 19613 5284 19625 5287
rect 18932 5256 19625 5284
rect 18932 5244 18938 5256
rect 19613 5253 19625 5256
rect 19659 5253 19671 5287
rect 19613 5247 19671 5253
rect 16574 5216 16580 5228
rect 15028 5188 16580 5216
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 15028 5157 15056 5188
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5216 18107 5219
rect 18138 5216 18144 5228
rect 18095 5188 18144 5216
rect 18095 5185 18107 5188
rect 18049 5179 18107 5185
rect 18138 5176 18144 5188
rect 18196 5176 18202 5228
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14976 5120 15025 5148
rect 14976 5108 14982 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 15102 5108 15108 5160
rect 15160 5148 15166 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15160 5120 15761 5148
rect 15160 5108 15166 5120
rect 15749 5117 15761 5120
rect 15795 5148 15807 5151
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 15795 5120 16773 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 16761 5117 16773 5120
rect 16807 5148 16819 5151
rect 17497 5151 17555 5157
rect 17497 5148 17509 5151
rect 16807 5120 17509 5148
rect 16807 5117 16819 5120
rect 16761 5111 16819 5117
rect 17497 5117 17509 5120
rect 17543 5148 17555 5151
rect 19426 5148 19432 5160
rect 17543 5120 19432 5148
rect 17543 5117 17555 5120
rect 17497 5111 17555 5117
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 14185 5083 14243 5089
rect 13688 5052 13733 5080
rect 13688 5040 13694 5052
rect 14185 5049 14197 5083
rect 14231 5080 14243 5083
rect 14734 5080 14740 5092
rect 14231 5052 14740 5080
rect 14231 5049 14243 5052
rect 14185 5043 14243 5049
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 16393 5083 16451 5089
rect 16393 5080 16405 5083
rect 15252 5052 16405 5080
rect 15252 5040 15258 5052
rect 16393 5049 16405 5052
rect 16439 5049 16451 5083
rect 16574 5080 16580 5092
rect 16535 5052 16580 5080
rect 16393 5043 16451 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11756 4984 11805 5012
rect 11756 4972 11762 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 11793 4975 11851 4981
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 14274 5012 14280 5024
rect 13035 4984 14280 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 14826 5012 14832 5024
rect 14787 4984 14832 5012
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 17862 5012 17868 5024
rect 17775 4984 17868 5012
rect 17862 4972 17868 4984
rect 17920 5012 17926 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 17920 4984 18429 5012
rect 17920 4972 17926 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 19242 5012 19248 5024
rect 19203 4984 19248 5012
rect 18417 4975 18475 4981
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 1104 4922 20884 4944
rect 1104 4870 8315 4922
rect 8367 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 15648 4922
rect 15700 4870 15712 4922
rect 15764 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 20884 4922
rect 1104 4848 20884 4870
rect 1535 4811 1593 4817
rect 1535 4777 1547 4811
rect 1581 4808 1593 4811
rect 1670 4808 1676 4820
rect 1581 4780 1676 4808
rect 1581 4777 1593 4780
rect 1535 4771 1593 4777
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 2866 4808 2872 4820
rect 2740 4780 2872 4808
rect 2740 4768 2746 4780
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3752 4780 3801 4808
rect 3752 4768 3758 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 5074 4808 5080 4820
rect 4028 4780 5080 4808
rect 4028 4768 4034 4780
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 5442 4808 5448 4820
rect 5355 4780 5448 4808
rect 5442 4768 5448 4780
rect 5500 4808 5506 4820
rect 5626 4808 5632 4820
rect 5500 4780 5632 4808
rect 5500 4768 5506 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6546 4808 6552 4820
rect 6507 4780 6552 4808
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 7190 4808 7196 4820
rect 7151 4780 7196 4808
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 7650 4808 7656 4820
rect 7300 4780 7656 4808
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1872 4672 1900 4768
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 3142 4740 3148 4752
rect 2455 4712 3004 4740
rect 3103 4712 3148 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 2038 4672 2044 4684
rect 1510 4644 2044 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2556 4675 2614 4681
rect 2556 4641 2568 4675
rect 2602 4672 2614 4675
rect 2682 4672 2688 4684
rect 2602 4644 2688 4672
rect 2602 4641 2614 4644
rect 2556 4635 2614 4641
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2976 4604 3004 4712
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3804 4712 4200 4740
rect 3804 4684 3832 4712
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 3513 4675 3571 4681
rect 3513 4672 3525 4675
rect 3476 4644 3525 4672
rect 3476 4632 3482 4644
rect 3513 4641 3525 4644
rect 3559 4672 3571 4675
rect 3786 4672 3792 4684
rect 3559 4644 3792 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 4062 4672 4068 4684
rect 4023 4644 4068 4672
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4172 4681 4200 4712
rect 4246 4700 4252 4752
rect 4304 4740 4310 4752
rect 4801 4743 4859 4749
rect 4801 4740 4813 4743
rect 4304 4712 4813 4740
rect 4304 4700 4310 4712
rect 4801 4709 4813 4712
rect 4847 4740 4859 4743
rect 5534 4740 5540 4752
rect 4847 4712 5540 4740
rect 4847 4709 4859 4712
rect 4801 4703 4859 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 5991 4743 6049 4749
rect 5991 4709 6003 4743
rect 6037 4740 6049 4743
rect 6454 4740 6460 4752
rect 6037 4712 6460 4740
rect 6037 4709 6049 4712
rect 5991 4703 6049 4709
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4641 4215 4675
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4157 4635 4215 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 5718 4672 5724 4684
rect 5675 4644 5724 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 5718 4632 5724 4644
rect 5776 4672 5782 4684
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 5776 4644 6837 4672
rect 5776 4632 5782 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 6825 4635 6883 4641
rect 3970 4604 3976 4616
rect 2976 4576 3976 4604
rect 2777 4567 2835 4573
rect 2314 4536 2320 4548
rect 2275 4508 2320 4536
rect 2314 4496 2320 4508
rect 2372 4496 2378 4548
rect 2792 4536 2820 4567
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 7300 4604 7328 4780
rect 7650 4768 7656 4780
rect 7708 4808 7714 4820
rect 7926 4808 7932 4820
rect 7708 4780 7932 4808
rect 7708 4768 7714 4780
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 8662 4808 8668 4820
rect 8527 4780 8668 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 10962 4808 10968 4820
rect 10919 4780 10968 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 10962 4768 10968 4780
rect 11020 4808 11026 4820
rect 11698 4808 11704 4820
rect 11020 4780 11704 4808
rect 11020 4768 11026 4780
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 15102 4808 15108 4820
rect 15063 4780 15108 4808
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15528 4780 15945 4808
rect 15528 4768 15534 4780
rect 15933 4777 15945 4780
rect 15979 4808 15991 4811
rect 16206 4808 16212 4820
rect 15979 4780 16212 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 16574 4808 16580 4820
rect 16535 4780 16580 4808
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 18325 4811 18383 4817
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 19242 4808 19248 4820
rect 18371 4780 19248 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 7558 4740 7564 4752
rect 7519 4712 7564 4740
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 7834 4700 7840 4752
rect 7892 4740 7898 4752
rect 8113 4743 8171 4749
rect 8113 4740 8125 4743
rect 7892 4712 8125 4740
rect 7892 4700 7898 4712
rect 8113 4709 8125 4712
rect 8159 4740 8171 4743
rect 8202 4740 8208 4752
rect 8159 4712 8208 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 8938 4700 8944 4752
rect 8996 4740 9002 4752
rect 9677 4743 9735 4749
rect 9677 4740 9689 4743
rect 8996 4712 9689 4740
rect 8996 4700 9002 4712
rect 9677 4709 9689 4712
rect 9723 4709 9735 4743
rect 11238 4740 11244 4752
rect 11199 4712 11244 4740
rect 9677 4703 9735 4709
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 11790 4740 11796 4752
rect 11751 4712 11796 4740
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 12983 4743 13041 4749
rect 12983 4709 12995 4743
rect 13029 4740 13041 4743
rect 13446 4740 13452 4752
rect 13029 4712 13452 4740
rect 13029 4709 13041 4712
rect 12983 4703 13041 4709
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 15194 4700 15200 4752
rect 15252 4740 15258 4752
rect 17767 4743 17825 4749
rect 15252 4712 15700 4740
rect 15252 4700 15258 4712
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 9950 4672 9956 4684
rect 9907 4644 9956 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 12492 4644 12633 4672
rect 12492 4632 12498 4644
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 13998 4672 14004 4684
rect 13955 4644 14004 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 13998 4632 14004 4644
rect 14056 4672 14062 4684
rect 15010 4672 15016 4684
rect 14056 4644 15016 4672
rect 14056 4632 14062 4644
rect 15010 4632 15016 4644
rect 15068 4672 15074 4684
rect 15286 4672 15292 4684
rect 15068 4644 15292 4672
rect 15068 4632 15074 4644
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7300 4576 7481 4604
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 11146 4604 11152 4616
rect 7469 4567 7527 4573
rect 7576 4576 10640 4604
rect 11107 4576 11152 4604
rect 2958 4536 2964 4548
rect 2792 4508 2964 4536
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 2498 4468 2504 4480
rect 1728 4440 2504 4468
rect 1728 4428 1734 4440
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 2685 4471 2743 4477
rect 2685 4437 2697 4471
rect 2731 4468 2743 4471
rect 2774 4468 2780 4480
rect 2731 4440 2780 4468
rect 2731 4437 2743 4440
rect 2685 4431 2743 4437
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 7576 4468 7604 4576
rect 7650 4496 7656 4548
rect 7708 4536 7714 4548
rect 9674 4536 9680 4548
rect 7708 4508 9680 4536
rect 7708 4496 7714 4508
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 8754 4468 8760 4480
rect 5500 4440 7604 4468
rect 8715 4440 8760 4468
rect 5500 4428 5506 4440
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 9214 4468 9220 4480
rect 9175 4440 9220 4468
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 9953 4471 10011 4477
rect 9953 4468 9965 4471
rect 9824 4440 9965 4468
rect 9824 4428 9830 4440
rect 9953 4437 9965 4440
rect 9999 4468 10011 4471
rect 10134 4468 10140 4480
rect 9999 4440 10140 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 10612 4468 10640 4576
rect 11146 4564 11152 4576
rect 11204 4604 11210 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 11204 4576 12541 4604
rect 11204 4564 11210 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 14734 4604 14740 4616
rect 14647 4576 14740 4604
rect 12529 4567 12587 4573
rect 14734 4564 14740 4576
rect 14792 4604 14798 4616
rect 15378 4604 15384 4616
rect 14792 4576 15384 4604
rect 14792 4564 14798 4576
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15672 4613 15700 4712
rect 17767 4709 17779 4743
rect 17813 4740 17825 4743
rect 17862 4740 17868 4752
rect 17813 4712 17868 4740
rect 17813 4709 17825 4712
rect 17767 4703 17825 4709
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 18598 4700 18604 4752
rect 18656 4740 18662 4752
rect 19153 4743 19211 4749
rect 19153 4740 19165 4743
rect 18656 4712 19165 4740
rect 18656 4700 18662 4712
rect 19153 4709 19165 4712
rect 19199 4740 19211 4743
rect 20070 4740 20076 4752
rect 19199 4712 20076 4740
rect 19199 4709 19211 4712
rect 19153 4703 19211 4709
rect 20070 4700 20076 4712
rect 20128 4740 20134 4752
rect 21542 4740 21548 4752
rect 20128 4712 21548 4740
rect 20128 4700 20134 4712
rect 21542 4700 21548 4712
rect 21600 4700 21606 4752
rect 19337 4675 19395 4681
rect 19337 4641 19349 4675
rect 19383 4672 19395 4675
rect 19426 4672 19432 4684
rect 19383 4644 19432 4672
rect 19383 4641 19395 4644
rect 19337 4635 19395 4641
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 18138 4604 18144 4616
rect 17451 4576 18144 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 11790 4536 11796 4548
rect 10836 4508 11796 4536
rect 10836 4496 10842 4508
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 14185 4539 14243 4545
rect 14185 4536 14197 4539
rect 13786 4508 14197 4536
rect 12526 4468 12532 4480
rect 10612 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 13538 4468 13544 4480
rect 13499 4440 13544 4468
rect 13538 4428 13544 4440
rect 13596 4468 13602 4480
rect 13786 4468 13814 4508
rect 14185 4505 14197 4508
rect 14231 4505 14243 4539
rect 14185 4499 14243 4505
rect 14826 4496 14832 4548
rect 14884 4536 14890 4548
rect 15565 4539 15623 4545
rect 15565 4536 15577 4539
rect 14884 4508 15577 4536
rect 14884 4496 14890 4508
rect 15565 4505 15577 4508
rect 15611 4536 15623 4539
rect 16022 4536 16028 4548
rect 15611 4508 16028 4536
rect 15611 4505 15623 4508
rect 15565 4499 15623 4505
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 13596 4440 13814 4468
rect 15454 4471 15512 4477
rect 13596 4428 13602 4440
rect 15454 4437 15466 4471
rect 15500 4468 15512 4471
rect 15930 4468 15936 4480
rect 15500 4440 15936 4468
rect 15500 4437 15512 4440
rect 15454 4431 15512 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 16908 4440 17049 4468
rect 16908 4428 16914 4440
rect 17037 4437 17049 4440
rect 17083 4437 17095 4471
rect 17037 4431 17095 4437
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 19429 4471 19487 4477
rect 19429 4468 19441 4471
rect 17184 4440 19441 4468
rect 17184 4428 17190 4440
rect 19429 4437 19441 4440
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 1104 4378 20884 4400
rect 1104 4326 4648 4378
rect 4700 4326 4712 4378
rect 4764 4326 4776 4378
rect 4828 4326 4840 4378
rect 4892 4326 11982 4378
rect 12034 4326 12046 4378
rect 12098 4326 12110 4378
rect 12162 4326 12174 4378
rect 12226 4326 19315 4378
rect 19367 4326 19379 4378
rect 19431 4326 19443 4378
rect 19495 4326 19507 4378
rect 19559 4326 20884 4378
rect 1104 4304 20884 4326
rect 2961 4267 3019 4273
rect 2961 4264 2973 4267
rect 1688 4236 2973 4264
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1688 4137 1716 4236
rect 2961 4233 2973 4236
rect 3007 4264 3019 4267
rect 3007 4236 3740 4264
rect 3007 4233 3019 4236
rect 2961 4227 3019 4233
rect 3142 4196 3148 4208
rect 3103 4168 3148 4196
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 3712 4196 3740 4236
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 3844 4236 4629 4264
rect 3844 4224 3850 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 4617 4227 4675 4233
rect 4861 4236 6561 4264
rect 4062 4196 4068 4208
rect 3712 4168 4068 4196
rect 4062 4156 4068 4168
rect 4120 4156 4126 4208
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 4861 4196 4889 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 8202 4264 8208 4276
rect 7055 4236 8208 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8996 4236 9045 4264
rect 8996 4224 9002 4236
rect 9033 4233 9045 4236
rect 9079 4233 9091 4267
rect 9033 4227 9091 4233
rect 9493 4267 9551 4273
rect 9493 4233 9505 4267
rect 9539 4264 9551 4267
rect 9950 4264 9956 4276
rect 9539 4236 9956 4264
rect 9539 4233 9551 4236
rect 9493 4227 9551 4233
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10560 4236 11554 4264
rect 10560 4224 10566 4236
rect 4488 4168 4889 4196
rect 5077 4199 5135 4205
rect 4488 4156 4494 4168
rect 5077 4165 5089 4199
rect 5123 4196 5135 4199
rect 5258 4196 5264 4208
rect 5123 4168 5264 4196
rect 5123 4165 5135 4168
rect 5077 4159 5135 4165
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 7745 4199 7803 4205
rect 7745 4196 7757 4199
rect 7248 4168 7757 4196
rect 7248 4156 7254 4168
rect 7745 4165 7757 4168
rect 7791 4165 7803 4199
rect 7745 4159 7803 4165
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 10229 4199 10287 4205
rect 10229 4196 10241 4199
rect 9824 4168 10241 4196
rect 9824 4156 9830 4168
rect 10229 4165 10241 4168
rect 10275 4165 10287 4199
rect 10229 4159 10287 4165
rect 11057 4199 11115 4205
rect 11057 4165 11069 4199
rect 11103 4196 11115 4199
rect 11238 4196 11244 4208
rect 11103 4168 11244 4196
rect 11103 4165 11115 4168
rect 11057 4159 11115 4165
rect 11238 4156 11244 4168
rect 11296 4156 11302 4208
rect 11526 4196 11554 4236
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11756 4236 12173 4264
rect 11756 4224 11762 4236
rect 12161 4233 12173 4236
rect 12207 4264 12219 4267
rect 12618 4264 12624 4276
rect 12207 4236 12624 4264
rect 12207 4233 12219 4236
rect 12161 4227 12219 4233
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 15565 4267 15623 4273
rect 15565 4233 15577 4267
rect 15611 4264 15623 4267
rect 15930 4264 15936 4276
rect 15611 4236 15936 4264
rect 15611 4233 15623 4236
rect 15565 4227 15623 4233
rect 15930 4224 15936 4236
rect 15988 4264 15994 4276
rect 17954 4264 17960 4276
rect 15988 4236 17960 4264
rect 15988 4224 15994 4236
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 19150 4264 19156 4276
rect 19111 4236 19156 4264
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19751 4267 19809 4273
rect 19751 4264 19763 4267
rect 19668 4236 19763 4264
rect 19668 4224 19674 4236
rect 19751 4233 19763 4236
rect 19797 4233 19809 4267
rect 20070 4264 20076 4276
rect 20031 4236 20076 4264
rect 19751 4227 19809 4233
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 11526 4168 13860 4196
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1544 4100 1685 4128
rect 1544 4088 1550 4100
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 2188 4100 3801 4128
rect 2188 4088 2194 4100
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 4338 4128 4344 4140
rect 4299 4100 4344 4128
rect 3789 4091 3847 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 5905 4131 5963 4137
rect 5321 4100 5672 4128
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2406 4060 2412 4072
rect 2363 4032 2412 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2866 4060 2872 4072
rect 2823 4032 2872 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4060 3019 4063
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3007 4032 3249 4060
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 3237 4023 3295 4029
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3513 4063 3571 4069
rect 3384 4032 3429 4060
rect 3384 4020 3390 4032
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 3694 4060 3700 4072
rect 3559 4032 3700 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 5321 4060 5349 4100
rect 5644 4072 5672 4100
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6270 4128 6276 4140
rect 5951 4100 6276 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 6840 4100 7481 4128
rect 5442 4060 5448 4072
rect 4126 4032 5349 4060
rect 5403 4032 5448 4060
rect 2222 3952 2228 4004
rect 2280 3992 2286 4004
rect 3602 3992 3608 4004
rect 2280 3964 3608 3992
rect 2280 3952 2286 3964
rect 3602 3952 3608 3964
rect 3660 3992 3666 4004
rect 4126 3992 4154 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5626 4060 5632 4072
rect 5539 4032 5632 4060
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 6840 4069 6868 4100
rect 7469 4097 7481 4100
rect 7515 4128 7527 4131
rect 7650 4128 7656 4140
rect 7515 4100 7656 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 7852 4100 9689 4128
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 3660 3964 4154 3992
rect 3660 3952 3666 3964
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 7852 3992 7880 4100
rect 9677 4097 9689 4100
rect 9723 4128 9735 4131
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 9723 4100 10609 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 11848 4100 12541 4128
rect 11848 4088 11854 4100
rect 12529 4097 12541 4100
rect 12575 4128 12587 4131
rect 12986 4128 12992 4140
rect 12575 4100 12992 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 10928 4032 11161 4060
rect 10928 4020 10934 4032
rect 11149 4029 11161 4032
rect 11195 4060 11207 4063
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11195 4032 11713 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 13832 4060 13860 4168
rect 18248 4168 18368 4196
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14366 4128 14372 4140
rect 13955 4100 14372 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 16776 4100 17877 4128
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 13832 4032 16221 4060
rect 11701 4023 11759 4029
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 5224 3964 7880 3992
rect 8021 3995 8079 4001
rect 5224 3952 5230 3964
rect 8021 3961 8033 3995
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 8113 3995 8171 4001
rect 8113 3961 8125 3995
rect 8159 3961 8171 3995
rect 8662 3992 8668 4004
rect 8575 3964 8668 3992
rect 8113 3955 8171 3961
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4338 3924 4344 3936
rect 3936 3896 4344 3924
rect 3936 3884 3942 3896
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 6273 3927 6331 3933
rect 6273 3893 6285 3927
rect 6319 3924 6331 3927
rect 6454 3924 6460 3936
rect 6319 3896 6460 3924
rect 6319 3893 6331 3896
rect 6273 3887 6331 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7834 3924 7840 3936
rect 7064 3896 7840 3924
rect 7064 3884 7070 3896
rect 7834 3884 7840 3896
rect 7892 3924 7898 3936
rect 8036 3924 8064 3955
rect 7892 3896 8064 3924
rect 8128 3924 8156 3955
rect 8662 3952 8668 3964
rect 8720 3992 8726 4004
rect 9674 3992 9680 4004
rect 8720 3964 9680 3992
rect 8720 3952 8726 3964
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 10134 3992 10140 4004
rect 9815 3964 10140 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 13173 3995 13231 4001
rect 12676 3964 12721 3992
rect 12676 3952 12682 3964
rect 13173 3961 13185 3995
rect 13219 3992 13231 3995
rect 14090 3992 14096 4004
rect 13219 3964 14096 3992
rect 13219 3961 13231 3964
rect 13173 3955 13231 3961
rect 14090 3952 14096 3964
rect 14148 3992 14154 4004
rect 14642 3992 14648 4004
rect 14148 3964 14648 3992
rect 14148 3952 14154 3964
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 16224 3992 16252 4023
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 16776 4069 16804 4100
rect 17865 4097 17877 4100
rect 17911 4128 17923 4131
rect 18248 4128 18276 4168
rect 17911 4100 18276 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16448 4032 16773 4060
rect 16448 4020 16454 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 18230 4060 18236 4072
rect 18191 4032 18236 4060
rect 16761 4023 16819 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18340 4060 18368 4168
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18340 4032 18521 4060
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 19680 4063 19738 4069
rect 19680 4029 19692 4063
rect 19726 4029 19738 4063
rect 19680 4023 19738 4029
rect 16574 3992 16580 4004
rect 16224 3964 16580 3992
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 16945 3995 17003 4001
rect 16945 3961 16957 3995
rect 16991 3992 17003 3995
rect 17310 3992 17316 4004
rect 16991 3964 17316 3992
rect 16991 3961 17003 3964
rect 16945 3955 17003 3961
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 18138 3952 18144 4004
rect 18196 3992 18202 4004
rect 18782 3992 18788 4004
rect 18196 3964 18788 3992
rect 18196 3952 18202 3964
rect 18782 3952 18788 3964
rect 18840 3952 18846 4004
rect 18874 3952 18880 4004
rect 18932 3992 18938 4004
rect 19695 3992 19723 4023
rect 20441 3995 20499 4001
rect 20441 3992 20453 3995
rect 18932 3964 20453 3992
rect 18932 3952 18938 3964
rect 20441 3961 20453 3964
rect 20487 3961 20499 3995
rect 20441 3955 20499 3961
rect 8754 3924 8760 3936
rect 8128 3896 8760 3924
rect 7892 3884 7898 3896
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 9548 3896 11345 3924
rect 9548 3884 9554 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 11333 3887 11391 3893
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 13446 3924 13452 3936
rect 11572 3896 13452 3924
rect 11572 3884 11578 3896
rect 13446 3884 13452 3896
rect 13504 3924 13510 3936
rect 14185 3927 14243 3933
rect 14185 3924 14197 3927
rect 13504 3896 14197 3924
rect 13504 3884 13510 3896
rect 14185 3893 14197 3896
rect 14231 3924 14243 3927
rect 14737 3927 14795 3933
rect 14737 3924 14749 3927
rect 14231 3896 14749 3924
rect 14231 3893 14243 3896
rect 14185 3887 14243 3893
rect 14737 3893 14749 3896
rect 14783 3924 14795 3927
rect 15102 3924 15108 3936
rect 14783 3896 15108 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15289 3927 15347 3933
rect 15289 3893 15301 3927
rect 15335 3924 15347 3927
rect 15470 3924 15476 3936
rect 15335 3896 15476 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 16022 3924 16028 3936
rect 15983 3896 16028 3924
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 16908 3896 17417 3924
rect 16908 3884 16914 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 1104 3834 20884 3856
rect 1104 3782 8315 3834
rect 8367 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 15648 3834
rect 15700 3782 15712 3834
rect 15764 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 20884 3834
rect 1104 3760 20884 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 5166 3720 5172 3732
rect 1443 3692 5172 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5534 3720 5540 3732
rect 5495 3692 5540 3720
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5684 3692 5917 3720
rect 5684 3680 5690 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 6362 3680 6368 3732
rect 6420 3720 6426 3732
rect 7558 3720 7564 3732
rect 6420 3692 7564 3720
rect 6420 3680 6426 3692
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8754 3720 8760 3732
rect 8619 3692 8760 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9306 3720 9312 3732
rect 9263 3692 9312 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10192 3692 10241 3720
rect 10192 3680 10198 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11790 3720 11796 3732
rect 11388 3692 11796 3720
rect 11388 3680 11394 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 12621 3723 12679 3729
rect 12621 3720 12633 3723
rect 12400 3692 12633 3720
rect 12400 3680 12406 3692
rect 12621 3689 12633 3692
rect 12667 3689 12679 3723
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12621 3683 12679 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 15010 3720 15016 3732
rect 14971 3692 15016 3720
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 16390 3720 16396 3732
rect 16351 3692 16396 3720
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 18046 3720 18052 3732
rect 16540 3692 18052 3720
rect 16540 3680 16546 3692
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 18230 3720 18236 3732
rect 18191 3692 18236 3720
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 18782 3720 18788 3732
rect 18739 3692 18788 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 2317 3655 2375 3661
rect 2317 3621 2329 3655
rect 2363 3652 2375 3655
rect 2774 3652 2780 3664
rect 2363 3624 2780 3652
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 3145 3655 3203 3661
rect 3145 3621 3157 3655
rect 3191 3652 3203 3655
rect 3510 3652 3516 3664
rect 3191 3624 3516 3652
rect 3191 3621 3203 3624
rect 3145 3615 3203 3621
rect 3510 3612 3516 3624
rect 3568 3652 3574 3664
rect 5442 3652 5448 3664
rect 3568 3624 5448 3652
rect 3568 3612 3574 3624
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2406 3584 2412 3596
rect 1995 3556 2412 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 3786 3584 3792 3596
rect 2731 3556 3792 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2700 3516 2728 3547
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 4062 3584 4068 3596
rect 3927 3556 4068 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4062 3544 4068 3556
rect 4120 3584 4126 3596
rect 4816 3593 4844 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 6178 3652 6184 3664
rect 6139 3624 6184 3652
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 6270 3612 6276 3664
rect 6328 3652 6334 3664
rect 6328 3624 6373 3652
rect 6328 3612 6334 3624
rect 7834 3612 7840 3664
rect 7892 3652 7898 3664
rect 7974 3655 8032 3661
rect 7974 3652 7986 3655
rect 7892 3624 7986 3652
rect 7892 3612 7898 3624
rect 7974 3621 7986 3624
rect 8020 3621 8032 3655
rect 11235 3655 11293 3661
rect 7974 3615 8032 3621
rect 8128 3624 10916 3652
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4120 3556 4261 3584
rect 4120 3544 4126 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 5350 3584 5356 3596
rect 5123 3556 5356 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 7374 3584 7380 3596
rect 6871 3556 7380 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 7374 3544 7380 3556
rect 7432 3584 7438 3596
rect 8128 3584 8156 3624
rect 7432 3556 8156 3584
rect 9677 3587 9735 3593
rect 7432 3544 7438 3556
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 10778 3584 10784 3596
rect 9723 3556 10784 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 10888 3584 10916 3624
rect 11235 3621 11247 3655
rect 11281 3652 11293 3655
rect 11514 3652 11520 3664
rect 11281 3624 11520 3652
rect 11281 3621 11293 3624
rect 11235 3615 11293 3621
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 13538 3652 13544 3664
rect 13499 3624 13544 3652
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 14090 3652 14096 3664
rect 14051 3624 14096 3652
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 14737 3655 14795 3661
rect 14737 3621 14749 3655
rect 14783 3652 14795 3655
rect 15194 3652 15200 3664
rect 14783 3624 15200 3652
rect 14783 3621 14795 3624
rect 14737 3615 14795 3621
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 15378 3652 15384 3664
rect 15339 3624 15384 3652
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 16025 3655 16083 3661
rect 15528 3624 15573 3652
rect 15528 3612 15534 3624
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16942 3652 16948 3664
rect 16071 3624 16948 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16942 3612 16948 3624
rect 17000 3612 17006 3664
rect 17286 3655 17344 3661
rect 17286 3652 17298 3655
rect 17230 3624 17298 3652
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 10888 3556 12081 3584
rect 12069 3553 12081 3556
rect 12115 3553 12127 3587
rect 12069 3547 12127 3553
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 16632 3556 16681 3584
rect 16632 3544 16638 3556
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 17230 3584 17258 3624
rect 17286 3621 17298 3624
rect 17332 3621 17344 3655
rect 18966 3652 18972 3664
rect 17286 3615 17344 3621
rect 18708 3624 18972 3652
rect 16908 3556 17258 3584
rect 17957 3587 18015 3593
rect 16908 3544 16914 3556
rect 17957 3553 17969 3587
rect 18003 3584 18015 3587
rect 18708 3584 18736 3624
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 18003 3556 18736 3584
rect 18003 3553 18015 3556
rect 17957 3547 18015 3553
rect 1728 3488 2728 3516
rect 5261 3519 5319 3525
rect 1728 3476 1734 3488
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 6914 3516 6920 3528
rect 5307 3488 6920 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 7156 3488 7665 3516
rect 7156 3476 7162 3488
rect 7653 3485 7665 3488
rect 7699 3516 7711 3519
rect 8110 3516 8116 3528
rect 7699 3488 8116 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10704 3488 10885 3516
rect 2501 3451 2559 3457
rect 2501 3417 2513 3451
rect 2547 3448 2559 3451
rect 2590 3448 2596 3460
rect 2547 3420 2596 3448
rect 2547 3417 2559 3420
rect 2501 3411 2559 3417
rect 2590 3408 2596 3420
rect 2648 3448 2654 3460
rect 3050 3448 3056 3460
rect 2648 3420 3056 3448
rect 2648 3408 2654 3420
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 3142 3408 3148 3460
rect 3200 3448 3206 3460
rect 7742 3448 7748 3460
rect 3200 3420 7748 3448
rect 3200 3408 3206 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 10704 3392 10732 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 12768 3488 13461 3516
rect 12768 3476 12774 3488
rect 13449 3485 13461 3488
rect 13495 3516 13507 3519
rect 14826 3516 14832 3528
rect 13495 3488 14832 3516
rect 13495 3485 13507 3488
rect 13449 3479 13507 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17310 3516 17316 3528
rect 17083 3488 17316 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3485 18935 3519
rect 19150 3516 19156 3528
rect 19111 3488 19156 3516
rect 18877 3479 18935 3485
rect 10778 3408 10784 3460
rect 10836 3448 10842 3460
rect 12618 3448 12624 3460
rect 10836 3420 12624 3448
rect 10836 3408 10842 3420
rect 12618 3408 12624 3420
rect 12676 3448 12682 3460
rect 16666 3448 16672 3460
rect 12676 3420 16672 3448
rect 12676 3408 12682 3420
rect 16666 3408 16672 3420
rect 16724 3448 16730 3460
rect 16724 3420 17080 3448
rect 16724 3408 16730 3420
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3326 3380 3332 3392
rect 2832 3352 3332 3380
rect 2832 3340 2838 3352
rect 3326 3340 3332 3352
rect 3384 3380 3390 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3384 3352 3433 3380
rect 3384 3340 3390 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 3421 3343 3479 3349
rect 7377 3383 7435 3389
rect 7377 3349 7389 3383
rect 7423 3380 7435 3383
rect 7466 3380 7472 3392
rect 7423 3352 7472 3380
rect 7423 3349 7435 3352
rect 7377 3343 7435 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 9861 3383 9919 3389
rect 9861 3349 9873 3383
rect 9907 3380 9919 3383
rect 10410 3380 10416 3392
rect 9907 3352 10416 3380
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10686 3380 10692 3392
rect 10647 3352 10692 3380
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 17052 3380 17080 3420
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 18892 3448 18920 3479
rect 19150 3476 19156 3488
rect 19208 3476 19214 3528
rect 19058 3448 19064 3460
rect 17184 3420 19064 3448
rect 17184 3408 17190 3420
rect 19058 3408 19064 3420
rect 19116 3408 19122 3460
rect 20070 3380 20076 3392
rect 17052 3352 20076 3380
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 1104 3290 20884 3312
rect 1104 3238 4648 3290
rect 4700 3238 4712 3290
rect 4764 3238 4776 3290
rect 4828 3238 4840 3290
rect 4892 3238 11982 3290
rect 12034 3238 12046 3290
rect 12098 3238 12110 3290
rect 12162 3238 12174 3290
rect 12226 3238 19315 3290
rect 19367 3238 19379 3290
rect 19431 3238 19443 3290
rect 19495 3238 19507 3290
rect 19559 3238 20884 3290
rect 1104 3216 20884 3238
rect 2406 3176 2412 3188
rect 2367 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3176 2470 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2464 3148 2697 3176
rect 2464 3136 2470 3148
rect 2685 3145 2697 3148
rect 2731 3176 2743 3179
rect 2869 3179 2927 3185
rect 2869 3176 2881 3179
rect 2731 3148 2881 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 2869 3145 2881 3148
rect 2915 3145 2927 3179
rect 2869 3139 2927 3145
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 5350 3176 5356 3188
rect 4571 3148 5356 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5500 3148 6193 3176
rect 5500 3136 5506 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10134 3176 10140 3188
rect 10091 3148 10140 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10413 3179 10471 3185
rect 10413 3145 10425 3179
rect 10459 3176 10471 3179
rect 10778 3176 10784 3188
rect 10459 3148 10784 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11514 3176 11520 3188
rect 11011 3148 11520 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 3053 3111 3111 3117
rect 3053 3108 3065 3111
rect 2832 3080 3065 3108
rect 2832 3068 2838 3080
rect 3053 3077 3065 3080
rect 3099 3077 3111 3111
rect 3053 3071 3111 3077
rect 3510 3068 3516 3120
rect 3568 3108 3574 3120
rect 3878 3108 3884 3120
rect 3568 3080 3884 3108
rect 3568 3068 3574 3080
rect 3878 3068 3884 3080
rect 3936 3108 3942 3120
rect 3973 3111 4031 3117
rect 3973 3108 3985 3111
rect 3936 3080 3985 3108
rect 3936 3068 3942 3080
rect 3973 3077 3985 3080
rect 4019 3077 4031 3111
rect 10686 3108 10692 3120
rect 3973 3071 4031 3077
rect 4126 3080 10692 3108
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 4126 3040 4154 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 2179 3012 4154 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4488 3012 4997 3040
rect 4488 3000 4494 3012
rect 4985 3009 4997 3012
rect 5031 3009 5043 3043
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 4985 3003 5043 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 8018 3040 8024 3052
rect 7979 3012 8024 3040
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9306 3040 9312 3052
rect 9171 3012 9312 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 1762 2972 1768 2984
rect 1719 2944 1768 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2314 2972 2320 2984
rect 1995 2944 2320 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 2682 2972 2688 2984
rect 2595 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2972 2746 2984
rect 2961 2975 3019 2981
rect 2961 2972 2973 2975
rect 2740 2944 2973 2972
rect 2740 2932 2746 2944
rect 2961 2941 2973 2944
rect 3007 2941 3019 2975
rect 2961 2935 3019 2941
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3510 2972 3516 2984
rect 3283 2944 3516 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3660 2944 3709 2972
rect 3660 2932 3666 2944
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 6454 2972 6460 2984
rect 4939 2944 6460 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 1912 2876 4016 2904
rect 1912 2864 1918 2876
rect 3988 2836 4016 2876
rect 5092 2836 5120 2944
rect 5321 2913 5349 2944
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 5306 2907 5364 2913
rect 5306 2873 5318 2907
rect 5352 2873 5364 2907
rect 6270 2904 6276 2916
rect 5306 2867 5364 2873
rect 5920 2876 6276 2904
rect 3988 2808 5120 2836
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5920 2845 5948 2876
rect 6270 2864 6276 2876
rect 6328 2904 6334 2916
rect 6549 2907 6607 2913
rect 6549 2904 6561 2907
rect 6328 2876 6561 2904
rect 6328 2864 6334 2876
rect 6549 2873 6561 2876
rect 6595 2904 6607 2907
rect 7009 2907 7067 2913
rect 7009 2904 7021 2907
rect 6595 2876 7021 2904
rect 6595 2873 6607 2876
rect 6549 2867 6607 2873
rect 7009 2873 7021 2876
rect 7055 2873 7067 2907
rect 7009 2867 7067 2873
rect 7466 2864 7472 2916
rect 7524 2904 7530 2916
rect 7524 2876 7569 2904
rect 7524 2864 7530 2876
rect 7834 2864 7840 2916
rect 7892 2904 7898 2916
rect 8389 2907 8447 2913
rect 8389 2904 8401 2907
rect 7892 2876 8401 2904
rect 7892 2864 7898 2876
rect 8389 2873 8401 2876
rect 8435 2904 8447 2907
rect 9033 2907 9091 2913
rect 9033 2904 9045 2907
rect 8435 2876 9045 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 9033 2873 9045 2876
rect 9079 2904 9091 2907
rect 9487 2907 9545 2913
rect 9487 2904 9499 2907
rect 9079 2876 9499 2904
rect 9079 2873 9091 2876
rect 9033 2867 9091 2873
rect 9487 2873 9499 2876
rect 9533 2904 9545 2907
rect 10686 2904 10692 2916
rect 9533 2876 10692 2904
rect 9533 2873 9545 2876
rect 9487 2867 9545 2873
rect 10686 2864 10692 2876
rect 10744 2904 10750 2916
rect 10980 2904 11008 3139
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 11848 3148 12081 3176
rect 11848 3136 11854 3148
rect 12069 3145 12081 3148
rect 12115 3176 12127 3179
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12115 3148 12173 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 13538 3176 13544 3188
rect 13499 3148 13544 3176
rect 12161 3139 12219 3145
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 15105 3179 15163 3185
rect 15105 3145 15117 3179
rect 15151 3176 15163 3179
rect 15470 3176 15476 3188
rect 15151 3148 15476 3176
rect 15151 3145 15163 3148
rect 15105 3139 15163 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 16632 3148 17417 3176
rect 16632 3136 16638 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17405 3139 17463 3145
rect 11425 3111 11483 3117
rect 11425 3077 11437 3111
rect 11471 3108 11483 3111
rect 15930 3108 15936 3120
rect 11471 3080 15936 3108
rect 11471 3077 11483 3080
rect 11425 3071 11483 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 12342 3040 12348 3052
rect 11664 3012 12348 3040
rect 11664 3000 11670 3012
rect 12342 3000 12348 3012
rect 12400 3040 12406 3052
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 12400 3012 12541 3040
rect 12400 3000 12406 3012
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 14090 3040 14096 3052
rect 13219 3012 14096 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 16942 3040 16948 3052
rect 14783 3012 16948 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17420 3040 17448 3139
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 19024 3148 19441 3176
rect 19024 3136 19030 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 19429 3139 19487 3145
rect 19058 3108 19064 3120
rect 19019 3080 19064 3108
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 17420 3012 18092 3040
rect 11238 2972 11244 2984
rect 11199 2944 11244 2972
rect 11238 2932 11244 2944
rect 11296 2972 11302 2984
rect 11422 2972 11428 2984
rect 11296 2944 11428 2972
rect 11296 2932 11302 2944
rect 11422 2932 11428 2944
rect 11480 2972 11486 2984
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11480 2944 11805 2972
rect 11480 2932 11486 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 18064 2981 18092 3012
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 19751 3043 19809 3049
rect 19751 3040 19763 3043
rect 18196 3012 19763 3040
rect 18196 3000 18202 3012
rect 19751 3009 19763 3012
rect 19797 3009 19809 3043
rect 19751 3003 19809 3009
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15344 2944 15577 2972
rect 15344 2932 15350 2944
rect 15565 2941 15577 2944
rect 15611 2972 15623 2975
rect 18049 2975 18107 2981
rect 15611 2944 17540 2972
rect 15611 2941 15623 2944
rect 15565 2935 15623 2941
rect 10744 2876 11008 2904
rect 12069 2907 12127 2913
rect 10744 2864 10750 2876
rect 12069 2873 12081 2907
rect 12115 2904 12127 2907
rect 12621 2907 12679 2913
rect 12621 2904 12633 2907
rect 12115 2876 12633 2904
rect 12115 2873 12127 2876
rect 12069 2867 12127 2873
rect 12621 2873 12633 2876
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 14185 2907 14243 2913
rect 14185 2873 14197 2907
rect 14231 2873 14243 2907
rect 14185 2867 14243 2873
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5500 2808 5917 2836
rect 5500 2796 5506 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 13909 2839 13967 2845
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 14200 2836 14228 2867
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 15381 2907 15439 2913
rect 15381 2904 15393 2907
rect 15160 2876 15393 2904
rect 15160 2864 15166 2876
rect 15381 2873 15393 2876
rect 15427 2904 15439 2907
rect 15886 2907 15944 2913
rect 15886 2904 15898 2907
rect 15427 2876 15898 2904
rect 15427 2873 15439 2876
rect 15381 2867 15439 2873
rect 15886 2873 15898 2876
rect 15932 2904 15944 2907
rect 16850 2904 16856 2916
rect 15932 2876 16856 2904
rect 15932 2873 15944 2876
rect 15886 2867 15944 2873
rect 16850 2864 16856 2876
rect 16908 2904 16914 2916
rect 17037 2907 17095 2913
rect 17037 2904 17049 2907
rect 16908 2876 17049 2904
rect 16908 2864 16914 2876
rect 17037 2873 17049 2876
rect 17083 2873 17095 2907
rect 17037 2867 17095 2873
rect 14550 2836 14556 2848
rect 13955 2808 14556 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 16482 2836 16488 2848
rect 16443 2808 16488 2836
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 17512 2836 17540 2944
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 19664 2975 19722 2981
rect 19664 2941 19676 2975
rect 19710 2972 19722 2975
rect 20070 2972 20076 2984
rect 19710 2944 20076 2972
rect 19710 2941 19722 2944
rect 19664 2935 19722 2941
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 18524 2904 18552 2935
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 17828 2876 18552 2904
rect 17828 2864 17834 2876
rect 18141 2839 18199 2845
rect 18141 2836 18153 2839
rect 17512 2808 18153 2836
rect 18141 2805 18153 2808
rect 18187 2805 18199 2839
rect 18141 2799 18199 2805
rect 1104 2746 20884 2768
rect 1104 2694 8315 2746
rect 8367 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 15648 2746
rect 15700 2694 15712 2746
rect 15764 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 20884 2746
rect 1104 2672 20884 2694
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 2406 2632 2412 2644
rect 2363 2604 2412 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 2406 2592 2412 2604
rect 2464 2632 2470 2644
rect 2866 2632 2872 2644
rect 2464 2604 2872 2632
rect 2464 2592 2470 2604
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3050 2592 3056 2644
rect 3108 2632 3114 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3108 2604 3801 2632
rect 3108 2592 3114 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 3789 2595 3847 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 5258 2632 5264 2644
rect 5123 2604 5264 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6362 2632 6368 2644
rect 6135 2604 6368 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6512 2604 6745 2632
rect 6512 2592 6518 2604
rect 6733 2601 6745 2604
rect 6779 2632 6791 2635
rect 6779 2604 7281 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 5442 2564 5448 2576
rect 1719 2536 5212 2564
rect 5403 2536 5448 2564
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1946 2496 1952 2508
rect 1510 2468 1952 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2406 2496 2412 2508
rect 2367 2468 2412 2496
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 2958 2496 2964 2508
rect 2731 2468 2964 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 3142 2496 3148 2508
rect 3103 2468 3148 2496
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 4090 2499 4148 2505
rect 4090 2465 4102 2499
rect 4136 2496 4148 2499
rect 4136 2468 4660 2496
rect 4136 2465 4148 2468
rect 4090 2459 4148 2465
rect 4632 2440 4660 2468
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5184 2428 5212 2536
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 7006 2564 7012 2576
rect 6043 2536 7012 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 7253 2573 7281 2604
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7524 2604 7849 2632
rect 7524 2592 7530 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 7837 2595 7895 2601
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8803 2635 8861 2641
rect 8803 2632 8815 2635
rect 7984 2604 8815 2632
rect 7984 2592 7990 2604
rect 8803 2601 8815 2604
rect 8849 2601 8861 2635
rect 8803 2595 8861 2601
rect 9214 2592 9220 2644
rect 9272 2632 9278 2644
rect 9907 2635 9965 2641
rect 9907 2632 9919 2635
rect 9272 2604 9919 2632
rect 9272 2592 9278 2604
rect 9907 2601 9919 2604
rect 9953 2601 9965 2635
rect 10686 2632 10692 2644
rect 10647 2604 10692 2632
rect 9907 2595 9965 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11698 2632 11704 2644
rect 11659 2604 11704 2632
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 13078 2632 13084 2644
rect 13039 2604 13084 2632
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 13446 2632 13452 2644
rect 13407 2604 13452 2632
rect 13446 2592 13452 2604
rect 13504 2632 13510 2644
rect 14550 2632 14556 2644
rect 13504 2604 13997 2632
rect 14511 2604 14556 2632
rect 13504 2592 13510 2604
rect 7253 2567 7337 2573
rect 7253 2536 7291 2567
rect 7279 2533 7291 2536
rect 7325 2564 7337 2567
rect 7742 2564 7748 2576
rect 7325 2536 7748 2564
rect 7325 2533 7337 2536
rect 7279 2527 7337 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 8110 2564 8116 2576
rect 8071 2536 8116 2564
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 10704 2564 10732 2592
rect 13969 2573 13997 2604
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 15286 2632 15292 2644
rect 15247 2604 15292 2632
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 16114 2632 16120 2644
rect 16075 2604 16120 2632
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 17310 2632 17316 2644
rect 17271 2604 17316 2632
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17770 2592 17776 2644
rect 17828 2632 17834 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 17828 2604 18061 2632
rect 17828 2592 17834 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 18049 2595 18107 2601
rect 11102 2567 11160 2573
rect 11102 2564 11114 2567
rect 10704 2536 11114 2564
rect 11102 2533 11114 2536
rect 11148 2533 11160 2567
rect 11102 2527 11160 2533
rect 13954 2567 14012 2573
rect 13954 2533 13966 2567
rect 14000 2533 14012 2567
rect 13954 2527 14012 2533
rect 15841 2567 15899 2573
rect 15841 2533 15853 2567
rect 15887 2564 15899 2567
rect 16482 2564 16488 2576
rect 15887 2536 16488 2564
rect 15887 2533 15899 2536
rect 15841 2527 15899 2533
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 17218 2524 17224 2576
rect 17276 2564 17282 2576
rect 17681 2567 17739 2573
rect 17681 2564 17693 2567
rect 17276 2536 17693 2564
rect 17276 2524 17282 2536
rect 17681 2533 17693 2536
rect 17727 2533 17739 2567
rect 18064 2564 18092 2595
rect 18064 2536 18828 2564
rect 17681 2527 17739 2533
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 6914 2456 6920 2468
rect 6972 2496 6978 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 6972 2468 8493 2496
rect 6972 2456 6978 2468
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8732 2499 8790 2505
rect 8732 2465 8744 2499
rect 8778 2496 8790 2499
rect 9122 2496 9128 2508
rect 8778 2468 9128 2496
rect 8778 2465 8790 2468
rect 8732 2459 8790 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9858 2505 9864 2508
rect 9836 2499 9864 2505
rect 9836 2496 9848 2499
rect 9771 2468 9848 2496
rect 9836 2465 9848 2468
rect 9916 2496 9922 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9916 2468 10241 2496
rect 9836 2459 9864 2465
rect 9858 2456 9864 2459
rect 9916 2456 9922 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 12688 2499 12746 2505
rect 12688 2465 12700 2499
rect 12734 2496 12746 2499
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 12734 2468 16037 2496
rect 12734 2465 12746 2468
rect 12688 2459 12746 2465
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 17696 2496 17724 2527
rect 18800 2505 18828 2536
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17696 2468 18337 2496
rect 16025 2459 16083 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 18785 2499 18843 2505
rect 18785 2465 18797 2499
rect 18831 2465 18843 2499
rect 18785 2459 18843 2465
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5184 2400 5365 2428
rect 5353 2397 5365 2400
rect 5399 2428 5411 2431
rect 10781 2431 10839 2437
rect 5399 2400 6316 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 2501 2363 2559 2369
rect 2501 2329 2513 2363
rect 2547 2360 2559 2363
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 2547 2332 6101 2360
rect 2547 2329 2559 2332
rect 2501 2323 2559 2329
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6288 2360 6316 2400
rect 10781 2397 10793 2431
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 6288 2332 9505 2360
rect 6089 2323 6147 2329
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 10796 2360 10824 2391
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13136 2400 13645 2428
rect 13136 2388 13142 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16393 2431 16451 2437
rect 16393 2428 16405 2431
rect 16172 2400 16405 2428
rect 16172 2388 16178 2400
rect 16393 2397 16405 2400
rect 16439 2397 16451 2431
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 16393 2391 16451 2397
rect 16500 2400 18889 2428
rect 12069 2363 12127 2369
rect 12069 2360 12081 2363
rect 10796 2332 12081 2360
rect 9493 2323 9551 2329
rect 12069 2329 12081 2332
rect 12115 2360 12127 2363
rect 16500 2360 16528 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 16942 2360 16948 2372
rect 12115 2332 16528 2360
rect 16903 2332 16948 2360
rect 12115 2329 12127 2332
rect 12069 2323 12127 2329
rect 16942 2320 16948 2332
rect 17000 2320 17006 2372
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 3510 2292 3516 2304
rect 3471 2264 3516 2292
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 12759 2295 12817 2301
rect 12759 2261 12771 2295
rect 12805 2292 12817 2295
rect 12986 2292 12992 2304
rect 12805 2264 12992 2292
rect 12805 2261 12817 2264
rect 12759 2255 12817 2261
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 16025 2295 16083 2301
rect 16025 2261 16037 2295
rect 16071 2292 16083 2295
rect 19150 2292 19156 2304
rect 16071 2264 19156 2292
rect 16071 2261 16083 2264
rect 16025 2255 16083 2261
rect 19150 2252 19156 2264
rect 19208 2292 19214 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 19208 2264 19349 2292
rect 19208 2252 19214 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 1104 2202 20884 2224
rect 1104 2150 4648 2202
rect 4700 2150 4712 2202
rect 4764 2150 4776 2202
rect 4828 2150 4840 2202
rect 4892 2150 11982 2202
rect 12034 2150 12046 2202
rect 12098 2150 12110 2202
rect 12162 2150 12174 2202
rect 12226 2150 19315 2202
rect 19367 2150 19379 2202
rect 19431 2150 19443 2202
rect 19495 2150 19507 2202
rect 19559 2150 20884 2202
rect 1104 2128 20884 2150
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 18138 2020 18144 2032
rect 10100 1992 18144 2020
rect 10100 1980 10106 1992
rect 18138 1980 18144 1992
rect 18196 1980 18202 2032
rect 11146 144 11152 196
rect 11204 184 11210 196
rect 11204 156 11278 184
rect 11204 144 11210 156
rect 11250 48 11278 156
rect 12986 76 12992 128
rect 13044 116 13050 128
rect 19150 116 19156 128
rect 13044 88 19156 116
rect 13044 76 13050 88
rect 19150 76 19156 88
rect 19208 76 19214 128
rect 16942 48 16948 60
rect 11250 20 16948 48
rect 16942 8 16948 20
rect 17000 8 17006 60
<< via1 >>
rect 16580 21496 16632 21548
rect 17316 21496 17368 21548
rect 4648 19558 4700 19610
rect 4712 19558 4764 19610
rect 4776 19558 4828 19610
rect 4840 19558 4892 19610
rect 11982 19558 12034 19610
rect 12046 19558 12098 19610
rect 12110 19558 12162 19610
rect 12174 19558 12226 19610
rect 19315 19558 19367 19610
rect 19379 19558 19431 19610
rect 19443 19558 19495 19610
rect 19507 19558 19559 19610
rect 11060 19388 11112 19440
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 10968 19116 11020 19168
rect 11612 19159 11664 19168
rect 11612 19125 11621 19159
rect 11621 19125 11655 19159
rect 11655 19125 11664 19159
rect 11612 19116 11664 19125
rect 12624 19116 12676 19168
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 13820 19116 13872 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 8315 19014 8367 19066
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 15648 19014 15700 19066
rect 15712 19014 15764 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 10692 18912 10744 18964
rect 19156 18912 19208 18964
rect 6552 18844 6604 18896
rect 10508 18844 10560 18896
rect 8208 18776 8260 18828
rect 10692 18819 10744 18828
rect 10692 18785 10710 18819
rect 10710 18785 10744 18819
rect 10692 18776 10744 18785
rect 11520 18776 11572 18828
rect 11796 18776 11848 18828
rect 13360 18776 13412 18828
rect 16028 18776 16080 18828
rect 8852 18572 8904 18624
rect 10876 18572 10928 18624
rect 11520 18572 11572 18624
rect 13728 18572 13780 18624
rect 14832 18572 14884 18624
rect 4648 18470 4700 18522
rect 4712 18470 4764 18522
rect 4776 18470 4828 18522
rect 4840 18470 4892 18522
rect 11982 18470 12034 18522
rect 12046 18470 12098 18522
rect 12110 18470 12162 18522
rect 12174 18470 12226 18522
rect 19315 18470 19367 18522
rect 19379 18470 19431 18522
rect 19443 18470 19495 18522
rect 19507 18470 19559 18522
rect 7748 18368 7800 18420
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 11796 18368 11848 18420
rect 7380 18300 7432 18352
rect 4436 18232 4488 18284
rect 15200 18368 15252 18420
rect 14372 18300 14424 18352
rect 14556 18300 14608 18352
rect 8760 18096 8812 18148
rect 11152 18164 11204 18216
rect 11612 18207 11664 18216
rect 11612 18173 11621 18207
rect 11621 18173 11655 18207
rect 11655 18173 11664 18207
rect 11612 18164 11664 18173
rect 13268 18164 13320 18216
rect 13544 18164 13596 18216
rect 10692 18096 10744 18148
rect 11888 18096 11940 18148
rect 14740 18096 14792 18148
rect 18512 18139 18564 18148
rect 18512 18105 18521 18139
rect 18521 18105 18555 18139
rect 18555 18105 18564 18139
rect 18512 18096 18564 18105
rect 8208 18028 8260 18080
rect 9404 18071 9456 18080
rect 9404 18037 9413 18071
rect 9413 18037 9447 18071
rect 9447 18037 9456 18071
rect 9404 18028 9456 18037
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 12808 18028 12860 18080
rect 13360 18028 13412 18080
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 16396 18028 16448 18080
rect 8315 17926 8367 17978
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 15648 17926 15700 17978
rect 15712 17926 15764 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 13084 17824 13136 17876
rect 9404 17756 9456 17808
rect 16764 17756 16816 17808
rect 6368 17688 6420 17740
rect 7748 17688 7800 17740
rect 8668 17688 8720 17740
rect 11704 17688 11756 17740
rect 13544 17731 13596 17740
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 17408 17688 17460 17740
rect 18696 17688 18748 17740
rect 19156 17688 19208 17740
rect 19708 17688 19760 17740
rect 13452 17620 13504 17672
rect 15384 17620 15436 17672
rect 17224 17552 17276 17604
rect 6552 17484 6604 17536
rect 7564 17484 7616 17536
rect 9128 17484 9180 17536
rect 11796 17484 11848 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 12716 17484 12768 17536
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 16028 17484 16080 17536
rect 17592 17484 17644 17536
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 18604 17484 18656 17536
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 4648 17382 4700 17434
rect 4712 17382 4764 17434
rect 4776 17382 4828 17434
rect 4840 17382 4892 17434
rect 11982 17382 12034 17434
rect 12046 17382 12098 17434
rect 12110 17382 12162 17434
rect 12174 17382 12226 17434
rect 19315 17382 19367 17434
rect 19379 17382 19431 17434
rect 19443 17382 19495 17434
rect 19507 17382 19559 17434
rect 6368 17323 6420 17332
rect 6368 17289 6377 17323
rect 6377 17289 6411 17323
rect 6411 17289 6420 17323
rect 6368 17280 6420 17289
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 9588 17280 9640 17332
rect 10508 17280 10560 17332
rect 19616 17280 19668 17332
rect 19708 17323 19760 17332
rect 19708 17289 19717 17323
rect 19717 17289 19751 17323
rect 19751 17289 19760 17323
rect 19708 17280 19760 17289
rect 112 17212 164 17264
rect 11336 17212 11388 17264
rect 11704 17212 11756 17264
rect 13360 17212 13412 17264
rect 16304 17255 16356 17264
rect 16304 17221 16313 17255
rect 16313 17221 16347 17255
rect 16347 17221 16356 17255
rect 16304 17212 16356 17221
rect 9404 17144 9456 17196
rect 10600 17144 10652 17196
rect 8024 17076 8076 17128
rect 9956 17076 10008 17128
rect 10508 17076 10560 17128
rect 12716 17144 12768 17196
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 7748 17051 7800 17060
rect 7748 17017 7757 17051
rect 7757 17017 7791 17051
rect 7791 17017 7800 17051
rect 7748 17008 7800 17017
rect 10784 17008 10836 17060
rect 12532 17076 12584 17128
rect 13820 17076 13872 17128
rect 14096 17144 14148 17196
rect 14372 17144 14424 17196
rect 12808 17008 12860 17060
rect 7288 16940 7340 16992
rect 9220 16940 9272 16992
rect 10048 16940 10100 16992
rect 11704 16940 11756 16992
rect 12716 16940 12768 16992
rect 13544 16940 13596 16992
rect 17776 17076 17828 17128
rect 18052 17119 18104 17128
rect 18052 17085 18096 17119
rect 18096 17085 18104 17119
rect 19064 17119 19116 17128
rect 18052 17076 18104 17085
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 18420 17008 18472 17060
rect 14372 16940 14424 16992
rect 15292 16940 15344 16992
rect 17408 16940 17460 16992
rect 18512 16940 18564 16992
rect 18696 16983 18748 16992
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 8315 16838 8367 16890
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 15648 16838 15700 16890
rect 15712 16838 15764 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 9772 16736 9824 16788
rect 12348 16779 12400 16788
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 13912 16779 13964 16788
rect 13912 16745 13921 16779
rect 13921 16745 13955 16779
rect 13955 16745 13964 16779
rect 13912 16736 13964 16745
rect 19524 16736 19576 16788
rect 2044 16668 2096 16720
rect 5540 16600 5592 16652
rect 6644 16600 6696 16652
rect 8760 16600 8812 16652
rect 10140 16600 10192 16652
rect 10232 16532 10284 16584
rect 12716 16600 12768 16652
rect 13728 16643 13780 16652
rect 13728 16609 13737 16643
rect 13737 16609 13771 16643
rect 13771 16609 13780 16643
rect 13728 16600 13780 16609
rect 14004 16600 14056 16652
rect 16120 16600 16172 16652
rect 18696 16600 18748 16652
rect 19616 16600 19668 16652
rect 12900 16532 12952 16584
rect 14924 16532 14976 16584
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 17132 16532 17184 16584
rect 5448 16396 5500 16448
rect 6736 16396 6788 16448
rect 6920 16396 6972 16448
rect 7932 16396 7984 16448
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 4648 16294 4700 16346
rect 4712 16294 4764 16346
rect 4776 16294 4828 16346
rect 4840 16294 4892 16346
rect 11982 16294 12034 16346
rect 12046 16294 12098 16346
rect 12110 16294 12162 16346
rect 12174 16294 12226 16346
rect 19315 16294 19367 16346
rect 19379 16294 19431 16346
rect 19443 16294 19495 16346
rect 19507 16294 19559 16346
rect 6644 16192 6696 16244
rect 9312 16192 9364 16244
rect 10600 16192 10652 16244
rect 13728 16192 13780 16244
rect 16764 16192 16816 16244
rect 19616 16235 19668 16244
rect 19616 16201 19625 16235
rect 19625 16201 19659 16235
rect 19659 16201 19668 16235
rect 19616 16192 19668 16201
rect 112 16124 164 16176
rect 1308 16056 1360 16108
rect 5908 16124 5960 16176
rect 7932 16124 7984 16176
rect 9036 16167 9088 16176
rect 9036 16133 9045 16167
rect 9045 16133 9079 16167
rect 9079 16133 9088 16167
rect 9036 16124 9088 16133
rect 6184 16056 6236 16108
rect 8760 16056 8812 16108
rect 9312 16056 9364 16108
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 2872 15852 2924 15904
rect 3976 15852 4028 15904
rect 4528 15988 4580 16040
rect 5724 15988 5776 16040
rect 6644 15988 6696 16040
rect 10140 15988 10192 16040
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 6828 15920 6880 15972
rect 8668 15920 8720 15972
rect 9496 15963 9548 15972
rect 9496 15929 9505 15963
rect 9505 15929 9539 15963
rect 9539 15929 9548 15963
rect 9496 15920 9548 15929
rect 12808 15988 12860 16040
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 11428 15920 11480 15972
rect 11612 15920 11664 15972
rect 4344 15852 4396 15904
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 8116 15852 8168 15904
rect 8852 15852 8904 15904
rect 10324 15852 10376 15904
rect 12716 15920 12768 15972
rect 16304 15988 16356 16040
rect 14280 15920 14332 15972
rect 16120 15920 16172 15972
rect 12808 15852 12860 15904
rect 14004 15852 14056 15904
rect 17316 15988 17368 16040
rect 16672 15963 16724 15972
rect 16672 15929 16681 15963
rect 16681 15929 16715 15963
rect 16715 15929 16724 15963
rect 16672 15920 16724 15929
rect 19708 15920 19760 15972
rect 16948 15852 17000 15904
rect 18880 15852 18932 15904
rect 8315 15750 8367 15802
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 15648 15750 15700 15802
rect 15712 15750 15764 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 18972 15648 19024 15700
rect 21548 15648 21600 15700
rect 3884 15580 3936 15632
rect 7932 15580 7984 15632
rect 5356 15555 5408 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 4988 15444 5040 15496
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 6460 15512 6512 15564
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 11336 15580 11388 15632
rect 9772 15555 9824 15564
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 15476 15512 15528 15564
rect 16120 15512 16172 15564
rect 16948 15512 17000 15564
rect 17776 15512 17828 15564
rect 19156 15512 19208 15564
rect 9036 15444 9088 15496
rect 3240 15376 3292 15428
rect 7104 15376 7156 15428
rect 11244 15444 11296 15496
rect 14188 15487 14240 15496
rect 14188 15453 14197 15487
rect 14197 15453 14231 15487
rect 14231 15453 14240 15487
rect 14188 15444 14240 15453
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 12900 15376 12952 15428
rect 13544 15376 13596 15428
rect 17408 15376 17460 15428
rect 4252 15308 4304 15360
rect 9312 15308 9364 15360
rect 14464 15351 14516 15360
rect 14464 15317 14473 15351
rect 14473 15317 14507 15351
rect 14507 15317 14516 15351
rect 14464 15308 14516 15317
rect 16304 15308 16356 15360
rect 17960 15308 18012 15360
rect 4648 15206 4700 15258
rect 4712 15206 4764 15258
rect 4776 15206 4828 15258
rect 4840 15206 4892 15258
rect 11982 15206 12034 15258
rect 12046 15206 12098 15258
rect 12110 15206 12162 15258
rect 12174 15206 12226 15258
rect 19315 15206 19367 15258
rect 19379 15206 19431 15258
rect 19443 15206 19495 15258
rect 19507 15206 19559 15258
rect 1860 14900 1912 14952
rect 2320 15104 2372 15156
rect 3240 15104 3292 15156
rect 7840 15104 7892 15156
rect 8208 15104 8260 15156
rect 9404 15104 9456 15156
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 14096 15104 14148 15156
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 19156 15147 19208 15156
rect 19156 15113 19165 15147
rect 19165 15113 19199 15147
rect 19199 15113 19208 15147
rect 19156 15104 19208 15113
rect 4528 15036 4580 15088
rect 4436 14968 4488 15020
rect 6460 15011 6512 15020
rect 6460 14977 6469 15011
rect 6469 14977 6503 15011
rect 6503 14977 6512 15011
rect 6460 14968 6512 14977
rect 10784 15036 10836 15088
rect 13728 15036 13780 15088
rect 14004 15036 14056 15088
rect 18328 15036 18380 15088
rect 8944 15011 8996 15020
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 3608 14900 3660 14952
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 3056 14875 3108 14884
rect 3056 14841 3065 14875
rect 3065 14841 3099 14875
rect 3099 14841 3108 14875
rect 3056 14832 3108 14841
rect 112 14764 164 14816
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 5356 14832 5408 14884
rect 7196 14900 7248 14952
rect 7932 14900 7984 14952
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 9312 14968 9364 15020
rect 9496 14968 9548 15020
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 14648 14968 14700 15020
rect 10508 14943 10560 14952
rect 10508 14909 10517 14943
rect 10517 14909 10551 14943
rect 10551 14909 10560 14943
rect 10508 14900 10560 14909
rect 10784 14900 10836 14952
rect 11336 14900 11388 14952
rect 13820 14900 13872 14952
rect 17776 14968 17828 15020
rect 12900 14875 12952 14884
rect 12900 14841 12909 14875
rect 12909 14841 12943 14875
rect 12943 14841 12952 14875
rect 12900 14832 12952 14841
rect 4528 14764 4580 14773
rect 5172 14764 5224 14816
rect 7012 14764 7064 14816
rect 9036 14764 9088 14816
rect 10416 14764 10468 14816
rect 11428 14764 11480 14816
rect 14648 14832 14700 14884
rect 17408 14900 17460 14952
rect 18236 14900 18288 14952
rect 18328 14900 18380 14952
rect 15936 14875 15988 14884
rect 15936 14841 15945 14875
rect 15945 14841 15979 14875
rect 15979 14841 15988 14875
rect 15936 14832 15988 14841
rect 18788 14832 18840 14884
rect 13544 14764 13596 14816
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 16948 14764 17000 14816
rect 17408 14764 17460 14816
rect 18144 14807 18196 14816
rect 18144 14773 18153 14807
rect 18153 14773 18187 14807
rect 18187 14773 18196 14807
rect 18144 14764 18196 14773
rect 8315 14662 8367 14714
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 15648 14662 15700 14714
rect 15712 14662 15764 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 5724 14560 5776 14612
rect 6644 14560 6696 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 12900 14603 12952 14612
rect 12900 14569 12909 14603
rect 12909 14569 12943 14603
rect 12943 14569 12952 14603
rect 12900 14560 12952 14569
rect 14648 14560 14700 14612
rect 4528 14492 4580 14544
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 2688 14424 2740 14476
rect 4988 14424 5040 14476
rect 7472 14492 7524 14544
rect 9312 14492 9364 14544
rect 9496 14492 9548 14544
rect 10508 14492 10560 14544
rect 8300 14467 8352 14476
rect 5264 14356 5316 14408
rect 6460 14356 6512 14408
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 7196 14356 7248 14408
rect 9312 14356 9364 14408
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 9956 14356 10008 14408
rect 10508 14356 10560 14408
rect 5356 14288 5408 14340
rect 2596 14263 2648 14272
rect 2596 14229 2605 14263
rect 2605 14229 2639 14263
rect 2639 14229 2648 14263
rect 2596 14220 2648 14229
rect 2780 14220 2832 14272
rect 8668 14288 8720 14340
rect 8852 14288 8904 14340
rect 11796 14492 11848 14544
rect 12348 14492 12400 14544
rect 13176 14535 13228 14544
rect 13176 14501 13185 14535
rect 13185 14501 13219 14535
rect 13219 14501 13228 14535
rect 13176 14492 13228 14501
rect 13820 14492 13872 14544
rect 15108 14492 15160 14544
rect 15936 14560 15988 14612
rect 16948 14603 17000 14612
rect 16948 14569 16957 14603
rect 16957 14569 16991 14603
rect 16991 14569 17000 14603
rect 16948 14560 17000 14569
rect 17868 14560 17920 14612
rect 18328 14492 18380 14544
rect 10784 14424 10836 14476
rect 11428 14424 11480 14476
rect 16488 14424 16540 14476
rect 16764 14424 16816 14476
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 18236 14424 18288 14476
rect 18972 14467 19024 14476
rect 18972 14433 18981 14467
rect 18981 14433 19015 14467
rect 19015 14433 19024 14467
rect 18972 14424 19024 14433
rect 11796 14356 11848 14408
rect 12624 14356 12676 14408
rect 12808 14356 12860 14408
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 15476 14356 15528 14408
rect 13728 14288 13780 14340
rect 14096 14288 14148 14340
rect 16120 14288 16172 14340
rect 10784 14220 10836 14272
rect 12716 14220 12768 14272
rect 13452 14220 13504 14272
rect 18328 14220 18380 14272
rect 4648 14118 4700 14170
rect 4712 14118 4764 14170
rect 4776 14118 4828 14170
rect 4840 14118 4892 14170
rect 11982 14118 12034 14170
rect 12046 14118 12098 14170
rect 12110 14118 12162 14170
rect 12174 14118 12226 14170
rect 19315 14118 19367 14170
rect 19379 14118 19431 14170
rect 19443 14118 19495 14170
rect 19507 14118 19559 14170
rect 2596 13948 2648 14000
rect 7656 14016 7708 14068
rect 8300 14016 8352 14068
rect 3516 13948 3568 14000
rect 5724 13948 5776 14000
rect 8668 13948 8720 14000
rect 8760 13948 8812 14000
rect 9588 13948 9640 14000
rect 9772 14016 9824 14068
rect 12900 14016 12952 14068
rect 13360 14016 13412 14068
rect 14648 14016 14700 14068
rect 15108 14059 15160 14068
rect 15108 14025 15117 14059
rect 15117 14025 15151 14059
rect 15151 14025 15160 14059
rect 15108 14016 15160 14025
rect 16488 14016 16540 14068
rect 9864 13991 9916 14000
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 3240 13880 3292 13932
rect 1676 13812 1728 13864
rect 2136 13812 2188 13864
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 2964 13812 3016 13864
rect 3516 13855 3568 13864
rect 2228 13787 2280 13796
rect 2228 13753 2237 13787
rect 2237 13753 2271 13787
rect 2271 13753 2280 13787
rect 2228 13744 2280 13753
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 2504 13676 2556 13728
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 4988 13812 5040 13864
rect 5356 13880 5408 13932
rect 7472 13880 7524 13932
rect 8852 13880 8904 13932
rect 9772 13880 9824 13932
rect 10324 13948 10376 14000
rect 10508 13948 10560 14000
rect 12808 13948 12860 14000
rect 15384 13948 15436 14000
rect 16764 13948 16816 14000
rect 20628 13948 20680 14000
rect 10784 13880 10836 13932
rect 11428 13923 11480 13932
rect 11428 13889 11437 13923
rect 11437 13889 11471 13923
rect 11471 13889 11480 13923
rect 11428 13880 11480 13889
rect 13268 13880 13320 13932
rect 3424 13744 3476 13796
rect 4528 13676 4580 13728
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 6092 13676 6144 13728
rect 7656 13812 7708 13864
rect 8760 13812 8812 13864
rect 12900 13812 12952 13864
rect 13452 13855 13504 13864
rect 13452 13821 13461 13855
rect 13461 13821 13495 13855
rect 13495 13821 13504 13855
rect 13452 13812 13504 13821
rect 13544 13812 13596 13864
rect 16120 13880 16172 13932
rect 16488 13880 16540 13932
rect 17408 13812 17460 13864
rect 18328 13880 18380 13932
rect 7748 13787 7800 13796
rect 7748 13753 7757 13787
rect 7757 13753 7791 13787
rect 7791 13753 7800 13787
rect 7748 13744 7800 13753
rect 8852 13676 8904 13728
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 10876 13676 10928 13728
rect 12072 13676 12124 13728
rect 12716 13676 12768 13728
rect 14648 13744 14700 13796
rect 15476 13744 15528 13796
rect 17500 13744 17552 13796
rect 18972 13812 19024 13864
rect 19156 13812 19208 13864
rect 16120 13676 16172 13728
rect 18144 13719 18196 13728
rect 18144 13685 18153 13719
rect 18153 13685 18187 13719
rect 18187 13685 18196 13719
rect 18144 13676 18196 13685
rect 19616 13676 19668 13728
rect 8315 13574 8367 13626
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 15648 13574 15700 13626
rect 15712 13574 15764 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 1768 13472 1820 13524
rect 3516 13472 3568 13524
rect 3792 13472 3844 13524
rect 2964 13379 3016 13388
rect 2964 13345 2973 13379
rect 2973 13345 3007 13379
rect 3007 13345 3016 13379
rect 2964 13336 3016 13345
rect 3424 13336 3476 13388
rect 3332 13268 3384 13320
rect 3976 13404 4028 13456
rect 4988 13472 5040 13524
rect 5632 13472 5684 13524
rect 9496 13515 9548 13524
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 5540 13404 5592 13456
rect 8760 13447 8812 13456
rect 8760 13413 8769 13447
rect 8769 13413 8803 13447
rect 8803 13413 8812 13447
rect 8760 13404 8812 13413
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 6092 13379 6144 13388
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 6460 13336 6512 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 8668 13336 8720 13388
rect 11428 13472 11480 13524
rect 13544 13472 13596 13524
rect 16580 13472 16632 13524
rect 18236 13472 18288 13524
rect 9956 13447 10008 13456
rect 9956 13413 9965 13447
rect 9965 13413 9999 13447
rect 9999 13413 10008 13447
rect 9956 13404 10008 13413
rect 12716 13404 12768 13456
rect 13176 13447 13228 13456
rect 13176 13413 13185 13447
rect 13185 13413 13219 13447
rect 13219 13413 13228 13447
rect 13176 13404 13228 13413
rect 14648 13404 14700 13456
rect 15200 13404 15252 13456
rect 17684 13404 17736 13456
rect 14004 13336 14056 13388
rect 18696 13336 18748 13388
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 4344 13268 4396 13320
rect 8024 13268 8076 13320
rect 9312 13268 9364 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 10600 13268 10652 13320
rect 11428 13268 11480 13320
rect 15108 13268 15160 13320
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16764 13311 16816 13320
rect 16028 13268 16080 13277
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 16948 13268 17000 13320
rect 17500 13268 17552 13320
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 19064 13268 19116 13320
rect 1676 13132 1728 13184
rect 6460 13200 6512 13252
rect 7656 13200 7708 13252
rect 9496 13200 9548 13252
rect 12072 13200 12124 13252
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 5356 13132 5408 13184
rect 6000 13132 6052 13184
rect 6092 13132 6144 13184
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 16304 13132 16356 13184
rect 16948 13132 17000 13184
rect 18236 13175 18288 13184
rect 18236 13141 18245 13175
rect 18245 13141 18279 13175
rect 18279 13141 18288 13175
rect 18236 13132 18288 13141
rect 4648 13030 4700 13082
rect 4712 13030 4764 13082
rect 4776 13030 4828 13082
rect 4840 13030 4892 13082
rect 11982 13030 12034 13082
rect 12046 13030 12098 13082
rect 12110 13030 12162 13082
rect 12174 13030 12226 13082
rect 19315 13030 19367 13082
rect 19379 13030 19431 13082
rect 19443 13030 19495 13082
rect 19507 13030 19559 13082
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 4160 12928 4212 12980
rect 5172 12928 5224 12980
rect 5816 12928 5868 12980
rect 8300 12928 8352 12980
rect 8760 12928 8812 12980
rect 9404 12928 9456 12980
rect 10876 12928 10928 12980
rect 13912 12971 13964 12980
rect 13912 12937 13921 12971
rect 13921 12937 13955 12971
rect 13955 12937 13964 12971
rect 13912 12928 13964 12937
rect 15200 12928 15252 12980
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 18880 12928 18932 12980
rect 6644 12860 6696 12912
rect 7104 12860 7156 12912
rect 9680 12860 9732 12912
rect 11428 12860 11480 12912
rect 11612 12860 11664 12912
rect 13360 12860 13412 12912
rect 2964 12792 3016 12844
rect 3424 12792 3476 12844
rect 4344 12792 4396 12844
rect 5356 12792 5408 12844
rect 5724 12792 5776 12844
rect 6736 12792 6788 12844
rect 8300 12792 8352 12844
rect 9496 12792 9548 12844
rect 12348 12792 12400 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13176 12792 13228 12844
rect 16120 12860 16172 12912
rect 16580 12860 16632 12912
rect 18604 12860 18656 12912
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 3148 12656 3200 12708
rect 4896 12699 4948 12708
rect 4896 12665 4905 12699
rect 4905 12665 4939 12699
rect 4939 12665 4948 12699
rect 4896 12656 4948 12665
rect 1308 12588 1360 12640
rect 4160 12588 4212 12640
rect 6092 12588 6144 12640
rect 6276 12631 6328 12640
rect 6276 12597 6285 12631
rect 6285 12597 6319 12631
rect 6319 12597 6328 12631
rect 6276 12588 6328 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 7840 12656 7892 12708
rect 6644 12588 6696 12597
rect 8668 12588 8720 12640
rect 8852 12588 8904 12640
rect 9956 12588 10008 12640
rect 11612 12588 11664 12640
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 12624 12699 12676 12708
rect 12624 12665 12633 12699
rect 12633 12665 12667 12699
rect 12667 12665 12676 12699
rect 12624 12656 12676 12665
rect 12716 12588 12768 12640
rect 16212 12792 16264 12844
rect 16856 12792 16908 12844
rect 17316 12792 17368 12844
rect 17500 12792 17552 12844
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 13820 12724 13872 12776
rect 16580 12767 16632 12776
rect 16580 12733 16589 12767
rect 16589 12733 16623 12767
rect 16623 12733 16632 12767
rect 16580 12724 16632 12733
rect 14004 12656 14056 12708
rect 14096 12588 14148 12640
rect 16856 12699 16908 12708
rect 15384 12588 15436 12640
rect 16856 12665 16865 12699
rect 16865 12665 16899 12699
rect 16899 12665 16908 12699
rect 16856 12656 16908 12665
rect 17316 12588 17368 12640
rect 18052 12588 18104 12640
rect 8315 12486 8367 12538
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 15648 12486 15700 12538
rect 15712 12486 15764 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 1768 12384 1820 12436
rect 2044 12316 2096 12368
rect 1584 12248 1636 12300
rect 3332 12384 3384 12436
rect 3424 12316 3476 12368
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 3976 12316 4028 12368
rect 5448 12384 5500 12436
rect 6092 12384 6144 12436
rect 6644 12384 6696 12436
rect 10416 12384 10468 12436
rect 11244 12384 11296 12436
rect 12348 12384 12400 12436
rect 14280 12427 14332 12436
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 17040 12384 17092 12436
rect 9220 12359 9272 12368
rect 9220 12325 9229 12359
rect 9229 12325 9263 12359
rect 9263 12325 9272 12359
rect 9220 12316 9272 12325
rect 9312 12316 9364 12368
rect 10600 12316 10652 12368
rect 6736 12248 6788 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 12164 12248 12216 12300
rect 12348 12248 12400 12300
rect 13728 12316 13780 12368
rect 15016 12316 15068 12368
rect 13268 12248 13320 12300
rect 17316 12384 17368 12436
rect 19156 12384 19208 12436
rect 17684 12316 17736 12368
rect 18696 12316 18748 12368
rect 2780 12180 2832 12232
rect 4528 12112 4580 12164
rect 4896 12112 4948 12164
rect 11244 12180 11296 12232
rect 14648 12180 14700 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 18972 12180 19024 12232
rect 10508 12112 10560 12164
rect 19064 12112 19116 12164
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 5172 12044 5224 12096
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 4648 11942 4700 11994
rect 4712 11942 4764 11994
rect 4776 11942 4828 11994
rect 4840 11942 4892 11994
rect 11982 11942 12034 11994
rect 12046 11942 12098 11994
rect 12110 11942 12162 11994
rect 12174 11942 12226 11994
rect 19315 11942 19367 11994
rect 19379 11942 19431 11994
rect 19443 11942 19495 11994
rect 19507 11942 19559 11994
rect 3148 11883 3200 11892
rect 3148 11849 3157 11883
rect 3157 11849 3191 11883
rect 3191 11849 3200 11883
rect 3148 11840 3200 11849
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 4988 11840 5040 11892
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 8024 11840 8076 11892
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 13268 11840 13320 11892
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 19156 11840 19208 11892
rect 3976 11772 4028 11824
rect 3424 11704 3476 11756
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 3148 11568 3200 11620
rect 6092 11772 6144 11824
rect 16304 11772 16356 11824
rect 18604 11772 18656 11824
rect 4344 11704 4396 11756
rect 5080 11704 5132 11756
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 10048 11704 10100 11756
rect 10600 11704 10652 11756
rect 8576 11636 8628 11688
rect 9312 11636 9364 11688
rect 11612 11704 11664 11756
rect 14280 11704 14332 11756
rect 11152 11636 11204 11688
rect 16948 11704 17000 11756
rect 18144 11704 18196 11756
rect 5080 11611 5132 11620
rect 5080 11577 5089 11611
rect 5089 11577 5123 11611
rect 5123 11577 5132 11611
rect 5080 11568 5132 11577
rect 7564 11611 7616 11620
rect 2320 11500 2372 11552
rect 2964 11500 3016 11552
rect 4988 11500 5040 11552
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 6644 11500 6696 11552
rect 7564 11577 7573 11611
rect 7573 11577 7607 11611
rect 7607 11577 7616 11611
rect 7564 11568 7616 11577
rect 9864 11568 9916 11620
rect 10508 11611 10560 11620
rect 10508 11577 10517 11611
rect 10517 11577 10551 11611
rect 10551 11577 10560 11611
rect 10508 11568 10560 11577
rect 8116 11500 8168 11552
rect 11612 11500 11664 11552
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 12624 11611 12676 11620
rect 12624 11577 12633 11611
rect 12633 11577 12667 11611
rect 12667 11577 12676 11611
rect 12624 11568 12676 11577
rect 13268 11568 13320 11620
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 16304 11568 16356 11620
rect 17040 11636 17092 11688
rect 18972 11636 19024 11688
rect 16764 11568 16816 11620
rect 17316 11568 17368 11620
rect 15108 11543 15160 11552
rect 14096 11500 14148 11509
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 19064 11500 19116 11552
rect 8315 11398 8367 11450
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 15648 11398 15700 11450
rect 15712 11398 15764 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 2044 11296 2096 11348
rect 2412 11339 2464 11348
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 3516 11296 3568 11348
rect 6460 11296 6512 11348
rect 6828 11296 6880 11348
rect 10048 11296 10100 11348
rect 11152 11296 11204 11348
rect 1952 11228 2004 11280
rect 3976 11228 4028 11280
rect 6092 11228 6144 11280
rect 6644 11228 6696 11280
rect 10508 11228 10560 11280
rect 10784 11228 10836 11280
rect 11244 11228 11296 11280
rect 12164 11296 12216 11348
rect 12624 11296 12676 11348
rect 13728 11296 13780 11348
rect 14188 11296 14240 11348
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 18144 11296 18196 11348
rect 18512 11296 18564 11348
rect 12348 11228 12400 11280
rect 15108 11228 15160 11280
rect 16028 11271 16080 11280
rect 16028 11237 16037 11271
rect 16037 11237 16071 11271
rect 16071 11237 16080 11271
rect 16028 11228 16080 11237
rect 17316 11228 17368 11280
rect 19064 11271 19116 11280
rect 19064 11237 19073 11271
rect 19073 11237 19107 11271
rect 19107 11237 19116 11271
rect 19064 11228 19116 11237
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 6920 11160 6972 11212
rect 9220 11160 9272 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 11336 11160 11388 11212
rect 17868 11160 17920 11212
rect 2872 11092 2924 11144
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 5724 11135 5776 11144
rect 2228 11024 2280 11076
rect 3608 11024 3660 11076
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 7380 11092 7432 11144
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 8024 11092 8076 11144
rect 10784 11092 10836 11144
rect 11704 11092 11756 11144
rect 12716 11092 12768 11144
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 15200 11092 15252 11144
rect 16948 11092 17000 11144
rect 17316 11092 17368 11144
rect 5080 11024 5132 11076
rect 12900 11024 12952 11076
rect 18880 11024 18932 11076
rect 19156 11092 19208 11144
rect 2320 10956 2372 11008
rect 3516 10956 3568 11008
rect 3700 10999 3752 11008
rect 3700 10965 3709 10999
rect 3709 10965 3743 10999
rect 3743 10965 3752 10999
rect 3700 10956 3752 10965
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 10600 10956 10652 11008
rect 11704 10956 11756 11008
rect 12348 10956 12400 11008
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 4648 10854 4700 10906
rect 4712 10854 4764 10906
rect 4776 10854 4828 10906
rect 4840 10854 4892 10906
rect 11982 10854 12034 10906
rect 12046 10854 12098 10906
rect 12110 10854 12162 10906
rect 12174 10854 12226 10906
rect 19315 10854 19367 10906
rect 19379 10854 19431 10906
rect 19443 10854 19495 10906
rect 19507 10854 19559 10906
rect 2780 10752 2832 10804
rect 3148 10752 3200 10804
rect 4160 10752 4212 10804
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 1952 10684 2004 10736
rect 3884 10684 3936 10736
rect 5908 10684 5960 10736
rect 3148 10616 3200 10668
rect 3700 10616 3752 10668
rect 8116 10752 8168 10804
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 10876 10752 10928 10804
rect 12348 10752 12400 10804
rect 12808 10752 12860 10804
rect 15108 10752 15160 10804
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 18052 10752 18104 10804
rect 6828 10684 6880 10736
rect 7380 10684 7432 10736
rect 17040 10727 17092 10736
rect 17040 10693 17049 10727
rect 17049 10693 17083 10727
rect 17083 10693 17092 10727
rect 17040 10684 17092 10693
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7564 10616 7616 10668
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11888 10616 11940 10668
rect 12808 10616 12860 10668
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 16580 10616 16632 10668
rect 17224 10616 17276 10668
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 2320 10548 2372 10600
rect 6092 10548 6144 10600
rect 6736 10548 6788 10600
rect 15016 10548 15068 10600
rect 2228 10523 2280 10532
rect 2228 10489 2237 10523
rect 2237 10489 2271 10523
rect 2271 10489 2280 10523
rect 2228 10480 2280 10489
rect 3240 10480 3292 10532
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 6644 10480 6696 10532
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 6276 10412 6328 10464
rect 6828 10412 6880 10464
rect 10876 10523 10928 10532
rect 10876 10489 10885 10523
rect 10885 10489 10919 10523
rect 10919 10489 10928 10523
rect 10876 10480 10928 10489
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 9680 10412 9732 10464
rect 10048 10412 10100 10464
rect 10508 10412 10560 10464
rect 11152 10412 11204 10464
rect 12348 10412 12400 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 16948 10480 17000 10532
rect 19064 10752 19116 10804
rect 18512 10684 18564 10736
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 14096 10412 14148 10421
rect 15200 10412 15252 10464
rect 17316 10412 17368 10464
rect 8315 10310 8367 10362
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 15648 10310 15700 10362
rect 15712 10310 15764 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 1492 10208 1544 10260
rect 2228 10208 2280 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 2320 10140 2372 10192
rect 3148 10183 3200 10192
rect 1676 10072 1728 10124
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3148 10149 3157 10183
rect 3157 10149 3191 10183
rect 3191 10149 3200 10183
rect 3148 10140 3200 10149
rect 3424 10183 3476 10192
rect 3424 10149 3433 10183
rect 3433 10149 3467 10183
rect 3467 10149 3476 10183
rect 3424 10140 3476 10149
rect 3700 10140 3752 10192
rect 3976 10140 4028 10192
rect 5080 10140 5132 10192
rect 7288 10208 7340 10260
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 11336 10208 11388 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 16396 10208 16448 10260
rect 16580 10208 16632 10260
rect 19708 10208 19760 10260
rect 21456 10208 21508 10260
rect 6460 10183 6512 10192
rect 6460 10149 6469 10183
rect 6469 10149 6503 10183
rect 6503 10149 6512 10183
rect 6460 10140 6512 10149
rect 8024 10183 8076 10192
rect 8024 10149 8033 10183
rect 8033 10149 8067 10183
rect 8067 10149 8076 10183
rect 8024 10140 8076 10149
rect 9404 10140 9456 10192
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 11152 10140 11204 10192
rect 12716 10140 12768 10192
rect 14096 10140 14148 10192
rect 17316 10140 17368 10192
rect 3240 10072 3292 10124
rect 12900 10072 12952 10124
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 3516 10004 3568 10056
rect 4252 10004 4304 10056
rect 5540 10004 5592 10056
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 7932 10047 7984 10056
rect 1768 9936 1820 9988
rect 5908 9936 5960 9988
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 11060 10004 11112 10056
rect 16672 10072 16724 10124
rect 16948 10072 17000 10124
rect 19064 10140 19116 10192
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 7932 9868 7984 9920
rect 15752 10004 15804 10056
rect 17776 10004 17828 10056
rect 18420 10004 18472 10056
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 13820 9936 13872 9988
rect 16120 9936 16172 9988
rect 13728 9868 13780 9920
rect 14464 9868 14516 9920
rect 4648 9766 4700 9818
rect 4712 9766 4764 9818
rect 4776 9766 4828 9818
rect 4840 9766 4892 9818
rect 11982 9766 12034 9818
rect 12046 9766 12098 9818
rect 12110 9766 12162 9818
rect 12174 9766 12226 9818
rect 19315 9766 19367 9818
rect 19379 9766 19431 9818
rect 19443 9766 19495 9818
rect 19507 9766 19559 9818
rect 3976 9664 4028 9716
rect 5264 9664 5316 9716
rect 9036 9707 9088 9716
rect 9036 9673 9045 9707
rect 9045 9673 9079 9707
rect 9079 9673 9088 9707
rect 9036 9664 9088 9673
rect 1492 9596 1544 9648
rect 2136 9596 2188 9648
rect 4528 9596 4580 9648
rect 5356 9596 5408 9648
rect 6460 9596 6512 9648
rect 1584 9528 1636 9580
rect 5080 9528 5132 9580
rect 5632 9528 5684 9580
rect 8024 9528 8076 9580
rect 9956 9664 10008 9716
rect 11152 9707 11204 9716
rect 11152 9673 11161 9707
rect 11161 9673 11195 9707
rect 11195 9673 11204 9707
rect 11152 9664 11204 9673
rect 15752 9707 15804 9716
rect 15752 9673 15761 9707
rect 15761 9673 15795 9707
rect 15795 9673 15804 9707
rect 15752 9664 15804 9673
rect 16672 9664 16724 9716
rect 19064 9707 19116 9716
rect 19064 9673 19073 9707
rect 19073 9673 19107 9707
rect 19107 9673 19116 9707
rect 19064 9664 19116 9673
rect 11060 9596 11112 9648
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 13452 9596 13504 9648
rect 15476 9596 15528 9648
rect 16396 9596 16448 9648
rect 17040 9639 17092 9648
rect 14740 9528 14792 9580
rect 15384 9528 15436 9580
rect 16120 9528 16172 9580
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 18420 9596 18472 9648
rect 17592 9528 17644 9580
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 18144 9528 18196 9537
rect 18880 9528 18932 9580
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 2872 9460 2924 9512
rect 2780 9392 2832 9444
rect 3332 9460 3384 9512
rect 7748 9460 7800 9512
rect 11152 9460 11204 9512
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 21548 9460 21600 9512
rect 4528 9392 4580 9444
rect 6920 9392 6972 9444
rect 7564 9435 7616 9444
rect 7564 9401 7573 9435
rect 7573 9401 7607 9435
rect 7607 9401 7616 9435
rect 7564 9392 7616 9401
rect 8852 9392 8904 9444
rect 10508 9392 10560 9444
rect 12900 9392 12952 9444
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 15200 9435 15252 9444
rect 3148 9324 3200 9376
rect 10232 9324 10284 9376
rect 10692 9324 10744 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 14096 9324 14148 9376
rect 14464 9324 14516 9376
rect 15200 9401 15209 9435
rect 15209 9401 15243 9435
rect 15243 9401 15252 9435
rect 15200 9392 15252 9401
rect 16580 9435 16632 9444
rect 16580 9401 16589 9435
rect 16589 9401 16623 9435
rect 16623 9401 16632 9435
rect 16580 9392 16632 9401
rect 15384 9324 15436 9376
rect 17316 9324 17368 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 19524 9324 19576 9376
rect 8315 9222 8367 9274
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 15648 9222 15700 9274
rect 15712 9222 15764 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 1400 9120 1452 9172
rect 1768 9120 1820 9172
rect 3332 9120 3384 9172
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 8024 9120 8076 9172
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 11612 9163 11664 9172
rect 1676 9052 1728 9104
rect 3884 9052 3936 9104
rect 4252 9095 4304 9104
rect 4252 9061 4261 9095
rect 4261 9061 4295 9095
rect 4295 9061 4304 9095
rect 4252 9052 4304 9061
rect 5448 9052 5500 9104
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 5632 9027 5684 9036
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 6644 8984 6696 9036
rect 7104 9052 7156 9104
rect 7564 9052 7616 9104
rect 9864 9052 9916 9104
rect 11612 9129 11621 9163
rect 11621 9129 11655 9163
rect 11655 9129 11664 9163
rect 11612 9120 11664 9129
rect 13636 9120 13688 9172
rect 14740 9163 14792 9172
rect 10692 9095 10744 9104
rect 10692 9061 10701 9095
rect 10701 9061 10735 9095
rect 10735 9061 10744 9095
rect 10692 9052 10744 9061
rect 11888 9052 11940 9104
rect 13176 9052 13228 9104
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 16580 9120 16632 9172
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 18144 9163 18196 9172
rect 18144 9129 18153 9163
rect 18153 9129 18187 9163
rect 18187 9129 18196 9163
rect 18144 9120 18196 9129
rect 13820 9095 13872 9104
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 14556 9052 14608 9104
rect 15016 9095 15068 9104
rect 15016 9061 15025 9095
rect 15025 9061 15059 9095
rect 15059 9061 15068 9095
rect 15016 9052 15068 9061
rect 15384 9052 15436 9104
rect 17316 9052 17368 9104
rect 18788 9095 18840 9104
rect 18788 9061 18797 9095
rect 18797 9061 18831 9095
rect 18831 9061 18840 9095
rect 18788 9052 18840 9061
rect 7932 8984 7984 9036
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 2228 8916 2280 8968
rect 2688 8916 2740 8968
rect 3332 8848 3384 8900
rect 2136 8780 2188 8832
rect 3240 8780 3292 8832
rect 3884 8780 3936 8832
rect 7840 8916 7892 8968
rect 10600 8916 10652 8968
rect 6920 8848 6972 8900
rect 11152 8891 11204 8900
rect 11152 8857 11161 8891
rect 11161 8857 11195 8891
rect 11195 8857 11204 8891
rect 15108 8916 15160 8968
rect 15844 8916 15896 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 17868 8916 17920 8968
rect 19524 8916 19576 8968
rect 11152 8848 11204 8857
rect 12624 8848 12676 8900
rect 14648 8848 14700 8900
rect 19064 8848 19116 8900
rect 6000 8780 6052 8832
rect 6368 8823 6420 8832
rect 6368 8789 6377 8823
rect 6377 8789 6411 8823
rect 6411 8789 6420 8823
rect 6368 8780 6420 8789
rect 11796 8780 11848 8832
rect 12716 8780 12768 8832
rect 4648 8678 4700 8730
rect 4712 8678 4764 8730
rect 4776 8678 4828 8730
rect 4840 8678 4892 8730
rect 11982 8678 12034 8730
rect 12046 8678 12098 8730
rect 12110 8678 12162 8730
rect 12174 8678 12226 8730
rect 19315 8678 19367 8730
rect 19379 8678 19431 8730
rect 19443 8678 19495 8730
rect 19507 8678 19559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2044 8576 2096 8628
rect 2964 8576 3016 8628
rect 4252 8576 4304 8628
rect 6276 8576 6328 8628
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 10232 8619 10284 8628
rect 10232 8585 10241 8619
rect 10241 8585 10275 8619
rect 10275 8585 10284 8619
rect 10232 8576 10284 8585
rect 10416 8576 10468 8628
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 16856 8576 16908 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 18788 8576 18840 8628
rect 19616 8619 19668 8628
rect 19616 8585 19625 8619
rect 19625 8585 19659 8619
rect 19659 8585 19668 8619
rect 19616 8576 19668 8585
rect 1584 8440 1636 8492
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 6092 8508 6144 8560
rect 6368 8508 6420 8560
rect 5448 8440 5500 8492
rect 7472 8440 7524 8492
rect 9128 8440 9180 8492
rect 10140 8440 10192 8492
rect 10600 8440 10652 8492
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 13268 8440 13320 8492
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 12532 8372 12584 8424
rect 15016 8440 15068 8492
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 3332 8304 3384 8356
rect 4068 8236 4120 8288
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 7564 8304 7616 8356
rect 5080 8236 5132 8288
rect 6000 8279 6052 8288
rect 6000 8245 6009 8279
rect 6009 8245 6043 8279
rect 6043 8245 6052 8279
rect 6000 8236 6052 8245
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 9036 8279 9088 8288
rect 7472 8236 7524 8245
rect 9036 8245 9045 8279
rect 9045 8245 9079 8279
rect 9079 8245 9088 8279
rect 10416 8304 10468 8356
rect 9036 8236 9088 8245
rect 9772 8236 9824 8288
rect 10140 8236 10192 8288
rect 11888 8236 11940 8288
rect 13452 8236 13504 8288
rect 13636 8236 13688 8288
rect 13820 8236 13872 8288
rect 15476 8236 15528 8288
rect 17316 8236 17368 8288
rect 18512 8236 18564 8288
rect 19064 8304 19116 8356
rect 8315 8134 8367 8186
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 15648 8134 15700 8186
rect 15712 8134 15764 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 1400 8032 1452 8084
rect 2780 8032 2832 8084
rect 1676 8007 1728 8016
rect 1676 7973 1685 8007
rect 1685 7973 1719 8007
rect 1719 7973 1728 8007
rect 1676 7964 1728 7973
rect 3332 7964 3384 8016
rect 2412 7896 2464 7948
rect 4712 8032 4764 8084
rect 5080 8032 5132 8084
rect 6276 8032 6328 8084
rect 8852 8032 8904 8084
rect 9128 8032 9180 8084
rect 9312 8032 9364 8084
rect 10232 8032 10284 8084
rect 13912 8032 13964 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16488 8032 16540 8084
rect 16948 8032 17000 8084
rect 17500 8032 17552 8084
rect 7564 7964 7616 8016
rect 11796 7964 11848 8016
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 15476 8007 15528 8016
rect 13820 7964 13872 7973
rect 15476 7973 15485 8007
rect 15485 7973 15519 8007
rect 15519 7973 15528 8007
rect 15476 7964 15528 7973
rect 17316 7964 17368 8016
rect 18512 7964 18564 8016
rect 4528 7896 4580 7948
rect 9772 7939 9824 7948
rect 9772 7905 9781 7939
rect 9781 7905 9815 7939
rect 9815 7905 9824 7939
rect 9772 7896 9824 7905
rect 6276 7828 6328 7880
rect 9128 7828 9180 7880
rect 9588 7828 9640 7880
rect 12624 7896 12676 7948
rect 16764 7896 16816 7948
rect 18420 7896 18472 7948
rect 1308 7692 1360 7744
rect 5356 7692 5408 7744
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 14832 7828 14884 7880
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 15200 7760 15252 7812
rect 17960 7828 18012 7880
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 18880 7828 18932 7880
rect 7012 7692 7064 7744
rect 7472 7692 7524 7744
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 4648 7590 4700 7642
rect 4712 7590 4764 7642
rect 4776 7590 4828 7642
rect 4840 7590 4892 7642
rect 11982 7590 12034 7642
rect 12046 7590 12098 7642
rect 12110 7590 12162 7642
rect 12174 7590 12226 7642
rect 19315 7590 19367 7642
rect 19379 7590 19431 7642
rect 19443 7590 19495 7642
rect 19507 7590 19559 7642
rect 1768 7488 1820 7540
rect 3332 7488 3384 7540
rect 4528 7488 4580 7540
rect 10048 7488 10100 7540
rect 12808 7531 12860 7540
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 15476 7488 15528 7540
rect 16304 7488 16356 7540
rect 16764 7488 16816 7540
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 18512 7488 18564 7540
rect 1308 7352 1360 7404
rect 6092 7420 6144 7472
rect 11888 7420 11940 7472
rect 13452 7420 13504 7472
rect 6000 7352 6052 7404
rect 6920 7352 6972 7404
rect 7288 7352 7340 7404
rect 11152 7352 11204 7404
rect 12348 7352 12400 7404
rect 18788 7420 18840 7472
rect 8576 7284 8628 7336
rect 2964 7216 3016 7268
rect 3332 7259 3384 7268
rect 3332 7225 3341 7259
rect 3341 7225 3375 7259
rect 3375 7225 3384 7259
rect 3332 7216 3384 7225
rect 5356 7259 5408 7268
rect 5356 7225 5365 7259
rect 5365 7225 5399 7259
rect 5399 7225 5408 7259
rect 5356 7216 5408 7225
rect 6920 7259 6972 7268
rect 1676 7148 1728 7200
rect 5080 7148 5132 7200
rect 6276 7148 6328 7200
rect 6920 7225 6929 7259
rect 6929 7225 6963 7259
rect 6963 7225 6972 7259
rect 6920 7216 6972 7225
rect 7012 7259 7064 7268
rect 7012 7225 7021 7259
rect 7021 7225 7055 7259
rect 7055 7225 7064 7259
rect 7012 7216 7064 7225
rect 7564 7216 7616 7268
rect 10508 7259 10560 7268
rect 10508 7225 10517 7259
rect 10517 7225 10551 7259
rect 10551 7225 10560 7259
rect 10508 7216 10560 7225
rect 9036 7148 9088 7200
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 12348 7216 12400 7268
rect 14004 7284 14056 7336
rect 16488 7327 16540 7336
rect 16488 7293 16497 7327
rect 16497 7293 16531 7327
rect 16531 7293 16540 7327
rect 16488 7284 16540 7293
rect 18696 7352 18748 7404
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 14464 7216 14516 7268
rect 18144 7216 18196 7268
rect 13268 7148 13320 7200
rect 13636 7148 13688 7200
rect 17316 7191 17368 7200
rect 17316 7157 17325 7191
rect 17325 7157 17359 7191
rect 17359 7157 17368 7191
rect 17316 7148 17368 7157
rect 18420 7148 18472 7200
rect 8315 7046 8367 7098
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 15648 7046 15700 7098
rect 15712 7046 15764 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 6920 6944 6972 6996
rect 7656 6944 7708 6996
rect 8944 6944 8996 6996
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 11888 6944 11940 6996
rect 13636 6944 13688 6996
rect 13820 6944 13872 6996
rect 14004 6944 14056 6996
rect 17408 6944 17460 6996
rect 18512 6944 18564 6996
rect 18696 6944 18748 6996
rect 1952 6919 2004 6928
rect 1952 6885 1961 6919
rect 1961 6885 1995 6919
rect 1995 6885 2004 6919
rect 1952 6876 2004 6885
rect 2228 6919 2280 6928
rect 2228 6885 2237 6919
rect 2237 6885 2271 6919
rect 2271 6885 2280 6919
rect 2228 6876 2280 6885
rect 3332 6876 3384 6928
rect 3792 6876 3844 6928
rect 1584 6808 1636 6860
rect 3884 6808 3936 6860
rect 5080 6876 5132 6928
rect 6644 6876 6696 6928
rect 12900 6919 12952 6928
rect 12900 6885 12909 6919
rect 12909 6885 12943 6919
rect 12943 6885 12952 6919
rect 12900 6876 12952 6885
rect 4160 6808 4212 6860
rect 6092 6851 6144 6860
rect 6092 6817 6101 6851
rect 6101 6817 6135 6851
rect 6135 6817 6144 6851
rect 6092 6808 6144 6817
rect 8668 6808 8720 6860
rect 8852 6808 8904 6860
rect 10876 6808 10928 6860
rect 11796 6851 11848 6860
rect 11796 6817 11805 6851
rect 11805 6817 11839 6851
rect 11839 6817 11848 6851
rect 11796 6808 11848 6817
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 15292 6808 15344 6860
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 16304 6808 16356 6860
rect 18788 6876 18840 6928
rect 17408 6808 17460 6860
rect 1676 6740 1728 6792
rect 5816 6740 5868 6792
rect 6368 6740 6420 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 10692 6740 10744 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 17776 6740 17828 6792
rect 2964 6672 3016 6724
rect 3332 6604 3384 6656
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 6184 6672 6236 6724
rect 7196 6672 7248 6724
rect 11060 6672 11112 6724
rect 14188 6672 14240 6724
rect 15384 6672 15436 6724
rect 18880 6740 18932 6792
rect 19616 6672 19668 6724
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 10600 6604 10652 6656
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 16488 6604 16540 6656
rect 4648 6502 4700 6554
rect 4712 6502 4764 6554
rect 4776 6502 4828 6554
rect 4840 6502 4892 6554
rect 11982 6502 12034 6554
rect 12046 6502 12098 6554
rect 12110 6502 12162 6554
rect 12174 6502 12226 6554
rect 19315 6502 19367 6554
rect 19379 6502 19431 6554
rect 19443 6502 19495 6554
rect 19507 6502 19559 6554
rect 2964 6400 3016 6452
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 3332 6400 3384 6409
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 8668 6400 8720 6452
rect 8852 6400 8904 6452
rect 13452 6443 13504 6452
rect 13452 6409 13461 6443
rect 13461 6409 13495 6443
rect 13495 6409 13504 6443
rect 13452 6400 13504 6409
rect 15292 6400 15344 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 17960 6400 18012 6452
rect 18788 6400 18840 6452
rect 3240 6332 3292 6384
rect 7012 6332 7064 6384
rect 7932 6375 7984 6384
rect 7932 6341 7941 6375
rect 7941 6341 7975 6375
rect 7975 6341 7984 6375
rect 11152 6375 11204 6384
rect 7932 6332 7984 6341
rect 4160 6264 4212 6316
rect 4988 6264 5040 6316
rect 7196 6264 7248 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 11152 6341 11161 6375
rect 11161 6341 11195 6375
rect 11195 6341 11204 6375
rect 11152 6332 11204 6341
rect 13360 6332 13412 6384
rect 15936 6375 15988 6384
rect 15936 6341 15945 6375
rect 15945 6341 15979 6375
rect 15979 6341 15988 6375
rect 15936 6332 15988 6341
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 1584 6060 1636 6112
rect 5080 6128 5132 6180
rect 5632 6128 5684 6180
rect 6828 6128 6880 6180
rect 7472 6171 7524 6180
rect 7472 6137 7481 6171
rect 7481 6137 7515 6171
rect 7515 6137 7524 6171
rect 7472 6128 7524 6137
rect 9036 6171 9088 6180
rect 9036 6137 9045 6171
rect 9045 6137 9079 6171
rect 9079 6137 9088 6171
rect 9036 6128 9088 6137
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 6000 6060 6052 6112
rect 8944 6060 8996 6112
rect 9772 6128 9824 6180
rect 10600 6196 10652 6248
rect 10876 6128 10928 6180
rect 11704 6196 11756 6248
rect 12532 6239 12584 6248
rect 12072 6128 12124 6180
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 12808 6196 12860 6248
rect 13728 6196 13780 6248
rect 14832 6239 14884 6248
rect 14832 6205 14841 6239
rect 14841 6205 14875 6239
rect 14875 6205 14884 6239
rect 14832 6196 14884 6205
rect 15476 6196 15528 6248
rect 19064 6264 19116 6316
rect 16304 6128 16356 6180
rect 16488 6171 16540 6180
rect 16488 6137 16497 6171
rect 16497 6137 16531 6171
rect 16531 6137 16540 6171
rect 16488 6128 16540 6137
rect 16764 6128 16816 6180
rect 17960 6128 18012 6180
rect 18972 6128 19024 6180
rect 19340 6171 19392 6180
rect 19340 6137 19349 6171
rect 19349 6137 19383 6171
rect 19383 6137 19392 6171
rect 19340 6128 19392 6137
rect 11704 6060 11756 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12348 6060 12400 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 8315 5958 8367 6010
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 15648 5958 15700 6010
rect 15712 5958 15764 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 3056 5856 3108 5908
rect 3700 5856 3752 5908
rect 3884 5899 3936 5908
rect 3884 5865 3893 5899
rect 3893 5865 3927 5899
rect 3927 5865 3936 5899
rect 3884 5856 3936 5865
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 5448 5856 5500 5908
rect 6184 5856 6236 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 2412 5788 2464 5840
rect 3792 5788 3844 5840
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 4988 5788 5040 5840
rect 8208 5856 8260 5908
rect 8852 5856 8904 5908
rect 9036 5899 9088 5908
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 9312 5856 9364 5908
rect 10876 5856 10928 5908
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 14924 5856 14976 5908
rect 16120 5856 16172 5908
rect 16304 5856 16356 5908
rect 17960 5899 18012 5908
rect 6828 5831 6880 5840
rect 6828 5797 6837 5831
rect 6837 5797 6871 5831
rect 6871 5797 6880 5831
rect 6828 5788 6880 5797
rect 4252 5720 4304 5772
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 3608 5652 3660 5704
rect 3792 5652 3844 5704
rect 5816 5652 5868 5704
rect 7748 5720 7800 5772
rect 12072 5788 12124 5840
rect 8300 5720 8352 5772
rect 9128 5720 9180 5772
rect 9496 5720 9548 5772
rect 9772 5720 9824 5772
rect 11336 5763 11388 5772
rect 6092 5652 6144 5704
rect 6736 5652 6788 5704
rect 6920 5652 6972 5704
rect 8852 5652 8904 5704
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 11428 5720 11480 5772
rect 11612 5720 11664 5772
rect 11704 5720 11756 5772
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 14464 5788 14516 5840
rect 16764 5788 16816 5840
rect 17960 5865 17969 5899
rect 17969 5865 18003 5899
rect 18003 5865 18012 5899
rect 17960 5856 18012 5865
rect 18144 5856 18196 5908
rect 17408 5831 17460 5840
rect 17408 5797 17411 5831
rect 17411 5797 17445 5831
rect 17445 5797 17460 5831
rect 17408 5788 17460 5797
rect 17868 5788 17920 5840
rect 19156 5788 19208 5840
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 14004 5695 14056 5704
rect 12256 5652 12308 5661
rect 14004 5661 14013 5695
rect 14013 5661 14047 5695
rect 14047 5661 14056 5695
rect 14004 5652 14056 5661
rect 15200 5652 15252 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 19064 5652 19116 5704
rect 19340 5695 19392 5704
rect 19340 5661 19349 5695
rect 19349 5661 19383 5695
rect 19383 5661 19392 5695
rect 19340 5652 19392 5661
rect 1676 5584 1728 5636
rect 2320 5516 2372 5568
rect 7288 5627 7340 5636
rect 7288 5593 7297 5627
rect 7297 5593 7331 5627
rect 7331 5593 7340 5627
rect 7288 5584 7340 5593
rect 6000 5516 6052 5568
rect 11612 5584 11664 5636
rect 14832 5584 14884 5636
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 16028 5516 16080 5568
rect 18972 5516 19024 5568
rect 4648 5414 4700 5466
rect 4712 5414 4764 5466
rect 4776 5414 4828 5466
rect 4840 5414 4892 5466
rect 11982 5414 12034 5466
rect 12046 5414 12098 5466
rect 12110 5414 12162 5466
rect 12174 5414 12226 5466
rect 19315 5414 19367 5466
rect 19379 5414 19431 5466
rect 19443 5414 19495 5466
rect 19507 5414 19559 5466
rect 2780 5312 2832 5364
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 5080 5312 5132 5364
rect 1952 5244 2004 5296
rect 8944 5312 8996 5364
rect 9772 5312 9824 5364
rect 10508 5312 10560 5364
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 11336 5312 11388 5364
rect 12348 5312 12400 5364
rect 14188 5312 14240 5364
rect 14464 5355 14516 5364
rect 14464 5321 14473 5355
rect 14473 5321 14507 5355
rect 14507 5321 14516 5355
rect 14464 5312 14516 5321
rect 15292 5312 15344 5364
rect 18972 5355 19024 5364
rect 18972 5321 18981 5355
rect 18981 5321 19015 5355
rect 19015 5321 19024 5355
rect 18972 5312 19024 5321
rect 6552 5244 6604 5296
rect 6828 5244 6880 5296
rect 2320 5108 2372 5160
rect 2412 5108 2464 5160
rect 3608 5176 3660 5228
rect 4068 5176 4120 5228
rect 4528 5176 4580 5228
rect 5172 5176 5224 5228
rect 6000 5176 6052 5228
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 3700 5151 3752 5160
rect 2780 5040 2832 5092
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 6736 5108 6788 5160
rect 3792 5040 3844 5092
rect 5080 5040 5132 5092
rect 8208 5244 8260 5296
rect 9404 5244 9456 5296
rect 11796 5244 11848 5296
rect 16028 5287 16080 5296
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 8300 5176 8352 5228
rect 9128 5176 9180 5228
rect 10968 5176 11020 5228
rect 12072 5176 12124 5228
rect 12348 5176 12400 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 13360 5176 13412 5228
rect 7748 5108 7800 5160
rect 11612 5108 11664 5160
rect 3424 4972 3476 5024
rect 8668 5040 8720 5092
rect 8852 5040 8904 5092
rect 10968 5083 11020 5092
rect 10968 5049 10977 5083
rect 10977 5049 11011 5083
rect 11011 5049 11020 5083
rect 10968 5040 11020 5049
rect 7196 4972 7248 5024
rect 7564 4972 7616 5024
rect 11704 4972 11756 5024
rect 13636 5083 13688 5092
rect 13636 5049 13645 5083
rect 13645 5049 13679 5083
rect 13679 5049 13688 5083
rect 16028 5253 16037 5287
rect 16037 5253 16071 5287
rect 16071 5253 16080 5287
rect 16028 5244 16080 5253
rect 18880 5244 18932 5296
rect 14924 5108 14976 5160
rect 16580 5176 16632 5228
rect 18144 5176 18196 5228
rect 15108 5108 15160 5160
rect 19432 5108 19484 5160
rect 13636 5040 13688 5049
rect 14740 5040 14792 5092
rect 15200 5040 15252 5092
rect 16580 5083 16632 5092
rect 16580 5049 16589 5083
rect 16589 5049 16623 5083
rect 16623 5049 16632 5083
rect 16580 5040 16632 5049
rect 14280 4972 14332 5024
rect 14832 5015 14884 5024
rect 14832 4981 14841 5015
rect 14841 4981 14875 5015
rect 14875 4981 14884 5015
rect 14832 4972 14884 4981
rect 17868 5015 17920 5024
rect 17868 4981 17877 5015
rect 17877 4981 17911 5015
rect 17911 4981 17920 5015
rect 17868 4972 17920 4981
rect 19248 5015 19300 5024
rect 19248 4981 19257 5015
rect 19257 4981 19291 5015
rect 19291 4981 19300 5015
rect 19248 4972 19300 4981
rect 8315 4870 8367 4922
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 15648 4870 15700 4922
rect 15712 4870 15764 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 1676 4768 1728 4820
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 2688 4768 2740 4820
rect 2872 4768 2924 4820
rect 3700 4768 3752 4820
rect 3976 4768 4028 4820
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 5448 4811 5500 4820
rect 5448 4777 5457 4811
rect 5457 4777 5491 4811
rect 5491 4777 5500 4811
rect 5448 4768 5500 4777
rect 5632 4768 5684 4820
rect 6552 4811 6604 4820
rect 6552 4777 6561 4811
rect 6561 4777 6595 4811
rect 6595 4777 6604 4811
rect 6552 4768 6604 4777
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 3148 4743 3200 4752
rect 2044 4632 2096 4684
rect 2688 4632 2740 4684
rect 3148 4709 3157 4743
rect 3157 4709 3191 4743
rect 3191 4709 3200 4743
rect 3148 4700 3200 4709
rect 3424 4632 3476 4684
rect 3792 4632 3844 4684
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4252 4700 4304 4752
rect 5540 4700 5592 4752
rect 6460 4700 6512 4752
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 5724 4632 5776 4684
rect 2320 4539 2372 4548
rect 2320 4505 2329 4539
rect 2329 4505 2363 4539
rect 2363 4505 2372 4539
rect 2320 4496 2372 4505
rect 3976 4564 4028 4616
rect 7656 4768 7708 4820
rect 7932 4768 7984 4820
rect 8668 4768 8720 4820
rect 10968 4768 11020 4820
rect 11704 4768 11756 4820
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 15476 4768 15528 4820
rect 16212 4768 16264 4820
rect 16580 4811 16632 4820
rect 16580 4777 16589 4811
rect 16589 4777 16623 4811
rect 16623 4777 16632 4811
rect 16580 4768 16632 4777
rect 19248 4768 19300 4820
rect 7564 4743 7616 4752
rect 7564 4709 7573 4743
rect 7573 4709 7607 4743
rect 7607 4709 7616 4743
rect 7564 4700 7616 4709
rect 7840 4700 7892 4752
rect 8208 4700 8260 4752
rect 8944 4700 8996 4752
rect 11244 4743 11296 4752
rect 11244 4709 11253 4743
rect 11253 4709 11287 4743
rect 11287 4709 11296 4743
rect 11244 4700 11296 4709
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 13452 4700 13504 4752
rect 15200 4700 15252 4752
rect 9956 4632 10008 4684
rect 12440 4632 12492 4684
rect 14004 4632 14056 4684
rect 15016 4632 15068 4684
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 11152 4607 11204 4616
rect 2964 4496 3016 4548
rect 1676 4428 1728 4480
rect 2504 4428 2556 4480
rect 2780 4428 2832 4480
rect 5448 4428 5500 4480
rect 7656 4496 7708 4548
rect 9680 4496 9732 4548
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 9772 4428 9824 4480
rect 10140 4428 10192 4480
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 15384 4564 15436 4616
rect 17868 4700 17920 4752
rect 18604 4700 18656 4752
rect 20076 4700 20128 4752
rect 21548 4700 21600 4752
rect 19432 4632 19484 4684
rect 18144 4564 18196 4616
rect 10784 4496 10836 4548
rect 11796 4496 11848 4548
rect 12532 4428 12584 4480
rect 13544 4471 13596 4480
rect 13544 4437 13553 4471
rect 13553 4437 13587 4471
rect 13587 4437 13596 4471
rect 14832 4496 14884 4548
rect 16028 4496 16080 4548
rect 13544 4428 13596 4437
rect 15936 4428 15988 4480
rect 16856 4428 16908 4480
rect 17132 4428 17184 4480
rect 4648 4326 4700 4378
rect 4712 4326 4764 4378
rect 4776 4326 4828 4378
rect 4840 4326 4892 4378
rect 11982 4326 12034 4378
rect 12046 4326 12098 4378
rect 12110 4326 12162 4378
rect 12174 4326 12226 4378
rect 19315 4326 19367 4378
rect 19379 4326 19431 4378
rect 19443 4326 19495 4378
rect 19507 4326 19559 4378
rect 1492 4088 1544 4140
rect 3148 4199 3200 4208
rect 3148 4165 3157 4199
rect 3157 4165 3191 4199
rect 3191 4165 3200 4199
rect 3148 4156 3200 4165
rect 3792 4224 3844 4276
rect 4068 4156 4120 4208
rect 4436 4156 4488 4208
rect 8208 4224 8260 4276
rect 8944 4224 8996 4276
rect 9956 4224 10008 4276
rect 10508 4224 10560 4276
rect 5264 4156 5316 4208
rect 7196 4156 7248 4208
rect 9772 4156 9824 4208
rect 11244 4156 11296 4208
rect 11704 4224 11756 4276
rect 12624 4224 12676 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 15936 4224 15988 4276
rect 17960 4224 18012 4276
rect 19156 4267 19208 4276
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 19616 4224 19668 4276
rect 20076 4267 20128 4276
rect 20076 4233 20085 4267
rect 20085 4233 20119 4267
rect 20119 4233 20128 4267
rect 20076 4224 20128 4233
rect 2136 4088 2188 4140
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 2412 4020 2464 4072
rect 2872 4020 2924 4072
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 3700 4020 3752 4072
rect 6276 4088 6328 4140
rect 5448 4063 5500 4072
rect 2228 3952 2280 4004
rect 3608 3952 3660 4004
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 7656 4088 7708 4140
rect 5172 3952 5224 4004
rect 11796 4088 11848 4140
rect 12992 4088 13044 4140
rect 10876 4020 10928 4072
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 8668 3995 8720 4004
rect 3884 3884 3936 3936
rect 4344 3884 4396 3936
rect 6460 3884 6512 3936
rect 7012 3884 7064 3936
rect 7840 3884 7892 3936
rect 8668 3961 8677 3995
rect 8677 3961 8711 3995
rect 8711 3961 8720 3995
rect 8668 3952 8720 3961
rect 9680 3952 9732 4004
rect 10140 3952 10192 4004
rect 12624 3995 12676 4004
rect 12624 3961 12633 3995
rect 12633 3961 12667 3995
rect 12667 3961 12676 3995
rect 12624 3952 12676 3961
rect 14096 3952 14148 4004
rect 14648 3952 14700 4004
rect 16396 4020 16448 4072
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 16580 3952 16632 4004
rect 17316 3952 17368 4004
rect 18144 3952 18196 4004
rect 18788 3995 18840 4004
rect 18788 3961 18797 3995
rect 18797 3961 18831 3995
rect 18831 3961 18840 3995
rect 18788 3952 18840 3961
rect 18880 3952 18932 4004
rect 8760 3884 8812 3936
rect 9496 3884 9548 3936
rect 11520 3884 11572 3936
rect 13452 3884 13504 3936
rect 15108 3884 15160 3936
rect 15476 3884 15528 3936
rect 16028 3927 16080 3936
rect 16028 3893 16037 3927
rect 16037 3893 16071 3927
rect 16071 3893 16080 3927
rect 16028 3884 16080 3893
rect 16856 3884 16908 3936
rect 8315 3782 8367 3834
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 15648 3782 15700 3834
rect 15712 3782 15764 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 5172 3680 5224 3732
rect 5540 3723 5592 3732
rect 5540 3689 5549 3723
rect 5549 3689 5583 3723
rect 5583 3689 5592 3723
rect 5540 3680 5592 3689
rect 5632 3680 5684 3732
rect 6368 3680 6420 3732
rect 7564 3680 7616 3732
rect 8760 3680 8812 3732
rect 9312 3680 9364 3732
rect 10140 3680 10192 3732
rect 11336 3680 11388 3732
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 12348 3680 12400 3732
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 15016 3723 15068 3732
rect 15016 3689 15025 3723
rect 15025 3689 15059 3723
rect 15059 3689 15068 3723
rect 15016 3680 15068 3689
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 16488 3680 16540 3732
rect 18052 3680 18104 3732
rect 18236 3723 18288 3732
rect 18236 3689 18245 3723
rect 18245 3689 18279 3723
rect 18279 3689 18288 3723
rect 18236 3680 18288 3689
rect 18788 3680 18840 3732
rect 2780 3612 2832 3664
rect 3516 3612 3568 3664
rect 2412 3587 2464 3596
rect 2412 3553 2421 3587
rect 2421 3553 2455 3587
rect 2455 3553 2464 3587
rect 2412 3544 2464 3553
rect 1676 3476 1728 3528
rect 3792 3544 3844 3596
rect 4068 3544 4120 3596
rect 5448 3612 5500 3664
rect 6184 3655 6236 3664
rect 6184 3621 6193 3655
rect 6193 3621 6227 3655
rect 6227 3621 6236 3655
rect 6184 3612 6236 3621
rect 6276 3655 6328 3664
rect 6276 3621 6285 3655
rect 6285 3621 6319 3655
rect 6319 3621 6328 3655
rect 6276 3612 6328 3621
rect 7840 3612 7892 3664
rect 5356 3544 5408 3596
rect 7380 3544 7432 3596
rect 10784 3544 10836 3596
rect 11520 3612 11572 3664
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 15200 3612 15252 3664
rect 15384 3655 15436 3664
rect 15384 3621 15393 3655
rect 15393 3621 15427 3655
rect 15427 3621 15436 3655
rect 15384 3612 15436 3621
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 16948 3612 17000 3664
rect 16580 3544 16632 3596
rect 16856 3544 16908 3596
rect 18972 3655 19024 3664
rect 18972 3621 18981 3655
rect 18981 3621 19015 3655
rect 19015 3621 19024 3655
rect 18972 3612 19024 3621
rect 6920 3476 6972 3528
rect 7104 3476 7156 3528
rect 8116 3476 8168 3528
rect 2596 3408 2648 3460
rect 3056 3408 3108 3460
rect 3148 3408 3200 3460
rect 7748 3408 7800 3460
rect 12716 3476 12768 3528
rect 14832 3476 14884 3528
rect 17316 3476 17368 3528
rect 19156 3519 19208 3528
rect 10784 3408 10836 3460
rect 12624 3408 12676 3460
rect 16672 3408 16724 3460
rect 2780 3340 2832 3392
rect 3332 3340 3384 3392
rect 7472 3340 7524 3392
rect 10416 3340 10468 3392
rect 10692 3383 10744 3392
rect 10692 3349 10701 3383
rect 10701 3349 10735 3383
rect 10735 3349 10744 3383
rect 10692 3340 10744 3349
rect 17132 3408 17184 3460
rect 19156 3485 19165 3519
rect 19165 3485 19199 3519
rect 19199 3485 19208 3519
rect 19156 3476 19208 3485
rect 19064 3408 19116 3460
rect 20076 3340 20128 3392
rect 4648 3238 4700 3290
rect 4712 3238 4764 3290
rect 4776 3238 4828 3290
rect 4840 3238 4892 3290
rect 11982 3238 12034 3290
rect 12046 3238 12098 3290
rect 12110 3238 12162 3290
rect 12174 3238 12226 3290
rect 19315 3238 19367 3290
rect 19379 3238 19431 3290
rect 19443 3238 19495 3290
rect 19507 3238 19559 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 5356 3136 5408 3188
rect 5448 3136 5500 3188
rect 10140 3136 10192 3188
rect 10784 3136 10836 3188
rect 2780 3068 2832 3120
rect 3516 3068 3568 3120
rect 3884 3068 3936 3120
rect 10692 3068 10744 3120
rect 4436 3000 4488 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 9312 3000 9364 3052
rect 1768 2932 1820 2984
rect 2320 2932 2372 2984
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 3516 2932 3568 2984
rect 3608 2932 3660 2984
rect 1860 2864 1912 2916
rect 6460 2932 6512 2984
rect 5448 2796 5500 2848
rect 6276 2864 6328 2916
rect 7472 2907 7524 2916
rect 7472 2873 7481 2907
rect 7481 2873 7515 2907
rect 7515 2873 7524 2907
rect 7472 2864 7524 2873
rect 7840 2864 7892 2916
rect 10692 2864 10744 2916
rect 11520 3136 11572 3188
rect 11796 3136 11848 3188
rect 13544 3179 13596 3188
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13544 3136 13596 3145
rect 15476 3136 15528 3188
rect 16580 3136 16632 3188
rect 17776 3179 17828 3188
rect 15936 3068 15988 3120
rect 11612 3000 11664 3052
rect 12348 3000 12400 3052
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 16948 3000 17000 3052
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18972 3136 19024 3188
rect 19064 3111 19116 3120
rect 19064 3077 19073 3111
rect 19073 3077 19107 3111
rect 19107 3077 19116 3111
rect 19064 3068 19116 3077
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 11428 2932 11480 2984
rect 15292 2932 15344 2984
rect 18144 3000 18196 3052
rect 15108 2864 15160 2916
rect 16856 2864 16908 2916
rect 14556 2796 14608 2848
rect 16488 2839 16540 2848
rect 16488 2805 16497 2839
rect 16497 2805 16531 2839
rect 16531 2805 16540 2839
rect 16488 2796 16540 2805
rect 20076 2975 20128 2984
rect 17776 2864 17828 2916
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 8315 2694 8367 2746
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 15648 2694 15700 2746
rect 15712 2694 15764 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 2412 2592 2464 2644
rect 2872 2592 2924 2644
rect 3056 2592 3108 2644
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 5264 2592 5316 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 6460 2592 6512 2644
rect 5448 2567 5500 2576
rect 1952 2456 2004 2508
rect 2412 2499 2464 2508
rect 2412 2465 2421 2499
rect 2421 2465 2455 2499
rect 2455 2465 2464 2499
rect 2412 2456 2464 2465
rect 2964 2456 3016 2508
rect 3148 2499 3200 2508
rect 3148 2465 3157 2499
rect 3157 2465 3191 2499
rect 3191 2465 3200 2499
rect 3148 2456 3200 2465
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5448 2533 5457 2567
rect 5457 2533 5491 2567
rect 5491 2533 5500 2567
rect 5448 2524 5500 2533
rect 7012 2524 7064 2576
rect 7472 2592 7524 2644
rect 7932 2592 7984 2644
rect 9220 2592 9272 2644
rect 10692 2635 10744 2644
rect 10692 2601 10701 2635
rect 10701 2601 10735 2635
rect 10735 2601 10744 2635
rect 10692 2592 10744 2601
rect 11704 2635 11756 2644
rect 11704 2601 11713 2635
rect 11713 2601 11747 2635
rect 11747 2601 11756 2635
rect 11704 2592 11756 2601
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 13084 2635 13136 2644
rect 13084 2601 13093 2635
rect 13093 2601 13127 2635
rect 13127 2601 13136 2635
rect 13084 2592 13136 2601
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 14556 2635 14608 2644
rect 13452 2592 13504 2601
rect 7748 2524 7800 2576
rect 8116 2567 8168 2576
rect 8116 2533 8125 2567
rect 8125 2533 8159 2567
rect 8159 2533 8168 2567
rect 8116 2524 8168 2533
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 15292 2635 15344 2644
rect 15292 2601 15301 2635
rect 15301 2601 15335 2635
rect 15335 2601 15344 2635
rect 15292 2592 15344 2601
rect 16120 2635 16172 2644
rect 16120 2601 16129 2635
rect 16129 2601 16163 2635
rect 16163 2601 16172 2635
rect 16120 2592 16172 2601
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 17776 2592 17828 2644
rect 16488 2567 16540 2576
rect 16488 2533 16497 2567
rect 16497 2533 16531 2567
rect 16531 2533 16540 2567
rect 16488 2524 16540 2533
rect 17224 2524 17276 2576
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 9128 2499 9180 2508
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 9128 2456 9180 2465
rect 9864 2499 9916 2508
rect 9864 2465 9882 2499
rect 9882 2465 9916 2499
rect 9864 2456 9916 2465
rect 13084 2388 13136 2440
rect 16120 2388 16172 2440
rect 16948 2363 17000 2372
rect 16948 2329 16957 2363
rect 16957 2329 16991 2363
rect 16991 2329 17000 2363
rect 16948 2320 17000 2329
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 12992 2252 13044 2304
rect 19156 2252 19208 2304
rect 4648 2150 4700 2202
rect 4712 2150 4764 2202
rect 4776 2150 4828 2202
rect 4840 2150 4892 2202
rect 11982 2150 12034 2202
rect 12046 2150 12098 2202
rect 12110 2150 12162 2202
rect 12174 2150 12226 2202
rect 19315 2150 19367 2202
rect 19379 2150 19431 2202
rect 19443 2150 19495 2202
rect 19507 2150 19559 2202
rect 10048 1980 10100 2032
rect 18144 1980 18196 2032
rect 11152 144 11204 196
rect 12992 76 13044 128
rect 19156 76 19208 128
rect 16948 8 17000 60
<< metal2 >>
rect 846 21570 902 22000
rect 2594 21570 2650 22000
rect 768 21542 902 21570
rect 110 17368 166 17377
rect 110 17303 166 17312
rect 124 17270 152 17303
rect 112 17264 164 17270
rect 112 17206 164 17212
rect 768 17105 796 21542
rect 846 21520 902 21542
rect 2332 21542 2650 21570
rect 1490 20496 1546 20505
rect 1490 20431 1546 20440
rect 1306 18728 1362 18737
rect 1306 18663 1362 18672
rect 754 17096 810 17105
rect 754 17031 810 17040
rect 112 16176 164 16182
rect 112 16118 164 16124
rect 124 15609 152 16118
rect 1320 16114 1348 18663
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 110 15600 166 15609
rect 110 15535 166 15544
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 112 14816 164 14822
rect 112 14758 164 14764
rect 124 11937 152 14758
rect 1308 12640 1360 12646
rect 1308 12582 1360 12588
rect 110 11928 166 11937
rect 110 11863 166 11872
rect 386 9208 442 9217
rect 386 9143 442 9152
rect 110 8528 166 8537
rect 110 8463 166 8472
rect 124 8265 152 8463
rect 110 8256 166 8265
rect 110 8191 166 8200
rect 400 82 428 9143
rect 1320 7750 1348 12582
rect 1412 9178 1440 15438
rect 1504 10266 1532 20431
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1688 13870 1716 14554
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13433 1624 13670
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1596 11354 1624 12242
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1688 11234 1716 13126
rect 1780 12782 1808 13466
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 12442 1808 12718
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1596 11206 1716 11234
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1412 8090 1440 9114
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 1320 7410 1348 7686
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1504 4146 1532 9590
rect 1596 9586 1624 11206
rect 1674 10704 1730 10713
rect 1674 10639 1730 10648
rect 1688 10606 1716 10639
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 1596 8634 1624 9415
rect 1688 9110 1716 10066
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1780 9178 1808 9930
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1676 9104 1728 9110
rect 1676 9046 1728 9052
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 6866 1624 8434
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1688 7206 1716 7958
rect 1780 7546 1808 9114
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6118 1624 6802
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1596 3233 1624 6054
rect 1688 5642 1716 6734
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1688 4826 1716 5578
rect 1872 4826 1900 14894
rect 2056 12782 2084 16662
rect 2332 15162 2360 21542
rect 2594 21520 2650 21542
rect 4434 21570 4490 22000
rect 6274 21570 6330 22000
rect 8114 21570 8170 22000
rect 9954 21570 10010 22000
rect 11794 21570 11850 22000
rect 13634 21570 13690 22000
rect 15474 21570 15530 22000
rect 4434 21542 4568 21570
rect 4434 21520 4490 21542
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 3976 15904 4028 15910
rect 4344 15904 4396 15910
rect 4028 15864 4108 15892
rect 3976 15846 4028 15852
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12374 2084 12718
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11286 1992 11630
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1964 6934 1992 10678
rect 2056 8634 2084 11290
rect 2148 9654 2176 13806
rect 2240 13802 2268 14418
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2608 14006 2636 14214
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2240 11082 2268 13738
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2332 11014 2360 11494
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10606 2360 10950
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2240 10266 2268 10474
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2332 10198 2360 10542
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2148 8838 2176 9454
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 1964 5302 1992 6870
rect 1952 5296 2004 5302
rect 1952 5238 2004 5244
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 3534 1716 4422
rect 1766 4312 1822 4321
rect 1766 4247 1822 4256
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1582 3224 1638 3233
rect 1582 3159 1638 3168
rect 1780 2990 1808 4247
rect 1768 2984 1820 2990
rect 2056 2961 2084 4626
rect 2148 4146 2176 8774
rect 2240 6934 2268 8910
rect 2424 7954 2452 11290
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2228 6928 2280 6934
rect 2228 6870 2280 6876
rect 2240 5778 2268 6870
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5846 2452 6190
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2240 4010 2268 5714
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5273 2360 5510
rect 2318 5264 2374 5273
rect 2318 5199 2374 5208
rect 2332 5166 2360 5199
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2332 4185 2360 4490
rect 2318 4176 2374 4185
rect 2318 4111 2374 4120
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2332 2990 2360 4111
rect 2424 4078 2452 5102
rect 2516 4486 2544 13670
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2424 3602 2452 4014
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2424 3194 2452 3538
rect 2608 3466 2636 13942
rect 2700 10130 2728 14418
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13870 2820 14214
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2792 11218 2820 12174
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10810 2820 11154
rect 2884 11150 2912 15846
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3252 15337 3280 15370
rect 3238 15328 3294 15337
rect 3238 15263 3294 15272
rect 3252 15162 3280 15263
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 2976 13870 3004 14894
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2976 12850 3004 13330
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2976 12306 3004 12786
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2976 11558 3004 12242
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 10804 2832 10810
rect 2832 10764 2912 10792
rect 2780 10746 2832 10752
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 8974 2728 10066
rect 2884 9518 2912 10764
rect 2962 9616 3018 9625
rect 2962 9551 3018 9560
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2792 8498 2820 9386
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2792 8090 2820 8434
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 7970 2912 9454
rect 2976 9042 3004 9551
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8634 3004 8978
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2792 7942 2912 7970
rect 2792 5778 2820 7942
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2976 6730 3004 7210
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6458 3004 6666
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2870 6352 2926 6361
rect 2870 6287 2926 6296
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2792 5370 2820 5714
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2700 4690 2728 4762
rect 2792 4729 2820 5034
rect 2884 4826 2912 6287
rect 3068 5914 3096 14826
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 11898 3188 12650
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3160 11626 3188 11834
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3160 10810 3188 11562
rect 3252 10962 3280 13874
rect 3528 13870 3556 13942
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13394 3464 13738
rect 3528 13530 3556 13806
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12442 3372 13262
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12850 3464 13126
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3436 12374 3464 12786
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11762 3464 12038
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3620 11506 3648 14894
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3436 11478 3648 11506
rect 3252 10934 3372 10962
rect 3148 10804 3200 10810
rect 3200 10764 3280 10792
rect 3148 10746 3200 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10198 3188 10610
rect 3252 10538 3280 10764
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3148 9376 3200 9382
rect 3252 9364 3280 10066
rect 3344 9518 3372 10934
rect 3436 10713 3464 11478
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3528 11014 3556 11290
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3422 10704 3478 10713
rect 3422 10639 3478 10648
rect 3436 10198 3464 10639
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3528 10062 3556 10950
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3200 9336 3280 9364
rect 3148 9318 3200 9324
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2962 5264 3018 5273
rect 2962 5199 3018 5208
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2778 4720 2834 4729
rect 2688 4684 2740 4690
rect 2778 4655 2834 4664
rect 2688 4626 2740 4632
rect 2792 4486 2820 4655
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 3670 2820 4422
rect 2884 4078 2912 4762
rect 2976 4554 3004 5199
rect 3160 4758 3188 9318
rect 3344 9178 3372 9454
rect 3332 9172 3384 9178
rect 3384 9132 3464 9160
rect 3332 9114 3384 9120
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 6390 3280 8774
rect 3344 8362 3372 8842
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3344 8022 3372 8298
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3344 7546 3372 7958
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3344 6934 3372 7210
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3344 6662 3372 6870
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6458 3372 6598
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3436 5030 3464 9132
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2792 3126 2820 3334
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2320 2984 2372 2990
rect 1768 2926 1820 2932
rect 2042 2952 2098 2961
rect 1860 2916 1912 2922
rect 2320 2926 2372 2932
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2042 2887 2098 2896
rect 1860 2858 1912 2864
rect 478 82 534 480
rect 400 54 534 82
rect 478 0 534 54
rect 1490 82 1546 480
rect 1872 82 1900 2858
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2424 2514 2452 2586
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 1964 2417 1992 2450
rect 1950 2408 2006 2417
rect 1950 2343 2006 2352
rect 1964 2310 1992 2343
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1490 54 1900 82
rect 2594 82 2650 480
rect 2700 82 2728 2926
rect 2792 1465 2820 3062
rect 2884 2650 2912 4014
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2976 2514 3004 4490
rect 3436 4298 3464 4626
rect 3160 4270 3464 4298
rect 3160 4214 3188 4270
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3332 4072 3384 4078
rect 3436 4060 3464 4270
rect 3384 4032 3464 4060
rect 3332 4014 3384 4020
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 3068 2650 3096 3402
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3160 2514 3188 3402
rect 3344 3398 3372 4014
rect 3528 3670 3556 9998
rect 3620 5710 3648 11018
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3712 10674 3740 10950
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3712 6746 3740 10134
rect 3804 6934 3832 13466
rect 3896 10742 3924 15574
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3988 12986 4016 13398
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3988 11830 4016 12310
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 4080 11665 4108 15864
rect 4344 15846 4396 15852
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 12986 4200 13262
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 11898 4200 12582
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3988 10470 4016 11222
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10198 4016 10406
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 3896 9110 3924 9959
rect 3988 9722 4016 10134
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3896 8981 3924 9046
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3896 6866 3924 8774
rect 4080 8294 4108 11591
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10810 4200 11086
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4264 10062 4292 15302
rect 4356 13326 4384 15846
rect 4448 15337 4476 18226
rect 4540 17649 4568 21542
rect 6274 21542 6592 21570
rect 6274 21520 6330 21542
rect 4622 19612 4918 19632
rect 4678 19610 4702 19612
rect 4758 19610 4782 19612
rect 4838 19610 4862 19612
rect 4700 19558 4702 19610
rect 4764 19558 4776 19610
rect 4838 19558 4840 19610
rect 4678 19556 4702 19558
rect 4758 19556 4782 19558
rect 4838 19556 4862 19558
rect 4622 19536 4918 19556
rect 6564 18902 6592 21542
rect 7760 21542 8170 21570
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 4622 18524 4918 18544
rect 4678 18522 4702 18524
rect 4758 18522 4782 18524
rect 4838 18522 4862 18524
rect 4700 18470 4702 18522
rect 4764 18470 4776 18522
rect 4838 18470 4840 18522
rect 4678 18468 4702 18470
rect 4758 18468 4782 18470
rect 4838 18468 4862 18470
rect 4622 18448 4918 18468
rect 7760 18426 7788 21542
rect 8114 21520 8170 21542
rect 9784 21542 10010 21570
rect 8289 19068 8585 19088
rect 8345 19066 8369 19068
rect 8425 19066 8449 19068
rect 8505 19066 8529 19068
rect 8367 19014 8369 19066
rect 8431 19014 8443 19066
rect 8505 19014 8507 19066
rect 8345 19012 8369 19014
rect 8425 19012 8449 19014
rect 8505 19012 8529 19014
rect 8289 18992 8585 19012
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 6366 17776 6422 17785
rect 6366 17711 6368 17720
rect 6420 17711 6422 17720
rect 6368 17682 6420 17688
rect 4526 17640 4582 17649
rect 4526 17575 4582 17584
rect 4622 17436 4918 17456
rect 4678 17434 4702 17436
rect 4758 17434 4782 17436
rect 4838 17434 4862 17436
rect 4700 17382 4702 17434
rect 4764 17382 4776 17434
rect 4838 17382 4840 17434
rect 4678 17380 4702 17382
rect 4758 17380 4782 17382
rect 4838 17380 4862 17382
rect 4622 17360 4918 17380
rect 6380 17338 6408 17682
rect 6642 17640 6698 17649
rect 6642 17575 6698 17584
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6368 17332 6420 17338
rect 6420 17292 6500 17320
rect 6368 17274 6420 17280
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 4622 16348 4918 16368
rect 4678 16346 4702 16348
rect 4758 16346 4782 16348
rect 4838 16346 4862 16348
rect 4700 16294 4702 16346
rect 4764 16294 4776 16346
rect 4838 16294 4840 16346
rect 4678 16292 4702 16294
rect 4758 16292 4782 16294
rect 4838 16292 4862 16294
rect 4622 16272 4918 16292
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4434 15328 4490 15337
rect 4434 15263 4490 15272
rect 4540 15094 4568 15982
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4622 15260 4918 15280
rect 4678 15258 4702 15260
rect 4758 15258 4782 15260
rect 4838 15258 4862 15260
rect 4700 15206 4702 15258
rect 4764 15206 4776 15258
rect 4838 15206 4840 15258
rect 4678 15204 4702 15206
rect 4758 15204 4782 15206
rect 4838 15204 4862 15206
rect 4622 15184 4918 15204
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4356 12850 4384 13262
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4264 8634 4292 9046
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3712 6718 3924 6746
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 5137 3648 5170
rect 3712 5166 3740 5850
rect 3804 5846 3832 6598
rect 3896 5914 3924 6718
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3700 5160 3752 5166
rect 3606 5128 3662 5137
rect 3700 5102 3752 5108
rect 3606 5063 3662 5072
rect 3712 4826 3740 5102
rect 3804 5098 3832 5646
rect 4080 5234 4108 8230
rect 4356 7392 4384 11698
rect 4448 9217 4476 14962
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14550 4568 14758
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4540 13734 4568 14486
rect 5000 14482 5028 15438
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4622 14172 4918 14192
rect 4678 14170 4702 14172
rect 4758 14170 4782 14172
rect 4838 14170 4862 14172
rect 4700 14118 4702 14170
rect 4764 14118 4776 14170
rect 4838 14118 4840 14170
rect 4678 14116 4702 14118
rect 4758 14116 4782 14118
rect 4838 14116 4862 14118
rect 4622 14096 4918 14116
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13433 4568 13670
rect 5000 13530 5028 13806
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4526 13424 4582 13433
rect 4526 13359 4582 13368
rect 4622 13084 4918 13104
rect 4678 13082 4702 13084
rect 4758 13082 4782 13084
rect 4838 13082 4862 13084
rect 4700 13030 4702 13082
rect 4764 13030 4776 13082
rect 4838 13030 4840 13082
rect 4678 13028 4702 13030
rect 4758 13028 4782 13030
rect 4838 13028 4862 13030
rect 4622 13008 4918 13028
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4908 12170 4936 12650
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4540 9654 4568 12106
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4622 11996 4918 12016
rect 4678 11994 4702 11996
rect 4758 11994 4782 11996
rect 4838 11994 4862 11996
rect 4700 11942 4702 11994
rect 4764 11942 4776 11994
rect 4838 11942 4840 11994
rect 4678 11940 4702 11942
rect 4758 11940 4782 11942
rect 4838 11940 4862 11942
rect 4622 11920 4918 11940
rect 5000 11898 5028 12038
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5000 11558 5028 11834
rect 5092 11762 5120 15642
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 12986 5212 14758
rect 5276 14521 5304 14894
rect 5368 14890 5396 15506
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5262 14512 5318 14521
rect 5262 14447 5318 14456
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5092 11082 5120 11562
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5184 10962 5212 12038
rect 5092 10934 5212 10962
rect 4622 10908 4918 10928
rect 4678 10906 4702 10908
rect 4758 10906 4782 10908
rect 4838 10906 4862 10908
rect 4700 10854 4702 10906
rect 4764 10854 4776 10906
rect 4838 10854 4840 10906
rect 4678 10852 4702 10854
rect 4758 10852 4782 10854
rect 4838 10852 4862 10854
rect 4622 10832 4918 10852
rect 5092 10198 5120 10934
rect 5276 10588 5304 14350
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 13938 5396 14282
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5460 13814 5488 16390
rect 5552 15910 5580 16594
rect 6472 16572 6500 17292
rect 6380 16544 6500 16572
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5368 13786 5488 13814
rect 5368 13190 5396 13786
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 11762 5396 12786
rect 5460 12442 5488 13670
rect 5552 13462 5580 15846
rect 5736 14618 5764 15982
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5184 10560 5304 10588
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 4622 9820 4918 9840
rect 4678 9818 4702 9820
rect 4758 9818 4782 9820
rect 4838 9818 4862 9820
rect 4700 9766 4702 9818
rect 4764 9766 4776 9818
rect 4838 9766 4840 9818
rect 4678 9764 4702 9766
rect 4758 9764 4782 9766
rect 4838 9764 4862 9766
rect 4622 9744 4918 9764
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4434 9208 4490 9217
rect 4434 9143 4490 9152
rect 4540 7954 4568 9386
rect 5092 9178 5120 9522
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4622 8732 4918 8752
rect 4678 8730 4702 8732
rect 4758 8730 4782 8732
rect 4838 8730 4862 8732
rect 4700 8678 4702 8730
rect 4764 8678 4776 8730
rect 4838 8678 4840 8730
rect 4678 8676 4702 8678
rect 4758 8676 4782 8678
rect 4838 8676 4862 8678
rect 4622 8656 4918 8676
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4724 8090 4752 8298
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8090 5120 8230
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4540 7546 4568 7890
rect 4622 7644 4918 7664
rect 4678 7642 4702 7644
rect 4758 7642 4782 7644
rect 4838 7642 4862 7644
rect 4700 7590 4702 7642
rect 4764 7590 4776 7642
rect 4838 7590 4840 7642
rect 4678 7588 4702 7590
rect 4758 7588 4782 7590
rect 4838 7588 4862 7590
rect 4622 7568 4918 7588
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4356 7364 4476 7392
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4172 6322 4200 6802
rect 4250 6760 4306 6769
rect 4250 6695 4306 6704
rect 4264 6662 4292 6695
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4172 6118 4200 6258
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3712 4078 3740 4762
rect 3804 4690 3832 5034
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 4282 3832 4626
rect 3988 4622 4016 4762
rect 4264 4758 4292 5714
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 4616 4028 4622
rect 4080 4593 4108 4626
rect 3976 4558 4028 4564
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 4080 4214 4108 4519
rect 4264 4321 4292 4694
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4250 4312 4306 4321
rect 4250 4247 4306 4256
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3528 2990 3556 3062
rect 3620 2990 3648 3946
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3792 3596 3844 3602
rect 3896 3584 3924 3878
rect 4080 3602 4108 4150
rect 4356 4146 4384 4626
rect 4448 4214 4476 7364
rect 5092 7206 5120 8026
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6934 5120 7142
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4622 6556 4918 6576
rect 4678 6554 4702 6556
rect 4758 6554 4782 6556
rect 4838 6554 4862 6556
rect 4700 6502 4702 6554
rect 4764 6502 4776 6554
rect 4838 6502 4840 6554
rect 4678 6500 4702 6502
rect 4758 6500 4782 6502
rect 4838 6500 4862 6502
rect 4622 6480 4918 6500
rect 5000 6322 5028 6598
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5000 5846 5028 6258
rect 5092 6186 5120 6870
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4540 5370 4568 5714
rect 4622 5468 4918 5488
rect 4678 5466 4702 5468
rect 4758 5466 4782 5468
rect 4838 5466 4862 5468
rect 4700 5414 4702 5466
rect 4764 5414 4776 5466
rect 4838 5414 4840 5466
rect 4678 5412 4702 5414
rect 4758 5412 4782 5414
rect 4838 5412 4862 5414
rect 4622 5392 4918 5412
rect 5092 5370 5120 6122
rect 5184 5914 5212 10560
rect 5356 10532 5408 10538
rect 5276 10492 5356 10520
rect 5276 9926 5304 10492
rect 5356 10474 5408 10480
rect 5460 10033 5488 10950
rect 5540 10056 5592 10062
rect 5446 10024 5502 10033
rect 5540 9998 5592 10004
rect 5446 9959 5502 9968
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 9722 5304 9862
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5356 9648 5408 9654
rect 5262 9616 5318 9625
rect 5356 9590 5408 9596
rect 5262 9551 5318 9560
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4250 4040 4306 4049
rect 4250 3975 4306 3984
rect 3844 3556 3924 3584
rect 3792 3538 3844 3544
rect 3896 3126 3924 3556
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3528 2310 3556 2926
rect 4264 2650 4292 3975
rect 4356 3942 4384 4082
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4448 3058 4476 4150
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 2594 54 2728 82
rect 3528 82 3556 2246
rect 3698 82 3754 480
rect 3528 54 3754 82
rect 4540 82 4568 5170
rect 5092 5098 5120 5306
rect 5184 5234 5212 5850
rect 5276 5681 5304 9551
rect 5368 7834 5396 9590
rect 5460 9110 5488 9959
rect 5552 9178 5580 9998
rect 5644 9586 5672 13466
rect 5736 13394 5764 13942
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5736 12850 5764 13330
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5736 10266 5764 11086
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8498 5488 9046
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8537 5672 8978
rect 5630 8528 5686 8537
rect 5448 8492 5500 8498
rect 5630 8463 5686 8472
rect 5448 8434 5500 8440
rect 5644 8430 5672 8463
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5368 7806 5488 7834
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7274 5396 7686
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5460 5914 5488 7806
rect 5828 6882 5856 12922
rect 5920 10742 5948 16118
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13394 6132 13670
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6104 13190 6132 13330
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5920 9994 5948 10678
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 6012 8922 6040 13126
rect 6104 12646 6132 13126
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6104 11830 6132 12378
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6104 11558 6132 11766
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11286 6132 11494
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6104 10606 6132 11222
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5736 6854 5856 6882
rect 5920 8894 6040 8922
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5262 5672 5318 5681
rect 5262 5607 5318 5616
rect 5262 5264 5318 5273
rect 5172 5228 5224 5234
rect 5262 5199 5318 5208
rect 5172 5170 5224 5176
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 5092 4826 5120 4927
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4622 4380 4918 4400
rect 4678 4378 4702 4380
rect 4758 4378 4782 4380
rect 4838 4378 4862 4380
rect 4700 4326 4702 4378
rect 4764 4326 4776 4378
rect 4838 4326 4840 4378
rect 4678 4324 4702 4326
rect 4758 4324 4782 4326
rect 4838 4324 4862 4326
rect 4622 4304 4918 4324
rect 5276 4214 5304 5199
rect 5644 4826 5672 6122
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5460 4486 5488 4762
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4480 5500 4486
rect 5354 4448 5410 4457
rect 5448 4422 5500 4428
rect 5354 4383 5410 4392
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3738 5212 3946
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 4622 3292 4918 3312
rect 4678 3290 4702 3292
rect 4758 3290 4782 3292
rect 4838 3290 4862 3292
rect 4700 3238 4702 3290
rect 4764 3238 4776 3290
rect 4838 3238 4840 3290
rect 4678 3236 4702 3238
rect 4758 3236 4782 3238
rect 4838 3236 4862 3238
rect 4622 3216 4918 3236
rect 5276 2650 5304 4150
rect 5368 3602 5396 4383
rect 5460 4078 5488 4422
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5552 3738 5580 4694
rect 5736 4690 5764 6854
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 5710 5856 6734
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5920 5216 5948 8894
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6012 8294 6040 8774
rect 6104 8566 6132 9862
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7410 6040 8230
rect 6104 7478 6132 8502
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6104 6866 6132 7414
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6196 6730 6224 16050
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6288 10470 6316 12582
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6380 10146 6408 16544
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6472 15026 6500 15506
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6472 13394 6500 14350
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6472 11354 6500 13194
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6288 10118 6408 10146
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6288 8634 6316 10118
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 8838 6408 9998
rect 6472 9654 6500 10134
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6288 8090 6316 8570
rect 6380 8566 6408 8774
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7206 6316 7822
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5574 6040 6054
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6000 5228 6052 5234
rect 5920 5188 6000 5216
rect 6000 5170 6052 5176
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 6104 4154 6132 5646
rect 6012 4126 6132 4154
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5644 3738 5672 4014
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 3194 5396 3538
rect 5460 3194 5488 3606
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5460 2582 5488 2790
rect 5448 2576 5500 2582
rect 4618 2544 4674 2553
rect 5448 2518 5500 2524
rect 4618 2479 4674 2488
rect 4632 2446 4660 2479
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4622 2204 4918 2224
rect 4678 2202 4702 2204
rect 4758 2202 4782 2204
rect 4838 2202 4862 2204
rect 4700 2150 4702 2202
rect 4764 2150 4776 2202
rect 4838 2150 4840 2202
rect 4678 2148 4702 2150
rect 4758 2148 4782 2150
rect 4838 2148 4862 2150
rect 4622 2128 4918 2148
rect 4802 82 4858 480
rect 4540 54 4858 82
rect 1490 0 1546 54
rect 2594 0 2650 54
rect 3698 0 3754 54
rect 4802 0 4858 54
rect 5906 82 5962 480
rect 6012 82 6040 4126
rect 6196 3670 6224 5850
rect 6288 4146 6316 7142
rect 6380 6798 6408 7686
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6564 5914 6592 17478
rect 6656 16658 6684 17575
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6656 16250 6684 16594
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6644 16040 6696 16046
rect 6642 16008 6644 16017
rect 6696 16008 6698 16017
rect 6642 15943 6698 15952
rect 6656 15910 6684 15943
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6656 12918 6684 14554
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6748 12850 6776 16390
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6656 12442 6684 12582
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6656 11898 6684 12378
rect 6748 12306 6776 12786
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6656 11558 6684 11834
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6840 11354 6868 15914
rect 6932 11762 6960 16390
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6656 11014 6684 11222
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10538 6684 10746
rect 6840 10742 6868 11290
rect 6932 11218 6960 11698
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6736 10600 6788 10606
rect 6788 10560 6960 10588
rect 6736 10542 6788 10548
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6734 9616 6790 9625
rect 6734 9551 6790 9560
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 8634 6684 8978
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6656 6458 6684 6870
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6748 5710 6776 9551
rect 6840 6186 6868 10406
rect 6932 9450 6960 10560
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7024 8956 7052 14758
rect 7116 13002 7144 15370
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7208 14414 7236 14894
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7116 12974 7236 13002
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7116 9110 7144 12854
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7208 8956 7236 12974
rect 7300 11132 7328 16934
rect 7392 11234 7420 18294
rect 8220 18086 8248 18770
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7484 13938 7512 14486
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7576 11744 7604 17478
rect 7760 17066 7788 17682
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7760 16969 7788 17002
rect 7746 16960 7802 16969
rect 7746 16895 7802 16904
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7944 16182 7972 16390
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7944 15638 7972 16118
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7668 13870 7696 14010
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7668 13258 7696 13806
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7576 11716 7696 11744
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7392 11206 7512 11234
rect 7380 11144 7432 11150
rect 7300 11104 7380 11132
rect 7380 11086 7432 11092
rect 7392 10742 7420 11086
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 10266 7328 10610
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7024 8928 7144 8956
rect 7208 8928 7420 8956
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6932 7410 6960 8842
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7024 7274 7052 7686
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6932 7002 6960 7210
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7024 6390 7052 6734
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6564 4826 6592 5238
rect 6748 5166 6776 5646
rect 6840 5302 6868 5782
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6932 5234 6960 5646
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6472 3942 6500 4694
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6288 2922 6316 3606
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6380 2650 6408 3674
rect 6472 2990 6500 3878
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6472 2650 6500 2926
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6932 2514 6960 3470
rect 7024 2582 7052 3878
rect 7116 3534 7144 8928
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 6798 7328 7346
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 6322 7236 6666
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7300 5234 7328 5578
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4826 7236 4966
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7208 4214 7236 4762
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7300 4154 7328 5170
rect 7392 4604 7420 8928
rect 7484 8498 7512 11206
rect 7576 10674 7604 11562
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 9110 7604 9386
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 7750 7512 8230
rect 7576 8022 7604 8298
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6186 7512 7686
rect 7576 7274 7604 7958
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7668 7002 7696 11716
rect 7760 10266 7788 13738
rect 7852 13569 7880 15098
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14618 7972 14894
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7944 14521 7972 14554
rect 7930 14512 7986 14521
rect 7930 14447 7986 14456
rect 7838 13560 7894 13569
rect 8036 13512 8064 17070
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 7838 13495 7894 13504
rect 7944 13484 8064 13512
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7852 11150 7880 12650
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7944 10996 7972 13484
rect 8022 13424 8078 13433
rect 8022 13359 8078 13368
rect 8036 13326 8064 13359
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12306 8064 13262
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11898 8064 12242
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8128 11642 8156 15846
rect 8220 15688 8248 18022
rect 8289 17980 8585 18000
rect 8345 17978 8369 17980
rect 8425 17978 8449 17980
rect 8505 17978 8529 17980
rect 8367 17926 8369 17978
rect 8431 17926 8443 17978
rect 8505 17926 8507 17978
rect 8345 17924 8369 17926
rect 8425 17924 8449 17926
rect 8505 17924 8529 17926
rect 8289 17904 8585 17924
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8680 17338 8708 17682
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8772 16969 8800 18090
rect 8758 16960 8814 16969
rect 8289 16892 8585 16912
rect 8758 16895 8814 16904
rect 8345 16890 8369 16892
rect 8425 16890 8449 16892
rect 8505 16890 8529 16892
rect 8367 16838 8369 16890
rect 8431 16838 8443 16890
rect 8505 16838 8507 16890
rect 8345 16836 8369 16838
rect 8425 16836 8449 16838
rect 8505 16836 8529 16838
rect 8289 16816 8585 16836
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8772 16114 8800 16594
rect 8864 16289 8892 18566
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9416 17814 9444 18022
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8850 16280 8906 16289
rect 8850 16215 8906 16224
rect 9048 16182 9076 16390
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8289 15804 8585 15824
rect 8345 15802 8369 15804
rect 8425 15802 8449 15804
rect 8505 15802 8529 15804
rect 8367 15750 8369 15802
rect 8431 15750 8443 15802
rect 8505 15750 8507 15802
rect 8345 15748 8369 15750
rect 8425 15748 8449 15750
rect 8505 15748 8529 15750
rect 8289 15728 8585 15748
rect 8680 15722 8708 15914
rect 8772 15892 8800 16050
rect 8852 15904 8904 15910
rect 8772 15864 8852 15892
rect 8852 15846 8904 15852
rect 8680 15694 8800 15722
rect 8220 15660 8340 15688
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8220 15162 8248 15506
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8312 15042 8340 15660
rect 8036 11614 8156 11642
rect 8220 15014 8340 15042
rect 8036 11150 8064 11614
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7852 10968 7972 10996
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 9518 7788 10202
rect 7748 9512 7800 9518
rect 7852 9489 7880 10968
rect 8128 10810 8156 11494
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9926 7972 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7748 9454 7800 9460
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7852 8974 7880 9415
rect 7944 9042 7972 9862
rect 8036 9586 8064 10134
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9178 8064 9522
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7944 6390 7972 8978
rect 8220 6916 8248 15014
rect 8289 14716 8585 14736
rect 8345 14714 8369 14716
rect 8425 14714 8449 14716
rect 8505 14714 8529 14716
rect 8367 14662 8369 14714
rect 8431 14662 8443 14714
rect 8505 14662 8507 14714
rect 8345 14660 8369 14662
rect 8425 14660 8449 14662
rect 8505 14660 8529 14662
rect 8289 14640 8585 14660
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8312 14074 8340 14418
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8680 14006 8708 14282
rect 8772 14006 8800 15694
rect 8864 15473 8892 15846
rect 9048 15502 9076 16118
rect 9036 15496 9088 15502
rect 8850 15464 8906 15473
rect 9036 15438 9088 15444
rect 8850 15399 8906 15408
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8864 14346 8892 14894
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8289 13628 8585 13648
rect 8345 13626 8369 13628
rect 8425 13626 8449 13628
rect 8505 13626 8529 13628
rect 8367 13574 8369 13626
rect 8431 13574 8443 13626
rect 8505 13574 8507 13626
rect 8345 13572 8369 13574
rect 8425 13572 8449 13574
rect 8505 13572 8529 13574
rect 8289 13552 8585 13572
rect 8680 13394 8708 13942
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 13462 8800 13806
rect 8864 13734 8892 13874
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8312 12986 8340 13330
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 12850 8340 12922
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8680 12646 8708 13330
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8289 12540 8585 12560
rect 8345 12538 8369 12540
rect 8425 12538 8449 12540
rect 8505 12538 8529 12540
rect 8367 12486 8369 12538
rect 8431 12486 8443 12538
rect 8505 12486 8507 12538
rect 8345 12484 8369 12486
rect 8425 12484 8449 12486
rect 8505 12484 8529 12486
rect 8289 12464 8585 12484
rect 8576 12300 8628 12306
rect 8680 12288 8708 12582
rect 8628 12260 8708 12288
rect 8576 12242 8628 12248
rect 8588 11694 8616 12242
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8289 11452 8585 11472
rect 8345 11450 8369 11452
rect 8425 11450 8449 11452
rect 8505 11450 8529 11452
rect 8367 11398 8369 11450
rect 8431 11398 8443 11450
rect 8505 11398 8507 11450
rect 8345 11396 8369 11398
rect 8425 11396 8449 11398
rect 8505 11396 8529 11398
rect 8289 11376 8585 11396
rect 8289 10364 8585 10384
rect 8345 10362 8369 10364
rect 8425 10362 8449 10364
rect 8505 10362 8529 10364
rect 8367 10310 8369 10362
rect 8431 10310 8443 10362
rect 8505 10310 8507 10362
rect 8345 10308 8369 10310
rect 8425 10308 8449 10310
rect 8505 10308 8529 10310
rect 8289 10288 8585 10308
rect 8289 9276 8585 9296
rect 8345 9274 8369 9276
rect 8425 9274 8449 9276
rect 8505 9274 8529 9276
rect 8367 9222 8369 9274
rect 8431 9222 8443 9274
rect 8505 9222 8507 9274
rect 8345 9220 8369 9222
rect 8425 9220 8449 9222
rect 8505 9220 8529 9222
rect 8289 9200 8585 9220
rect 8289 8188 8585 8208
rect 8345 8186 8369 8188
rect 8425 8186 8449 8188
rect 8505 8186 8529 8188
rect 8367 8134 8369 8186
rect 8431 8134 8443 8186
rect 8505 8134 8507 8186
rect 8345 8132 8369 8134
rect 8425 8132 8449 8134
rect 8505 8132 8529 8134
rect 8289 8112 8585 8132
rect 8666 7984 8722 7993
rect 8666 7919 8722 7928
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 7342 8616 7686
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8289 7100 8585 7120
rect 8345 7098 8369 7100
rect 8425 7098 8449 7100
rect 8505 7098 8529 7100
rect 8367 7046 8369 7098
rect 8431 7046 8443 7098
rect 8505 7046 8507 7098
rect 8345 7044 8369 7046
rect 8425 7044 8449 7046
rect 8505 7044 8529 7046
rect 8289 7024 8585 7044
rect 8128 6888 8248 6916
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7576 4758 7604 4966
rect 7668 4826 7696 5510
rect 7760 5166 7788 5714
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7392 4576 7604 4604
rect 7300 4126 7420 4154
rect 7392 3602 7420 4126
rect 7576 3738 7604 4576
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7668 4146 7696 4490
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7194 3496 7250 3505
rect 7194 3431 7250 3440
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 5906 54 6040 82
rect 7010 82 7066 480
rect 7208 82 7236 3431
rect 7392 3058 7420 3538
rect 7760 3466 7788 5102
rect 7852 5001 7880 5170
rect 7838 4992 7894 5001
rect 7838 4927 7894 4936
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 7852 3942 7880 4694
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7484 2922 7512 3334
rect 7852 2922 7880 3606
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7484 2650 7512 2858
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7748 2576 7800 2582
rect 7852 2564 7880 2858
rect 7944 2650 7972 4762
rect 8128 4049 8156 6888
rect 8680 6866 8708 7919
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8680 6458 8708 6802
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8289 6012 8585 6032
rect 8345 6010 8369 6012
rect 8425 6010 8449 6012
rect 8505 6010 8529 6012
rect 8367 5958 8369 6010
rect 8431 5958 8443 6010
rect 8505 5958 8507 6010
rect 8345 5956 8369 5958
rect 8425 5956 8449 5958
rect 8505 5956 8529 5958
rect 8289 5936 8585 5956
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8220 5817 8248 5850
rect 8206 5808 8262 5817
rect 8206 5743 8262 5752
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8220 4758 8248 5238
rect 8312 5234 8340 5714
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8289 4924 8585 4944
rect 8345 4922 8369 4924
rect 8425 4922 8449 4924
rect 8505 4922 8529 4924
rect 8367 4870 8369 4922
rect 8431 4870 8443 4922
rect 8505 4870 8507 4922
rect 8345 4868 8369 4870
rect 8425 4868 8449 4870
rect 8505 4868 8529 4870
rect 8289 4848 8585 4868
rect 8680 4826 8708 5034
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8208 4752 8260 4758
rect 8772 4729 8800 12922
rect 8864 12646 8892 13670
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 10470 8892 12582
rect 8956 10674 8984 14962
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9450 8892 10406
rect 8956 10266 8984 10610
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9048 9722 9076 14758
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 9140 8498 9168 17478
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9404 17196 9456 17202
rect 9324 17156 9404 17184
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 12866 9260 16934
rect 9324 16833 9352 17156
rect 9404 17138 9456 17144
rect 9310 16824 9366 16833
rect 9310 16759 9366 16768
rect 9324 16250 9352 16759
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9324 15366 9352 16050
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9312 15360 9364 15366
rect 9402 15328 9458 15337
rect 9364 15308 9402 15314
rect 9312 15302 9402 15308
rect 9324 15286 9402 15302
rect 9402 15263 9458 15272
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9324 14550 9352 14962
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9324 13326 9352 14350
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9416 12986 9444 15098
rect 9508 15026 9536 15914
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9496 14544 9548 14550
rect 9600 14521 9628 17274
rect 9496 14486 9548 14492
rect 9586 14512 9642 14521
rect 9508 13734 9536 14486
rect 9586 14447 9642 14456
rect 9692 14396 9720 17614
rect 9784 16794 9812 21542
rect 9954 21520 10010 21542
rect 11532 21542 11850 21570
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10704 18970 10732 19110
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10520 17338 10548 18838
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10704 18426 10732 18770
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10692 18420 10744 18426
rect 10612 18380 10692 18408
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10520 17134 10548 17274
rect 10612 17202 10640 18380
rect 10692 18362 10744 18368
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9784 15162 9812 15506
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9968 14414 9996 17070
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9772 14408 9824 14414
rect 9692 14368 9772 14396
rect 9956 14408 10008 14414
rect 9772 14350 9824 14356
rect 9862 14376 9918 14385
rect 9784 14074 9812 14350
rect 9956 14350 10008 14356
rect 9862 14311 9918 14320
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9876 14006 9904 14311
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9508 13530 9536 13670
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9232 12838 9444 12866
rect 9508 12850 9536 13194
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12374 9260 12718
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9218 12200 9274 12209
rect 9218 12135 9274 12144
rect 9232 11218 9260 12135
rect 9324 11898 9352 12310
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 6866 8892 8026
rect 9048 7206 9076 8230
rect 9140 8090 9168 8434
rect 9324 8090 9352 11630
rect 9416 10198 9444 12838
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8864 6458 8892 6802
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8956 6322 8984 6938
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9048 6186 9076 7142
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8864 5710 8892 5850
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5098 8892 5646
rect 8956 5370 8984 6054
rect 9048 5914 9076 6122
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9140 5778 9168 7822
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8956 4758 8984 5306
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8944 4752 8996 4758
rect 8208 4694 8260 4700
rect 8758 4720 8814 4729
rect 8944 4694 8996 4700
rect 8758 4655 8814 4664
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8114 4040 8170 4049
rect 8036 3998 8114 4026
rect 8036 3058 8064 3998
rect 8114 3975 8170 3984
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8128 2582 8156 3470
rect 7800 2536 7880 2564
rect 8116 2576 8168 2582
rect 7748 2518 7800 2524
rect 8116 2518 8168 2524
rect 7010 54 7236 82
rect 8114 82 8170 480
rect 8220 82 8248 4218
rect 8574 4040 8630 4049
rect 8668 4004 8720 4010
rect 8630 3984 8668 3992
rect 8574 3975 8668 3984
rect 8588 3964 8668 3975
rect 8668 3946 8720 3952
rect 8772 3942 8800 4422
rect 8956 4282 8984 4694
rect 9140 4468 9168 5170
rect 9220 4480 9272 4486
rect 9140 4440 9220 4468
rect 9220 4422 9272 4428
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8289 3836 8585 3856
rect 8345 3834 8369 3836
rect 8425 3834 8449 3836
rect 8505 3834 8529 3836
rect 8367 3782 8369 3834
rect 8431 3782 8443 3834
rect 8505 3782 8507 3834
rect 8345 3780 8369 3782
rect 8425 3780 8449 3782
rect 8505 3780 8529 3782
rect 8289 3760 8585 3780
rect 8772 3738 8800 3878
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 9126 2952 9182 2961
rect 9126 2887 9182 2896
rect 8289 2748 8585 2768
rect 8345 2746 8369 2748
rect 8425 2746 8449 2748
rect 8505 2746 8529 2748
rect 8367 2694 8369 2746
rect 8431 2694 8443 2746
rect 8505 2694 8507 2746
rect 8345 2692 8369 2694
rect 8425 2692 8449 2694
rect 8505 2692 8529 2694
rect 8289 2672 8585 2692
rect 9140 2514 9168 2887
rect 9232 2650 9260 4422
rect 9324 3738 9352 5850
rect 9508 5778 9536 12786
rect 9600 7886 9628 13942
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12918 9720 13262
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5302 9444 5510
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9692 4554 9720 10406
rect 9784 8294 9812 13874
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 12646 9996 13398
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 10060 11762 10088 16934
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10152 16046 10180 16594
rect 10232 16584 10284 16590
rect 10520 16561 10548 17070
rect 10232 16526 10284 16532
rect 10506 16552 10562 16561
rect 10244 16114 10272 16526
rect 10506 16487 10562 16496
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9876 10810 9904 11562
rect 10060 11354 10088 11698
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10060 10470 10088 11154
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9864 10192 9916 10198
rect 10152 10146 10180 15982
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 14006 10364 15846
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10428 13852 10456 14758
rect 10520 14550 10548 14894
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 14006 10548 14350
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 9864 10134 9916 10140
rect 9876 9110 9904 10134
rect 10060 10118 10180 10146
rect 10336 13824 10456 13852
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9968 9178 9996 9658
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9862 8936 9918 8945
rect 9862 8871 9918 8880
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7206 9812 7890
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6186 9812 7142
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9784 5370 9812 5714
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 4321 9812 4422
rect 9770 4312 9826 4321
rect 9770 4247 9826 4256
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9680 4004 9732 4010
rect 9784 3992 9812 4150
rect 9732 3964 9812 3992
rect 9680 3946 9732 3952
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9324 3058 9352 3674
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 8114 54 8248 82
rect 9218 82 9274 480
rect 9508 82 9536 3878
rect 9876 2514 9904 8871
rect 10060 7546 10088 10118
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 8498 10180 9998
rect 10336 9674 10364 13824
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10244 9646 10364 9674
rect 10244 9382 10272 9646
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 8634 10272 9318
rect 10428 8634 10456 12378
rect 10520 12306 10548 13942
rect 10612 13326 10640 16186
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12374 10640 13126
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11626 10548 12106
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10612 11665 10640 11698
rect 10598 11656 10654 11665
rect 10508 11620 10560 11626
rect 10598 11591 10654 11600
rect 10508 11562 10560 11568
rect 10520 11286 10548 11562
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 9450 10548 10406
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 7540 10100 7546
rect 9968 7500 10048 7528
rect 9968 4690 9996 7500
rect 10048 7482 10100 7488
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9968 4282 9996 4626
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 10060 2038 10088 6598
rect 10152 4486 10180 8230
rect 10244 8090 10272 8570
rect 10428 8362 10456 8570
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10520 7274 10548 9386
rect 10612 8974 10640 10950
rect 10704 9466 10732 18090
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10796 16969 10824 17002
rect 10782 16960 10838 16969
rect 10782 16895 10838 16904
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10796 15706 10824 15982
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10796 15094 10824 15642
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10796 14482 10824 14894
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13938 10824 14214
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13814 10916 18566
rect 10796 13786 10916 13814
rect 10796 11286 10824 13786
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13190 10916 13670
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12986 10916 13126
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10674 10824 11086
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10888 10538 10916 10746
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10704 9438 10824 9466
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9110 10732 9318
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8498 10640 8910
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6254 10640 6598
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10520 4282 10548 5306
rect 10612 4593 10640 6190
rect 10704 5370 10732 6734
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10598 4584 10654 4593
rect 10796 4554 10824 9438
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10888 6186 10916 6802
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5914 10916 6122
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10874 5672 10930 5681
rect 10874 5607 10930 5616
rect 10598 4519 10654 4528
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10888 4078 10916 5607
rect 10980 5234 11008 19110
rect 11072 10062 11100 19382
rect 11532 18834 11560 21542
rect 11794 21520 11850 21542
rect 13372 21542 13690 21570
rect 11956 19612 12252 19632
rect 12012 19610 12036 19612
rect 12092 19610 12116 19612
rect 12172 19610 12196 19612
rect 12034 19558 12036 19610
rect 12098 19558 12110 19610
rect 12172 19558 12174 19610
rect 12012 19556 12036 19558
rect 12092 19556 12116 19558
rect 12172 19556 12196 19558
rect 11956 19536 12252 19556
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11164 11694 11192 18158
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11348 15638 11376 17206
rect 11428 15972 11480 15978
rect 11428 15914 11480 15920
rect 11440 15881 11468 15914
rect 11426 15872 11482 15881
rect 11426 15807 11482 15816
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 12442 11284 15438
rect 11348 14958 11376 15574
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11348 14793 11376 14894
rect 11440 14822 11468 15506
rect 11428 14816 11480 14822
rect 11334 14784 11390 14793
rect 11428 14758 11480 14764
rect 11334 14719 11390 14728
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 11898 11284 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11164 10470 11192 11290
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11072 9654 11100 9998
rect 11164 9722 11192 10134
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 11164 9518 11192 9551
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11164 8498 11192 8842
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7002 11100 7686
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 4826 11008 5034
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11072 4154 11100 6666
rect 11164 6390 11192 7346
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11256 6168 11284 11222
rect 11348 11218 11376 14554
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11440 13938 11468 14418
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11440 13530 11468 13874
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12918 11468 13262
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10266 11376 11154
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11164 6140 11284 6168
rect 11164 4622 11192 6140
rect 11440 5914 11468 12854
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11348 5370 11376 5714
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11256 4214 11284 4694
rect 11244 4208 11296 4214
rect 11072 4126 11192 4154
rect 11244 4150 11296 4156
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3738 10180 3946
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10152 3194 10180 3674
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 3466 10824 3538
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 9218 54 9536 82
rect 10322 82 10378 480
rect 10428 82 10456 3334
rect 10704 3126 10732 3334
rect 10796 3194 10824 3402
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10704 2650 10732 2858
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10322 54 10456 82
rect 10888 82 10916 4014
rect 11164 202 11192 4126
rect 11256 3720 11284 4150
rect 11336 3732 11388 3738
rect 11256 3692 11336 3720
rect 11336 3674 11388 3680
rect 11440 2990 11468 5714
rect 11532 4154 11560 18566
rect 11624 18222 11652 19110
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11808 18426 11836 18770
rect 11956 18524 12252 18544
rect 12012 18522 12036 18524
rect 12092 18522 12116 18524
rect 12172 18522 12196 18524
rect 12034 18470 12036 18522
rect 12098 18470 12110 18522
rect 12172 18470 12174 18522
rect 12012 18468 12036 18470
rect 12092 18468 12116 18470
rect 12172 18468 12196 18470
rect 11956 18448 12252 18468
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17270 11744 17682
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11716 17105 11744 17206
rect 11702 17096 11758 17105
rect 11702 17031 11758 17040
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11624 12918 11652 15914
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 11762 11652 12582
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 9178 11652 11494
rect 11716 11150 11744 16934
rect 11808 14550 11836 17478
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11716 6882 11744 10950
rect 11808 8838 11836 14350
rect 11900 10674 11928 18090
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 11956 17436 12252 17456
rect 12012 17434 12036 17436
rect 12092 17434 12116 17436
rect 12172 17434 12196 17436
rect 12034 17382 12036 17434
rect 12098 17382 12110 17434
rect 12172 17382 12174 17434
rect 12012 17380 12036 17382
rect 12092 17380 12116 17382
rect 12172 17380 12196 17382
rect 11956 17360 12252 17380
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 11956 16348 12252 16368
rect 12012 16346 12036 16348
rect 12092 16346 12116 16348
rect 12172 16346 12196 16348
rect 12034 16294 12036 16346
rect 12098 16294 12110 16346
rect 12172 16294 12174 16346
rect 12012 16292 12036 16294
rect 12092 16292 12116 16294
rect 12172 16292 12196 16294
rect 11956 16272 12252 16292
rect 11956 15260 12252 15280
rect 12012 15258 12036 15260
rect 12092 15258 12116 15260
rect 12172 15258 12196 15260
rect 12034 15206 12036 15258
rect 12098 15206 12110 15258
rect 12172 15206 12174 15258
rect 12012 15204 12036 15206
rect 12092 15204 12116 15206
rect 12172 15204 12196 15206
rect 11956 15184 12252 15204
rect 12360 15178 12388 16730
rect 12452 15960 12480 18022
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17134 12572 17478
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12452 15932 12572 15960
rect 12360 15150 12480 15178
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 11956 14172 12252 14192
rect 12012 14170 12036 14172
rect 12092 14170 12116 14172
rect 12172 14170 12196 14172
rect 12034 14118 12036 14170
rect 12098 14118 12110 14170
rect 12172 14118 12174 14170
rect 12012 14116 12036 14118
rect 12092 14116 12116 14118
rect 12172 14116 12196 14118
rect 11956 14096 12252 14116
rect 12070 13968 12126 13977
rect 12070 13903 12126 13912
rect 12084 13734 12112 13903
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13258 12112 13670
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11956 13084 12252 13104
rect 12012 13082 12036 13084
rect 12092 13082 12116 13084
rect 12172 13082 12196 13084
rect 12034 13030 12036 13082
rect 12098 13030 12110 13082
rect 12172 13030 12174 13082
rect 12012 13028 12036 13030
rect 12092 13028 12116 13030
rect 12172 13028 12196 13030
rect 11956 13008 12252 13028
rect 12360 12850 12388 14486
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12306 12204 12582
rect 12360 12442 12388 12786
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 11956 11996 12252 12016
rect 12012 11994 12036 11996
rect 12092 11994 12116 11996
rect 12172 11994 12196 11996
rect 12034 11942 12036 11994
rect 12098 11942 12110 11994
rect 12172 11942 12174 11994
rect 12012 11940 12036 11942
rect 12092 11940 12116 11942
rect 12172 11940 12196 11942
rect 11956 11920 12252 11940
rect 12164 11552 12216 11558
rect 12360 11540 12388 12242
rect 12216 11512 12388 11540
rect 12164 11494 12216 11500
rect 12176 11354 12204 11494
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 11014 12388 11222
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 11956 10908 12252 10928
rect 12012 10906 12036 10908
rect 12092 10906 12116 10908
rect 12172 10906 12196 10908
rect 12034 10854 12036 10906
rect 12098 10854 12110 10906
rect 12172 10854 12174 10906
rect 12012 10852 12036 10854
rect 12092 10852 12116 10854
rect 12172 10852 12196 10854
rect 11956 10832 12252 10852
rect 12360 10810 12388 10950
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 12360 10470 12388 10746
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 11956 9820 12252 9840
rect 12012 9818 12036 9820
rect 12092 9818 12116 9820
rect 12172 9818 12196 9820
rect 12034 9766 12036 9818
rect 12098 9766 12110 9818
rect 12172 9766 12174 9818
rect 12012 9764 12036 9766
rect 12092 9764 12116 9766
rect 12172 9764 12196 9766
rect 11956 9744 12252 9764
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11900 8294 11928 9046
rect 11956 8732 12252 8752
rect 12012 8730 12036 8732
rect 12092 8730 12116 8732
rect 12172 8730 12196 8732
rect 12034 8678 12036 8730
rect 12098 8678 12110 8730
rect 12172 8678 12174 8730
rect 12012 8676 12036 8678
rect 12092 8676 12116 8678
rect 12172 8676 12196 8678
rect 11956 8656 12252 8676
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11808 7188 11836 7958
rect 11900 7478 11928 8230
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 11956 7644 12252 7664
rect 12012 7642 12036 7644
rect 12092 7642 12116 7644
rect 12172 7642 12196 7644
rect 12034 7590 12036 7642
rect 12098 7590 12110 7642
rect 12172 7590 12174 7642
rect 12012 7588 12036 7590
rect 12092 7588 12116 7590
rect 12172 7588 12196 7590
rect 11956 7568 12252 7588
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 12360 7410 12388 7686
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 11888 7200 11940 7206
rect 11808 7160 11888 7188
rect 11888 7142 11940 7148
rect 11900 7002 11928 7142
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11624 6854 11744 6882
rect 11796 6860 11848 6866
rect 11624 5778 11652 6854
rect 11796 6802 11848 6808
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6254 11744 6734
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11704 6112 11756 6118
rect 11808 6100 11836 6802
rect 11956 6556 12252 6576
rect 12012 6554 12036 6556
rect 12092 6554 12116 6556
rect 12172 6554 12196 6556
rect 12034 6502 12036 6554
rect 12098 6502 12110 6554
rect 12172 6502 12174 6554
rect 12012 6500 12036 6502
rect 12092 6500 12116 6502
rect 12172 6500 12196 6502
rect 11956 6480 12252 6500
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 11756 6072 11836 6100
rect 11704 6054 11756 6060
rect 11716 5778 11744 6054
rect 12084 5846 12112 6122
rect 12360 6118 12388 7210
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11624 5166 11652 5578
rect 11612 5160 11664 5166
rect 11716 5137 11744 5714
rect 12268 5710 12296 6054
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 11956 5468 12252 5488
rect 12012 5466 12036 5468
rect 12092 5466 12116 5468
rect 12172 5466 12196 5468
rect 12034 5414 12036 5466
rect 12098 5414 12110 5466
rect 12172 5414 12174 5466
rect 12012 5412 12036 5414
rect 12092 5412 12116 5414
rect 12172 5412 12196 5414
rect 11956 5392 12252 5412
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11612 5102 11664 5108
rect 11702 5128 11758 5137
rect 11702 5063 11758 5072
rect 11716 5030 11744 5063
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11716 4282 11744 4762
rect 11808 4758 11836 5238
rect 12360 5234 12388 5306
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12084 4826 12112 5170
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 12452 4690 12480 15150
rect 12544 10266 12572 15932
rect 12636 14414 12664 19110
rect 13372 18834 13400 21542
rect 13634 21520 13690 21542
rect 15212 21542 15530 21570
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17202 12756 17478
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12820 17066 12848 18022
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16658 12756 16934
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 15978 12756 16594
rect 12820 16046 12848 17002
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 14414 12848 15846
rect 12912 15434 12940 16526
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12912 14618 12940 14826
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12716 14272 12768 14278
rect 12622 14240 12678 14249
rect 12716 14214 12768 14220
rect 12622 14175 12678 14184
rect 12636 12832 12664 14175
rect 12728 13814 12756 14214
rect 12820 14006 12848 14350
rect 12912 14074 12940 14554
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12900 13864 12952 13870
rect 12728 13786 12848 13814
rect 12900 13806 12952 13812
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13462 12756 13670
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12820 12850 12848 13786
rect 12808 12844 12860 12850
rect 12636 12804 12756 12832
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12102 12664 12650
rect 12728 12646 12756 12804
rect 12808 12786 12860 12792
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11626 12664 12038
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12636 11354 12664 11562
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12728 11234 12756 12582
rect 12636 11206 12756 11234
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12544 9586 12572 10202
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12636 9466 12664 11206
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10198 12756 11086
rect 12820 10810 12848 12786
rect 12912 11082 12940 13806
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12808 10668 12860 10674
rect 13004 10656 13032 17138
rect 12808 10610 12860 10616
rect 12912 10628 13032 10656
rect 12820 10266 12848 10610
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12806 10160 12862 10169
rect 12912 10130 12940 10628
rect 12990 10568 13046 10577
rect 12990 10503 13046 10512
rect 12806 10095 12862 10104
rect 12900 10124 12952 10130
rect 12544 9438 12664 9466
rect 12544 8430 12572 9438
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12636 8634 12664 8842
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6254 12572 6598
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11532 4126 11652 4154
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11532 3670 11560 3878
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3194 11560 3606
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11624 3058 11652 4126
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11256 2417 11284 2926
rect 11716 2650 11744 4218
rect 11808 4146 11836 4490
rect 11956 4380 12252 4400
rect 12012 4378 12036 4380
rect 12092 4378 12116 4380
rect 12172 4378 12196 4380
rect 12034 4326 12036 4378
rect 12098 4326 12110 4378
rect 12172 4326 12174 4378
rect 12012 4324 12036 4326
rect 12092 4324 12116 4326
rect 12172 4324 12196 4326
rect 11956 4304 12252 4324
rect 12452 4154 12480 4626
rect 12544 4486 12572 6190
rect 12636 4593 12664 7890
rect 12622 4584 12678 4593
rect 12622 4519 12678 4528
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 12360 4126 12480 4154
rect 12360 3738 12388 4126
rect 12636 4010 12664 4218
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 11808 3194 11836 3674
rect 12728 3534 12756 8774
rect 12820 7546 12848 10095
rect 12900 10066 12952 10072
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 6934 12940 9386
rect 13004 8634 13032 10503
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5914 12848 6190
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3738 13032 4082
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 11956 3292 12252 3312
rect 12012 3290 12036 3292
rect 12092 3290 12116 3292
rect 12172 3290 12196 3292
rect 12034 3238 12036 3290
rect 12098 3238 12110 3290
rect 12172 3238 12174 3290
rect 12012 3236 12036 3238
rect 12092 3236 12116 3238
rect 12172 3236 12196 3238
rect 11956 3216 12252 3236
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 2650 12388 2994
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 11242 2408 11298 2417
rect 11242 2343 11298 2352
rect 11956 2204 12252 2224
rect 12012 2202 12036 2204
rect 12092 2202 12116 2204
rect 12172 2202 12196 2204
rect 12034 2150 12036 2202
rect 12098 2150 12110 2202
rect 12172 2150 12174 2202
rect 12012 2148 12036 2150
rect 12092 2148 12116 2150
rect 12172 2148 12196 2150
rect 11956 2128 12252 2148
rect 11152 196 11204 202
rect 11152 138 11204 144
rect 11426 82 11482 480
rect 10888 54 11482 82
rect 5906 0 5962 54
rect 7010 0 7066 54
rect 8114 0 8170 54
rect 9218 0 9274 54
rect 10322 0 10378 54
rect 11426 0 11482 54
rect 12530 82 12586 480
rect 12636 82 12664 3402
rect 13096 2650 13124 17818
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13188 13462 13216 14486
rect 13280 14249 13308 18158
rect 13372 18086 13400 18770
rect 13556 18222 13584 19110
rect 13728 18624 13780 18630
rect 13648 18584 13728 18612
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13266 14240 13322 14249
rect 13266 14175 13322 14184
rect 13372 14074 13400 17206
rect 13464 16454 13492 17614
rect 13556 16998 13584 17682
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16046 13492 16390
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13464 14385 13492 15982
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13556 14929 13584 15370
rect 13542 14920 13598 14929
rect 13542 14855 13598 14864
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13450 14376 13506 14385
rect 13450 14311 13506 14320
rect 13464 14278 13492 14311
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13188 9450 13216 12786
rect 13280 12306 13308 13874
rect 13556 13870 13584 14758
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13464 13274 13492 13806
rect 13556 13530 13584 13806
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13464 13246 13584 13274
rect 13556 13190 13584 13246
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13280 11898 13308 12242
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13280 11150 13308 11562
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13372 10996 13400 12854
rect 13280 10968 13400 10996
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 9110 13216 9386
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13280 8498 13308 10968
rect 13358 10840 13414 10849
rect 13358 10775 13414 10784
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13280 5778 13308 7142
rect 13372 6390 13400 10775
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13464 9654 13492 10066
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8294 13492 9318
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13464 6866 13492 7414
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13464 6458 13492 6802
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13280 5234 13308 5714
rect 13372 5234 13400 6326
rect 13556 5914 13584 13126
rect 13648 9178 13676 18584
rect 13728 18566 13780 18572
rect 13832 17241 13860 19110
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13818 17232 13874 17241
rect 14108 17202 14136 17478
rect 14384 17202 14412 18294
rect 13818 17167 13874 17176
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 13820 17128 13872 17134
rect 13872 17088 14044 17116
rect 13820 17070 13872 17076
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13740 16250 13768 16594
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15094 13768 15506
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13820 14952 13872 14958
rect 13726 14920 13782 14929
rect 13820 14894 13872 14900
rect 13726 14855 13782 14864
rect 13740 14346 13768 14855
rect 13832 14550 13860 14894
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13740 12374 13768 14282
rect 13818 13288 13874 13297
rect 13818 13223 13874 13232
rect 13832 12782 13860 13223
rect 13924 12986 13952 16730
rect 14016 16658 14044 17088
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14016 15910 14044 16594
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 14016 15570 14044 15846
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14016 15094 14044 15506
rect 14108 15162 14136 17138
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 14108 14346 14136 15098
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 14108 13433 14136 14282
rect 14094 13424 14150 13433
rect 14004 13388 14056 13394
rect 14094 13359 14150 13368
rect 14004 13330 14056 13336
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13740 11354 13768 12310
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 10169 13768 11290
rect 13726 10160 13782 10169
rect 13726 10095 13782 10104
rect 13832 9994 13860 12718
rect 14016 12714 14044 13330
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14108 11558 14136 12582
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 10470 14136 11494
rect 14200 11354 14228 15438
rect 14292 12442 14320 15914
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14292 11762 14320 12378
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14200 10674 14228 11290
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10198 14136 10406
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7206 13676 8230
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5794 13676 6938
rect 13740 6254 13768 9862
rect 14108 9382 14136 10134
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13832 8294 13860 9046
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8022 13860 8230
rect 13924 8090 13952 8366
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13832 7002 13860 7958
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 7002 14044 7278
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13464 5766 13676 5794
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13464 4758 13492 5766
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13636 5092 13688 5098
rect 13556 5052 13636 5080
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13464 4282 13492 4694
rect 13556 4486 13584 5052
rect 13636 5034 13688 5040
rect 14016 4690 14044 5646
rect 14200 5370 14228 6666
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13464 3942 13492 4218
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 2650 13492 3878
rect 13556 3670 13584 4422
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14108 3670 14136 3946
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 13556 3194 13584 3606
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 14108 3058 14136 3606
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13096 2446 13124 2586
rect 13358 2544 13414 2553
rect 13358 2479 13414 2488
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13004 134 13032 2246
rect 12530 54 12664 82
rect 12992 128 13044 134
rect 12992 70 13044 76
rect 13372 82 13400 2479
rect 13634 82 13690 480
rect 13372 54 13690 82
rect 14292 82 14320 4966
rect 14384 4146 14412 16934
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14476 15026 14504 15302
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9382 14504 9862
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14568 9110 14596 18294
rect 14660 17649 14688 19110
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14646 17640 14702 17649
rect 14646 17575 14702 17584
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14660 14890 14688 14962
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14660 14618 14688 14826
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14660 14074 14688 14554
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13462 14688 13738
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14660 11014 14688 12174
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14660 8906 14688 10950
rect 14752 9586 14780 18090
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14752 9178 14780 9522
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14844 7886 14872 18566
rect 15212 18426 15240 21542
rect 15474 21520 15530 21542
rect 16580 21548 16632 21554
rect 17314 21548 17370 22000
rect 19154 21570 19210 22000
rect 20994 21570 21050 22000
rect 17314 21520 17316 21548
rect 16580 21490 16632 21496
rect 17368 21520 17370 21548
rect 18984 21542 19210 21570
rect 17316 21490 17368 21496
rect 15622 19068 15918 19088
rect 15678 19066 15702 19068
rect 15758 19066 15782 19068
rect 15838 19066 15862 19068
rect 15700 19014 15702 19066
rect 15764 19014 15776 19066
rect 15838 19014 15840 19066
rect 15678 19012 15702 19014
rect 15758 19012 15782 19014
rect 15838 19012 15862 19014
rect 15622 18992 15918 19012
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 16040 18086 16068 18770
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 15622 17980 15918 18000
rect 15678 17978 15702 17980
rect 15758 17978 15782 17980
rect 15838 17978 15862 17980
rect 15700 17926 15702 17978
rect 15764 17926 15776 17978
rect 15838 17926 15840 17978
rect 15678 17924 15702 17926
rect 15758 17924 15782 17926
rect 15838 17924 15862 17926
rect 15622 17904 15918 17924
rect 16040 17785 16068 18022
rect 16026 17776 16082 17785
rect 16026 17711 16082 17720
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14476 5846 14504 7210
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6254 14872 6598
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14936 5914 14964 16526
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15120 14074 15148 14486
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15304 13546 15332 16934
rect 15396 14414 15424 17614
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15622 16892 15918 16912
rect 15678 16890 15702 16892
rect 15758 16890 15782 16892
rect 15838 16890 15862 16892
rect 15700 16838 15702 16890
rect 15764 16838 15776 16890
rect 15838 16838 15840 16890
rect 15678 16836 15702 16838
rect 15758 16836 15782 16838
rect 15838 16836 15862 16838
rect 15622 16816 15918 16836
rect 15622 15804 15918 15824
rect 15678 15802 15702 15804
rect 15758 15802 15782 15804
rect 15838 15802 15862 15804
rect 15700 15750 15702 15802
rect 15764 15750 15776 15802
rect 15838 15750 15840 15802
rect 15678 15748 15702 15750
rect 15758 15748 15782 15750
rect 15838 15748 15862 15750
rect 15622 15728 15918 15748
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15488 14822 15516 15506
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14414 15516 14758
rect 15622 14716 15918 14736
rect 15678 14714 15702 14716
rect 15758 14714 15782 14716
rect 15838 14714 15862 14716
rect 15700 14662 15702 14714
rect 15764 14662 15776 14714
rect 15838 14662 15840 14714
rect 15678 14660 15702 14662
rect 15758 14660 15782 14662
rect 15838 14660 15862 14662
rect 15622 14640 15918 14660
rect 15948 14618 15976 14826
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15396 14006 15424 14350
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 16040 13814 16068 17478
rect 16316 17270 16344 17682
rect 16304 17264 16356 17270
rect 16304 17206 16356 17212
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16132 15978 16160 16594
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16120 15972 16172 15978
rect 16172 15932 16252 15960
rect 16120 15914 16172 15920
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16132 14346 16160 15506
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16132 13938 16160 14282
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15948 13786 16068 13814
rect 15120 13518 15332 13546
rect 15120 13326 15148 13518
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15120 12442 15148 13262
rect 15212 12986 15240 13398
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15028 11354 15056 12310
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15028 10606 15056 11290
rect 15120 11286 15148 11494
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15120 10810 15148 11222
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15212 10470 15240 11086
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 9450 15240 10406
rect 15290 10160 15346 10169
rect 15290 10095 15346 10104
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 15028 8498 15056 9046
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15120 8090 15148 8910
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15212 7818 15240 9386
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15304 6866 15332 10095
rect 15396 9586 15424 12582
rect 15488 9654 15516 13738
rect 15622 13628 15918 13648
rect 15678 13626 15702 13628
rect 15758 13626 15782 13628
rect 15838 13626 15862 13628
rect 15700 13574 15702 13626
rect 15764 13574 15776 13626
rect 15838 13574 15840 13626
rect 15678 13572 15702 13574
rect 15758 13572 15782 13574
rect 15838 13572 15862 13574
rect 15622 13552 15918 13572
rect 15622 12540 15918 12560
rect 15678 12538 15702 12540
rect 15758 12538 15782 12540
rect 15838 12538 15862 12540
rect 15700 12486 15702 12538
rect 15764 12486 15776 12538
rect 15838 12486 15840 12538
rect 15678 12484 15702 12486
rect 15758 12484 15782 12486
rect 15838 12484 15862 12486
rect 15622 12464 15918 12484
rect 15622 11452 15918 11472
rect 15678 11450 15702 11452
rect 15758 11450 15782 11452
rect 15838 11450 15862 11452
rect 15700 11398 15702 11450
rect 15764 11398 15776 11450
rect 15838 11398 15840 11450
rect 15678 11396 15702 11398
rect 15758 11396 15782 11398
rect 15838 11396 15862 11398
rect 15622 11376 15918 11396
rect 15622 10364 15918 10384
rect 15678 10362 15702 10364
rect 15758 10362 15782 10364
rect 15838 10362 15862 10364
rect 15700 10310 15702 10362
rect 15764 10310 15776 10362
rect 15838 10310 15840 10362
rect 15678 10308 15702 10310
rect 15758 10308 15782 10310
rect 15838 10308 15862 10310
rect 15622 10288 15918 10308
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9722 15792 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15764 9489 15792 9658
rect 15750 9480 15806 9489
rect 15750 9415 15806 9424
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9110 15424 9318
rect 15622 9276 15918 9296
rect 15678 9274 15702 9276
rect 15758 9274 15782 9276
rect 15838 9274 15862 9276
rect 15700 9222 15702 9274
rect 15764 9222 15776 9274
rect 15838 9222 15840 9274
rect 15678 9220 15702 9222
rect 15758 9220 15782 9222
rect 15838 9220 15862 9222
rect 15622 9200 15918 9220
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15396 8634 15424 9046
rect 15844 8968 15896 8974
rect 15948 8956 15976 13786
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12238 16068 13262
rect 16132 12918 16160 13670
rect 16224 12968 16252 15932
rect 16316 15366 16344 15982
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 13190 16344 15302
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16224 12940 16344 12968
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11286 16068 12174
rect 16118 11384 16174 11393
rect 16118 11319 16174 11328
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16132 9994 16160 11319
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 15896 8928 15976 8956
rect 16028 8968 16080 8974
rect 15844 8910 15896 8916
rect 16028 8910 16080 8916
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 16040 8498 16068 8910
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 8022 15516 8230
rect 15622 8188 15918 8208
rect 15678 8186 15702 8188
rect 15758 8186 15782 8188
rect 15838 8186 15862 8188
rect 15700 8134 15702 8186
rect 15764 8134 15776 8186
rect 15838 8134 15840 8186
rect 15678 8132 15702 8134
rect 15758 8132 15782 8134
rect 15838 8132 15862 8134
rect 15622 8112 15918 8132
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 6458 15332 6802
rect 15396 6730 15424 7822
rect 15488 7546 15516 7958
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15622 7100 15918 7120
rect 15678 7098 15702 7100
rect 15758 7098 15782 7100
rect 15838 7098 15862 7100
rect 15700 7046 15702 7098
rect 15764 7046 15776 7098
rect 15838 7046 15840 7098
rect 15678 7044 15702 7046
rect 15758 7044 15782 7046
rect 15838 7044 15862 7046
rect 15622 7024 15918 7044
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15948 6390 15976 6802
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 16026 6352 16082 6361
rect 16026 6287 16082 6296
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14476 5370 14504 5782
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14660 4010 14688 5510
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4622 14780 5034
rect 14844 5030 14872 5578
rect 14936 5166 14964 5850
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5273 15240 5646
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15198 5264 15254 5273
rect 15198 5199 15254 5208
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 4729 14872 4966
rect 15120 4826 15148 5102
rect 15212 5098 15240 5199
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15212 4758 15240 5034
rect 15200 4752 15252 4758
rect 14830 4720 14886 4729
rect 15200 4694 15252 4700
rect 14830 4655 14886 4664
rect 15016 4684 15068 4690
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14844 4554 14872 4655
rect 15016 4626 15068 4632
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 15028 3738 15056 4626
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14568 2650 14596 2790
rect 14844 2650 14872 3470
rect 15120 2922 15148 3878
rect 15212 3670 15240 4694
rect 15304 4690 15332 5306
rect 15488 4826 15516 6190
rect 15622 6012 15918 6032
rect 15678 6010 15702 6012
rect 15758 6010 15782 6012
rect 15838 6010 15862 6012
rect 15700 5958 15702 6010
rect 15764 5958 15776 6010
rect 15838 5958 15840 6010
rect 15678 5956 15702 5958
rect 15758 5956 15782 5958
rect 15838 5956 15862 5958
rect 15622 5936 15918 5956
rect 16040 5574 16068 6287
rect 16132 5914 16160 9522
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16224 5658 16252 12786
rect 16316 11830 16344 12940
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16304 11620 16356 11626
rect 16304 11562 16356 11568
rect 16316 7546 16344 11562
rect 16408 10266 16436 18022
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 14074 16528 14418
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16408 9654 16436 10202
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16500 8090 16528 13874
rect 16592 13530 16620 21490
rect 17328 21459 17356 21490
rect 17498 18728 17554 18737
rect 17498 18663 17554 18672
rect 16762 18048 16818 18057
rect 16762 17983 16818 17992
rect 16776 17814 16804 17983
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16592 12782 16620 12854
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16592 10266 16620 10610
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16684 10130 16712 15914
rect 16776 14482 16804 16186
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16776 13326 16804 13942
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16868 12850 16896 16526
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15570 16988 15846
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16960 14822 16988 15506
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16960 13326 16988 14554
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16684 9722 16712 10066
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16592 9178 16620 9386
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16670 8936 16726 8945
rect 16670 8871 16726 8880
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16316 6866 16344 7482
rect 16500 7342 16528 8026
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6186 16528 6598
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16316 5914 16344 6122
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16132 5630 16252 5658
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16040 5302 16068 5510
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15622 4924 15918 4944
rect 15678 4922 15702 4924
rect 15758 4922 15782 4924
rect 15838 4922 15862 4924
rect 15700 4870 15702 4922
rect 15764 4870 15776 4922
rect 15838 4870 15840 4922
rect 15678 4868 15702 4870
rect 15758 4868 15782 4870
rect 15838 4868 15862 4870
rect 15622 4848 15918 4868
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15292 4684 15344 4690
rect 16040 4672 16068 5238
rect 15292 4626 15344 4632
rect 15948 4644 16068 4672
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15396 3670 15424 4558
rect 15948 4486 15976 4644
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15948 4282 15976 4422
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16040 3942 16068 4490
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15488 3670 15516 3878
rect 15622 3836 15918 3856
rect 15678 3834 15702 3836
rect 15758 3834 15782 3836
rect 15838 3834 15862 3836
rect 15700 3782 15702 3834
rect 15764 3782 15776 3834
rect 15838 3782 15840 3834
rect 15678 3780 15702 3782
rect 15758 3780 15782 3782
rect 15838 3780 15862 3782
rect 15622 3760 15918 3780
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15488 3194 15516 3606
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15936 3120 15988 3126
rect 16040 3097 16068 3878
rect 15936 3062 15988 3068
rect 16026 3088 16082 3097
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15304 2650 15332 2926
rect 15622 2748 15918 2768
rect 15678 2746 15702 2748
rect 15758 2746 15782 2748
rect 15838 2746 15862 2748
rect 15700 2694 15702 2746
rect 15764 2694 15776 2746
rect 15838 2694 15840 2746
rect 15678 2692 15702 2694
rect 15758 2692 15782 2694
rect 15838 2692 15862 2694
rect 15622 2672 15918 2692
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 14738 82 14794 480
rect 14292 54 14794 82
rect 12530 0 12586 54
rect 13634 0 13690 54
rect 14738 0 14794 54
rect 15842 82 15898 480
rect 15948 82 15976 3062
rect 16026 3023 16082 3032
rect 16132 2650 16160 5630
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16224 4060 16252 4762
rect 16396 4072 16448 4078
rect 16224 4032 16396 4060
rect 16396 4014 16448 4020
rect 16408 3738 16436 4014
rect 16500 3738 16528 6122
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16592 5098 16620 5170
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4826 16620 5034
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16592 3602 16620 3946
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16592 3194 16620 3538
rect 16684 3466 16712 8871
rect 16776 7954 16804 11562
rect 16868 9042 16896 12650
rect 16960 11762 16988 13126
rect 17052 12442 17080 15438
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16960 11150 16988 11698
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 17052 10742 17080 11630
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16960 10130 16988 10474
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 17052 9654 17080 10678
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8634 16896 8978
rect 17144 8956 17172 16526
rect 17236 10674 17264 17546
rect 17420 16998 17448 17682
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17316 16040 17368 16046
rect 17420 16017 17448 16934
rect 17316 15982 17368 15988
rect 17406 16008 17462 16017
rect 17328 12850 17356 15982
rect 17406 15943 17462 15952
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17420 15162 17448 15370
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17420 14958 17448 15098
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 14482 17448 14758
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17420 13870 17448 14418
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17512 13802 17540 18663
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18524 18057 18552 18090
rect 18510 18048 18566 18057
rect 18510 17983 18566 17992
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18708 17649 18736 17682
rect 18694 17640 18750 17649
rect 18694 17575 18750 17584
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17406 13696 17462 13705
rect 17406 13631 17462 13640
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 12442 17356 12582
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 11898 17356 12378
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17328 11626 17356 11834
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17328 11286 17356 11562
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17328 10554 17356 11086
rect 17052 8928 17172 8956
rect 17236 10526 17356 10554
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16776 7546 16804 7890
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16776 5846 16804 6122
rect 16764 5840 16816 5846
rect 16764 5782 16816 5788
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 3942 16896 4422
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3602 16896 3878
rect 16960 3670 16988 8026
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16868 2922 16896 3538
rect 16960 3058 16988 3606
rect 17052 3448 17080 8928
rect 17130 4584 17186 4593
rect 17130 4519 17186 4528
rect 17144 4486 17172 4519
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17132 3460 17184 3466
rect 17052 3420 17132 3448
rect 17132 3402 17184 3408
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16132 2446 16160 2586
rect 16500 2582 16528 2790
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16960 2378 16988 2994
rect 17236 2582 17264 10526
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10198 17356 10406
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17328 9382 17356 10134
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 9110 17356 9318
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17328 8294 17356 9046
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17328 8022 17356 8230
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17328 7206 17356 7958
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17328 6848 17356 7142
rect 17420 7002 17448 13631
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17512 12986 17540 13262
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 8090 17540 12786
rect 17604 9586 17632 17478
rect 18064 17134 18092 17478
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17788 15570 17816 17070
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17788 15473 17816 15506
rect 17774 15464 17830 15473
rect 17774 15399 17830 15408
rect 17788 15162 17816 15399
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17776 15156 17828 15162
rect 17696 15116 17776 15144
rect 17696 13569 17724 15116
rect 17776 15098 17828 15104
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17682 13560 17738 13569
rect 17682 13495 17738 13504
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17696 12374 17724 13398
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17788 10062 17816 14962
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17880 11218 17908 14554
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10810 17908 11154
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9178 17816 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8634 17908 8910
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17972 7886 18000 15302
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18340 14958 18368 15030
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 13841 18184 14758
rect 18248 14482 18276 14894
rect 18340 14550 18368 14894
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18142 13832 18198 13841
rect 18142 13767 18198 13776
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 11354 18092 12582
rect 18156 11762 18184 13670
rect 18248 13530 18276 14418
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 13938 18368 14214
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18236 13184 18288 13190
rect 18340 13172 18368 13874
rect 18288 13144 18368 13172
rect 18236 13126 18288 13132
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18156 11354 18184 11698
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18064 10810 18092 11290
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18156 9178 18184 9522
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17408 6860 17460 6866
rect 17328 6820 17408 6848
rect 17408 6802 17460 6808
rect 17420 6118 17448 6802
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17788 6458 17816 6734
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17972 6186 18000 6394
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5846 17448 6054
rect 17972 5914 18000 6122
rect 18156 5914 18184 7210
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17880 5030 17908 5782
rect 18156 5234 18184 5850
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17880 4758 17908 4966
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17774 4176 17830 4185
rect 17774 4111 17830 4120
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17328 3534 17356 3946
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17328 2650 17356 3470
rect 17788 3194 17816 4111
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17788 2922 17816 3130
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17788 2650 17816 2858
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 17972 1329 18000 4218
rect 18156 4010 18184 4558
rect 18248 4078 18276 13126
rect 18432 10062 18460 17002
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18524 11354 18552 16934
rect 18616 12918 18644 17478
rect 18708 16998 18736 17575
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18708 16658 18736 16934
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18708 12374 18736 13330
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18524 10742 18552 11290
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18432 9654 18460 9998
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18432 7954 18460 8570
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18524 8022 18552 8230
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18432 7546 18460 7890
rect 18524 7750 18552 7958
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 7546 18552 7686
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18432 7206 18460 7482
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18524 7002 18552 7482
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18616 4758 18644 11766
rect 18800 9194 18828 14826
rect 18892 13326 18920 15846
rect 18984 15706 19012 21542
rect 19154 21520 19210 21542
rect 20640 21542 21050 21570
rect 19614 20496 19670 20505
rect 19614 20431 19670 20440
rect 19289 19612 19585 19632
rect 19345 19610 19369 19612
rect 19425 19610 19449 19612
rect 19505 19610 19529 19612
rect 19367 19558 19369 19610
rect 19431 19558 19443 19610
rect 19505 19558 19507 19610
rect 19345 19556 19369 19558
rect 19425 19556 19449 19558
rect 19505 19556 19529 19558
rect 19289 19536 19585 19556
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19168 17746 19196 18906
rect 19289 18524 19585 18544
rect 19345 18522 19369 18524
rect 19425 18522 19449 18524
rect 19505 18522 19529 18524
rect 19367 18470 19369 18522
rect 19431 18470 19443 18522
rect 19505 18470 19507 18522
rect 19345 18468 19369 18470
rect 19425 18468 19449 18470
rect 19505 18468 19529 18470
rect 19289 18448 19585 18468
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19076 17134 19104 17478
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18984 13870 19012 14418
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 19076 13326 19104 17070
rect 19168 15570 19196 17682
rect 19289 17436 19585 17456
rect 19345 17434 19369 17436
rect 19425 17434 19449 17436
rect 19505 17434 19529 17436
rect 19367 17382 19369 17434
rect 19431 17382 19443 17434
rect 19505 17382 19507 17434
rect 19345 17380 19369 17382
rect 19425 17380 19449 17382
rect 19505 17380 19529 17382
rect 19289 17360 19585 17380
rect 19628 17338 19656 20431
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19720 17338 19748 17682
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19522 16960 19578 16969
rect 19522 16895 19578 16904
rect 19536 16794 19564 16895
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19289 16348 19585 16368
rect 19345 16346 19369 16348
rect 19425 16346 19449 16348
rect 19505 16346 19529 16348
rect 19367 16294 19369 16346
rect 19431 16294 19443 16346
rect 19505 16294 19507 16346
rect 19345 16292 19369 16294
rect 19425 16292 19449 16294
rect 19505 16292 19529 16294
rect 19289 16272 19585 16292
rect 19628 16250 19656 16594
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19708 15972 19760 15978
rect 19708 15914 19760 15920
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19168 15162 19196 15506
rect 19289 15260 19585 15280
rect 19345 15258 19369 15260
rect 19425 15258 19449 15260
rect 19505 15258 19529 15260
rect 19367 15206 19369 15258
rect 19431 15206 19443 15258
rect 19505 15206 19507 15258
rect 19345 15204 19369 15206
rect 19425 15204 19449 15206
rect 19505 15204 19529 15206
rect 19289 15184 19585 15204
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19168 15065 19196 15098
rect 19154 15056 19210 15065
rect 19154 14991 19210 15000
rect 19154 14512 19210 14521
rect 19154 14447 19210 14456
rect 19168 13870 19196 14447
rect 19289 14172 19585 14192
rect 19345 14170 19369 14172
rect 19425 14170 19449 14172
rect 19505 14170 19529 14172
rect 19367 14118 19369 14170
rect 19431 14118 19443 14170
rect 19505 14118 19507 14170
rect 19345 14116 19369 14118
rect 19425 14116 19449 14118
rect 19505 14116 19529 14118
rect 19289 14096 19585 14116
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 18892 12986 18920 13262
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18984 12238 19012 12786
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18984 11694 19012 12174
rect 19076 12170 19104 13262
rect 19289 13084 19585 13104
rect 19345 13082 19369 13084
rect 19425 13082 19449 13084
rect 19505 13082 19529 13084
rect 19367 13030 19369 13082
rect 19431 13030 19443 13082
rect 19505 13030 19507 13082
rect 19345 13028 19369 13030
rect 19425 13028 19449 13030
rect 19505 13028 19529 13030
rect 19289 13008 19585 13028
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 19076 11642 19104 12106
rect 19168 11898 19196 12378
rect 19289 11996 19585 12016
rect 19345 11994 19369 11996
rect 19425 11994 19449 11996
rect 19505 11994 19529 11996
rect 19367 11942 19369 11994
rect 19431 11942 19443 11994
rect 19505 11942 19507 11994
rect 19345 11940 19369 11942
rect 19425 11940 19449 11942
rect 19505 11940 19529 11942
rect 19289 11920 19585 11940
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19076 11614 19196 11642
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11286 19104 11494
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18892 10674 18920 11018
rect 19076 10810 19104 11222
rect 19168 11150 19196 11614
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19289 10908 19585 10928
rect 19345 10906 19369 10908
rect 19425 10906 19449 10908
rect 19505 10906 19529 10908
rect 19367 10854 19369 10906
rect 19431 10854 19443 10906
rect 19505 10854 19507 10906
rect 19345 10852 19369 10854
rect 19425 10852 19449 10854
rect 19505 10852 19529 10854
rect 19289 10832 19585 10852
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 10062 18920 10610
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18892 9586 18920 9998
rect 19076 9722 19104 10134
rect 19289 9820 19585 9840
rect 19345 9818 19369 9820
rect 19425 9818 19449 9820
rect 19505 9818 19529 9820
rect 19367 9766 19369 9818
rect 19431 9766 19443 9818
rect 19505 9766 19507 9818
rect 19345 9764 19369 9766
rect 19425 9764 19449 9766
rect 19505 9764 19529 9766
rect 19289 9744 19585 9764
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 18708 9166 18828 9194
rect 18708 7410 18736 9166
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18800 8634 18828 9046
rect 19536 8974 19564 9318
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 19076 8362 19104 8842
rect 19289 8732 19585 8752
rect 19345 8730 19369 8732
rect 19425 8730 19449 8732
rect 19505 8730 19529 8732
rect 19367 8678 19369 8730
rect 19431 8678 19443 8730
rect 19505 8678 19507 8730
rect 19345 8676 19369 8678
rect 19425 8676 19449 8678
rect 19505 8676 19529 8678
rect 19289 8656 19585 8676
rect 19628 8634 19656 13670
rect 19720 10266 19748 15914
rect 20640 14006 20668 21542
rect 20994 21520 21050 21542
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21560 15609 21588 15642
rect 21546 15600 21602 15609
rect 21546 15535 21602 15544
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 20074 9616 20130 9625
rect 20074 9551 20130 9560
rect 20088 9518 20116 9551
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18800 7478 18828 7822
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18892 7410 18920 7822
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18708 7002 18736 7346
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18800 6458 18828 6870
rect 18892 6798 18920 7346
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18892 5710 18920 6734
rect 19076 6322 19104 8298
rect 19289 7644 19585 7664
rect 19345 7642 19369 7644
rect 19425 7642 19449 7644
rect 19505 7642 19529 7644
rect 19367 7590 19369 7642
rect 19431 7590 19443 7642
rect 19505 7590 19507 7642
rect 19345 7588 19369 7590
rect 19425 7588 19449 7590
rect 19505 7588 19529 7590
rect 19289 7568 19585 7588
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19289 6556 19585 6576
rect 19345 6554 19369 6556
rect 19425 6554 19449 6556
rect 19505 6554 19529 6556
rect 19367 6502 19369 6554
rect 19431 6502 19443 6554
rect 19505 6502 19507 6554
rect 19345 6500 19369 6502
rect 19425 6500 19449 6502
rect 19505 6500 19529 6502
rect 19289 6480 19585 6500
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 5302 18920 5646
rect 18984 5574 19012 6122
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 5370 19012 5510
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18616 4629 18644 4694
rect 19076 4154 19104 5646
rect 19168 5012 19196 5782
rect 19352 5710 19380 6122
rect 19628 6118 19656 6666
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19289 5468 19585 5488
rect 19345 5466 19369 5468
rect 19425 5466 19449 5468
rect 19505 5466 19529 5468
rect 19367 5414 19369 5466
rect 19431 5414 19443 5466
rect 19505 5414 19507 5466
rect 19345 5412 19369 5414
rect 19425 5412 19449 5414
rect 19505 5412 19529 5414
rect 19289 5392 19585 5412
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19248 5024 19300 5030
rect 19168 4984 19248 5012
rect 19248 4966 19300 4972
rect 19260 4826 19288 4966
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19444 4690 19472 5102
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19444 4593 19472 4626
rect 19154 4584 19210 4593
rect 19154 4519 19210 4528
rect 19430 4584 19486 4593
rect 19430 4519 19486 4528
rect 19168 4282 19196 4519
rect 19289 4380 19585 4400
rect 19345 4378 19369 4380
rect 19425 4378 19449 4380
rect 19505 4378 19529 4380
rect 19367 4326 19369 4378
rect 19431 4326 19443 4378
rect 19505 4326 19507 4378
rect 19345 4324 19369 4326
rect 19425 4324 19449 4326
rect 19505 4324 19529 4326
rect 19289 4304 19585 4324
rect 19628 4282 19656 6054
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20088 4282 20116 4694
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 19076 4126 19196 4154
rect 20088 4153 20116 4218
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18248 3738 18276 4014
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18800 3738 18828 3946
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18064 3040 18092 3674
rect 18892 3505 18920 3946
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18878 3496 18934 3505
rect 18878 3431 18934 3440
rect 18984 3194 19012 3606
rect 19168 3534 19196 4126
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 19076 3126 19104 3402
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18144 3052 18196 3058
rect 18064 3012 18144 3040
rect 18144 2994 18196 3000
rect 19168 2310 19196 3470
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 19289 3292 19585 3312
rect 19345 3290 19369 3292
rect 19425 3290 19449 3292
rect 19505 3290 19529 3292
rect 19367 3238 19369 3290
rect 19431 3238 19443 3290
rect 19505 3238 19507 3290
rect 19345 3236 19369 3238
rect 19425 3236 19449 3238
rect 19505 3236 19529 3238
rect 19289 3216 19585 3236
rect 20088 2990 20116 3334
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19289 2204 19585 2224
rect 19345 2202 19369 2204
rect 19425 2202 19449 2204
rect 19505 2202 19529 2204
rect 19367 2150 19369 2202
rect 19431 2150 19443 2202
rect 19505 2150 19507 2202
rect 19345 2148 19369 2150
rect 19425 2148 19449 2150
rect 19505 2148 19529 2150
rect 19289 2128 19585 2148
rect 18144 2032 18196 2038
rect 18144 1974 18196 1980
rect 17958 1320 18014 1329
rect 17958 1255 18014 1264
rect 15842 54 15976 82
rect 16946 60 17002 480
rect 15842 0 15898 54
rect 16946 8 16948 60
rect 17000 8 17002 60
rect 16946 0 17002 8
rect 18050 82 18106 480
rect 18156 82 18184 1974
rect 20350 1456 20406 1465
rect 20350 1391 20406 1400
rect 18050 54 18184 82
rect 19154 128 19210 480
rect 19154 76 19156 128
rect 19208 76 19210 128
rect 18050 0 18106 54
rect 19154 0 19210 76
rect 20258 82 20314 480
rect 20364 82 20392 1391
rect 20258 54 20392 82
rect 21362 82 21418 480
rect 21468 82 21496 10202
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21560 8265 21588 9454
rect 21546 8256 21602 8265
rect 21546 8191 21602 8200
rect 21546 6352 21602 6361
rect 21546 6287 21602 6296
rect 21560 4758 21588 6287
rect 21548 4752 21600 4758
rect 21548 4694 21600 4700
rect 21362 54 21496 82
rect 20258 0 20314 54
rect 21362 0 21418 54
<< via2 >>
rect 110 17312 166 17368
rect 1490 20440 1546 20496
rect 1306 18672 1362 18728
rect 754 17040 810 17096
rect 110 15544 166 15600
rect 110 11872 166 11928
rect 386 9152 442 9208
rect 110 8472 166 8528
rect 110 8200 166 8256
rect 1582 13368 1638 13424
rect 1674 10648 1730 10704
rect 1582 9424 1638 9480
rect 1766 4256 1822 4312
rect 1582 3168 1638 3224
rect 2318 5208 2374 5264
rect 2318 4120 2374 4176
rect 3238 15272 3294 15328
rect 2962 9560 3018 9616
rect 2870 6296 2926 6352
rect 3422 10648 3478 10704
rect 2962 5208 3018 5264
rect 2778 4664 2834 4720
rect 2042 2896 2098 2952
rect 1950 2352 2006 2408
rect 4066 11600 4122 11656
rect 3882 9968 3938 10024
rect 4622 19610 4678 19612
rect 4702 19610 4758 19612
rect 4782 19610 4838 19612
rect 4862 19610 4918 19612
rect 4622 19558 4648 19610
rect 4648 19558 4678 19610
rect 4702 19558 4712 19610
rect 4712 19558 4758 19610
rect 4782 19558 4828 19610
rect 4828 19558 4838 19610
rect 4862 19558 4892 19610
rect 4892 19558 4918 19610
rect 4622 19556 4678 19558
rect 4702 19556 4758 19558
rect 4782 19556 4838 19558
rect 4862 19556 4918 19558
rect 4622 18522 4678 18524
rect 4702 18522 4758 18524
rect 4782 18522 4838 18524
rect 4862 18522 4918 18524
rect 4622 18470 4648 18522
rect 4648 18470 4678 18522
rect 4702 18470 4712 18522
rect 4712 18470 4758 18522
rect 4782 18470 4828 18522
rect 4828 18470 4838 18522
rect 4862 18470 4892 18522
rect 4892 18470 4918 18522
rect 4622 18468 4678 18470
rect 4702 18468 4758 18470
rect 4782 18468 4838 18470
rect 4862 18468 4918 18470
rect 8289 19066 8345 19068
rect 8369 19066 8425 19068
rect 8449 19066 8505 19068
rect 8529 19066 8585 19068
rect 8289 19014 8315 19066
rect 8315 19014 8345 19066
rect 8369 19014 8379 19066
rect 8379 19014 8425 19066
rect 8449 19014 8495 19066
rect 8495 19014 8505 19066
rect 8529 19014 8559 19066
rect 8559 19014 8585 19066
rect 8289 19012 8345 19014
rect 8369 19012 8425 19014
rect 8449 19012 8505 19014
rect 8529 19012 8585 19014
rect 6366 17740 6422 17776
rect 6366 17720 6368 17740
rect 6368 17720 6420 17740
rect 6420 17720 6422 17740
rect 4526 17584 4582 17640
rect 4622 17434 4678 17436
rect 4702 17434 4758 17436
rect 4782 17434 4838 17436
rect 4862 17434 4918 17436
rect 4622 17382 4648 17434
rect 4648 17382 4678 17434
rect 4702 17382 4712 17434
rect 4712 17382 4758 17434
rect 4782 17382 4828 17434
rect 4828 17382 4838 17434
rect 4862 17382 4892 17434
rect 4892 17382 4918 17434
rect 4622 17380 4678 17382
rect 4702 17380 4758 17382
rect 4782 17380 4838 17382
rect 4862 17380 4918 17382
rect 6642 17584 6698 17640
rect 4622 16346 4678 16348
rect 4702 16346 4758 16348
rect 4782 16346 4838 16348
rect 4862 16346 4918 16348
rect 4622 16294 4648 16346
rect 4648 16294 4678 16346
rect 4702 16294 4712 16346
rect 4712 16294 4758 16346
rect 4782 16294 4828 16346
rect 4828 16294 4838 16346
rect 4862 16294 4892 16346
rect 4892 16294 4918 16346
rect 4622 16292 4678 16294
rect 4702 16292 4758 16294
rect 4782 16292 4838 16294
rect 4862 16292 4918 16294
rect 4434 15272 4490 15328
rect 4622 15258 4678 15260
rect 4702 15258 4758 15260
rect 4782 15258 4838 15260
rect 4862 15258 4918 15260
rect 4622 15206 4648 15258
rect 4648 15206 4678 15258
rect 4702 15206 4712 15258
rect 4712 15206 4758 15258
rect 4782 15206 4828 15258
rect 4828 15206 4838 15258
rect 4862 15206 4892 15258
rect 4892 15206 4918 15258
rect 4622 15204 4678 15206
rect 4702 15204 4758 15206
rect 4782 15204 4838 15206
rect 4862 15204 4918 15206
rect 3606 5072 3662 5128
rect 4622 14170 4678 14172
rect 4702 14170 4758 14172
rect 4782 14170 4838 14172
rect 4862 14170 4918 14172
rect 4622 14118 4648 14170
rect 4648 14118 4678 14170
rect 4702 14118 4712 14170
rect 4712 14118 4758 14170
rect 4782 14118 4828 14170
rect 4828 14118 4838 14170
rect 4862 14118 4892 14170
rect 4892 14118 4918 14170
rect 4622 14116 4678 14118
rect 4702 14116 4758 14118
rect 4782 14116 4838 14118
rect 4862 14116 4918 14118
rect 4526 13368 4582 13424
rect 4622 13082 4678 13084
rect 4702 13082 4758 13084
rect 4782 13082 4838 13084
rect 4862 13082 4918 13084
rect 4622 13030 4648 13082
rect 4648 13030 4678 13082
rect 4702 13030 4712 13082
rect 4712 13030 4758 13082
rect 4782 13030 4828 13082
rect 4828 13030 4838 13082
rect 4862 13030 4892 13082
rect 4892 13030 4918 13082
rect 4622 13028 4678 13030
rect 4702 13028 4758 13030
rect 4782 13028 4838 13030
rect 4862 13028 4918 13030
rect 4622 11994 4678 11996
rect 4702 11994 4758 11996
rect 4782 11994 4838 11996
rect 4862 11994 4918 11996
rect 4622 11942 4648 11994
rect 4648 11942 4678 11994
rect 4702 11942 4712 11994
rect 4712 11942 4758 11994
rect 4782 11942 4828 11994
rect 4828 11942 4838 11994
rect 4862 11942 4892 11994
rect 4892 11942 4918 11994
rect 4622 11940 4678 11942
rect 4702 11940 4758 11942
rect 4782 11940 4838 11942
rect 4862 11940 4918 11942
rect 5262 14456 5318 14512
rect 4622 10906 4678 10908
rect 4702 10906 4758 10908
rect 4782 10906 4838 10908
rect 4862 10906 4918 10908
rect 4622 10854 4648 10906
rect 4648 10854 4678 10906
rect 4702 10854 4712 10906
rect 4712 10854 4758 10906
rect 4782 10854 4828 10906
rect 4828 10854 4838 10906
rect 4862 10854 4892 10906
rect 4892 10854 4918 10906
rect 4622 10852 4678 10854
rect 4702 10852 4758 10854
rect 4782 10852 4838 10854
rect 4862 10852 4918 10854
rect 4622 9818 4678 9820
rect 4702 9818 4758 9820
rect 4782 9818 4838 9820
rect 4862 9818 4918 9820
rect 4622 9766 4648 9818
rect 4648 9766 4678 9818
rect 4702 9766 4712 9818
rect 4712 9766 4758 9818
rect 4782 9766 4828 9818
rect 4828 9766 4838 9818
rect 4862 9766 4892 9818
rect 4892 9766 4918 9818
rect 4622 9764 4678 9766
rect 4702 9764 4758 9766
rect 4782 9764 4838 9766
rect 4862 9764 4918 9766
rect 4434 9152 4490 9208
rect 4622 8730 4678 8732
rect 4702 8730 4758 8732
rect 4782 8730 4838 8732
rect 4862 8730 4918 8732
rect 4622 8678 4648 8730
rect 4648 8678 4678 8730
rect 4702 8678 4712 8730
rect 4712 8678 4758 8730
rect 4782 8678 4828 8730
rect 4828 8678 4838 8730
rect 4862 8678 4892 8730
rect 4892 8678 4918 8730
rect 4622 8676 4678 8678
rect 4702 8676 4758 8678
rect 4782 8676 4838 8678
rect 4862 8676 4918 8678
rect 4622 7642 4678 7644
rect 4702 7642 4758 7644
rect 4782 7642 4838 7644
rect 4862 7642 4918 7644
rect 4622 7590 4648 7642
rect 4648 7590 4678 7642
rect 4702 7590 4712 7642
rect 4712 7590 4758 7642
rect 4782 7590 4828 7642
rect 4828 7590 4838 7642
rect 4862 7590 4892 7642
rect 4892 7590 4918 7642
rect 4622 7588 4678 7590
rect 4702 7588 4758 7590
rect 4782 7588 4838 7590
rect 4862 7588 4918 7590
rect 4250 6704 4306 6760
rect 4066 4528 4122 4584
rect 4250 4256 4306 4312
rect 4622 6554 4678 6556
rect 4702 6554 4758 6556
rect 4782 6554 4838 6556
rect 4862 6554 4918 6556
rect 4622 6502 4648 6554
rect 4648 6502 4678 6554
rect 4702 6502 4712 6554
rect 4712 6502 4758 6554
rect 4782 6502 4828 6554
rect 4828 6502 4838 6554
rect 4862 6502 4892 6554
rect 4892 6502 4918 6554
rect 4622 6500 4678 6502
rect 4702 6500 4758 6502
rect 4782 6500 4838 6502
rect 4862 6500 4918 6502
rect 4622 5466 4678 5468
rect 4702 5466 4758 5468
rect 4782 5466 4838 5468
rect 4862 5466 4918 5468
rect 4622 5414 4648 5466
rect 4648 5414 4678 5466
rect 4702 5414 4712 5466
rect 4712 5414 4758 5466
rect 4782 5414 4828 5466
rect 4828 5414 4838 5466
rect 4862 5414 4892 5466
rect 4892 5414 4918 5466
rect 4622 5412 4678 5414
rect 4702 5412 4758 5414
rect 4782 5412 4838 5414
rect 4862 5412 4918 5414
rect 5446 9968 5502 10024
rect 5262 9560 5318 9616
rect 4250 3984 4306 4040
rect 2778 1400 2834 1456
rect 5630 8472 5686 8528
rect 5262 5616 5318 5672
rect 5262 5208 5318 5264
rect 5078 4936 5134 4992
rect 4622 4378 4678 4380
rect 4702 4378 4758 4380
rect 4782 4378 4838 4380
rect 4862 4378 4918 4380
rect 4622 4326 4648 4378
rect 4648 4326 4678 4378
rect 4702 4326 4712 4378
rect 4712 4326 4758 4378
rect 4782 4326 4828 4378
rect 4828 4326 4838 4378
rect 4862 4326 4892 4378
rect 4892 4326 4918 4378
rect 4622 4324 4678 4326
rect 4702 4324 4758 4326
rect 4782 4324 4838 4326
rect 4862 4324 4918 4326
rect 5354 4392 5410 4448
rect 4622 3290 4678 3292
rect 4702 3290 4758 3292
rect 4782 3290 4838 3292
rect 4862 3290 4918 3292
rect 4622 3238 4648 3290
rect 4648 3238 4678 3290
rect 4702 3238 4712 3290
rect 4712 3238 4758 3290
rect 4782 3238 4828 3290
rect 4828 3238 4838 3290
rect 4862 3238 4892 3290
rect 4892 3238 4918 3290
rect 4622 3236 4678 3238
rect 4702 3236 4758 3238
rect 4782 3236 4838 3238
rect 4862 3236 4918 3238
rect 4618 2488 4674 2544
rect 4622 2202 4678 2204
rect 4702 2202 4758 2204
rect 4782 2202 4838 2204
rect 4862 2202 4918 2204
rect 4622 2150 4648 2202
rect 4648 2150 4678 2202
rect 4702 2150 4712 2202
rect 4712 2150 4758 2202
rect 4782 2150 4828 2202
rect 4828 2150 4838 2202
rect 4862 2150 4892 2202
rect 4892 2150 4918 2202
rect 4622 2148 4678 2150
rect 4702 2148 4758 2150
rect 4782 2148 4838 2150
rect 4862 2148 4918 2150
rect 6642 15988 6644 16008
rect 6644 15988 6696 16008
rect 6696 15988 6698 16008
rect 6642 15952 6698 15988
rect 6734 9560 6790 9616
rect 7746 16904 7802 16960
rect 7930 14456 7986 14512
rect 7838 13504 7894 13560
rect 8022 13368 8078 13424
rect 8289 17978 8345 17980
rect 8369 17978 8425 17980
rect 8449 17978 8505 17980
rect 8529 17978 8585 17980
rect 8289 17926 8315 17978
rect 8315 17926 8345 17978
rect 8369 17926 8379 17978
rect 8379 17926 8425 17978
rect 8449 17926 8495 17978
rect 8495 17926 8505 17978
rect 8529 17926 8559 17978
rect 8559 17926 8585 17978
rect 8289 17924 8345 17926
rect 8369 17924 8425 17926
rect 8449 17924 8505 17926
rect 8529 17924 8585 17926
rect 8758 16904 8814 16960
rect 8289 16890 8345 16892
rect 8369 16890 8425 16892
rect 8449 16890 8505 16892
rect 8529 16890 8585 16892
rect 8289 16838 8315 16890
rect 8315 16838 8345 16890
rect 8369 16838 8379 16890
rect 8379 16838 8425 16890
rect 8449 16838 8495 16890
rect 8495 16838 8505 16890
rect 8529 16838 8559 16890
rect 8559 16838 8585 16890
rect 8289 16836 8345 16838
rect 8369 16836 8425 16838
rect 8449 16836 8505 16838
rect 8529 16836 8585 16838
rect 8850 16224 8906 16280
rect 8289 15802 8345 15804
rect 8369 15802 8425 15804
rect 8449 15802 8505 15804
rect 8529 15802 8585 15804
rect 8289 15750 8315 15802
rect 8315 15750 8345 15802
rect 8369 15750 8379 15802
rect 8379 15750 8425 15802
rect 8449 15750 8495 15802
rect 8495 15750 8505 15802
rect 8529 15750 8559 15802
rect 8559 15750 8585 15802
rect 8289 15748 8345 15750
rect 8369 15748 8425 15750
rect 8449 15748 8505 15750
rect 8529 15748 8585 15750
rect 7838 9424 7894 9480
rect 8289 14714 8345 14716
rect 8369 14714 8425 14716
rect 8449 14714 8505 14716
rect 8529 14714 8585 14716
rect 8289 14662 8315 14714
rect 8315 14662 8345 14714
rect 8369 14662 8379 14714
rect 8379 14662 8425 14714
rect 8449 14662 8495 14714
rect 8495 14662 8505 14714
rect 8529 14662 8559 14714
rect 8559 14662 8585 14714
rect 8289 14660 8345 14662
rect 8369 14660 8425 14662
rect 8449 14660 8505 14662
rect 8529 14660 8585 14662
rect 8850 15408 8906 15464
rect 8289 13626 8345 13628
rect 8369 13626 8425 13628
rect 8449 13626 8505 13628
rect 8529 13626 8585 13628
rect 8289 13574 8315 13626
rect 8315 13574 8345 13626
rect 8369 13574 8379 13626
rect 8379 13574 8425 13626
rect 8449 13574 8495 13626
rect 8495 13574 8505 13626
rect 8529 13574 8559 13626
rect 8559 13574 8585 13626
rect 8289 13572 8345 13574
rect 8369 13572 8425 13574
rect 8449 13572 8505 13574
rect 8529 13572 8585 13574
rect 8289 12538 8345 12540
rect 8369 12538 8425 12540
rect 8449 12538 8505 12540
rect 8529 12538 8585 12540
rect 8289 12486 8315 12538
rect 8315 12486 8345 12538
rect 8369 12486 8379 12538
rect 8379 12486 8425 12538
rect 8449 12486 8495 12538
rect 8495 12486 8505 12538
rect 8529 12486 8559 12538
rect 8559 12486 8585 12538
rect 8289 12484 8345 12486
rect 8369 12484 8425 12486
rect 8449 12484 8505 12486
rect 8529 12484 8585 12486
rect 8289 11450 8345 11452
rect 8369 11450 8425 11452
rect 8449 11450 8505 11452
rect 8529 11450 8585 11452
rect 8289 11398 8315 11450
rect 8315 11398 8345 11450
rect 8369 11398 8379 11450
rect 8379 11398 8425 11450
rect 8449 11398 8495 11450
rect 8495 11398 8505 11450
rect 8529 11398 8559 11450
rect 8559 11398 8585 11450
rect 8289 11396 8345 11398
rect 8369 11396 8425 11398
rect 8449 11396 8505 11398
rect 8529 11396 8585 11398
rect 8289 10362 8345 10364
rect 8369 10362 8425 10364
rect 8449 10362 8505 10364
rect 8529 10362 8585 10364
rect 8289 10310 8315 10362
rect 8315 10310 8345 10362
rect 8369 10310 8379 10362
rect 8379 10310 8425 10362
rect 8449 10310 8495 10362
rect 8495 10310 8505 10362
rect 8529 10310 8559 10362
rect 8559 10310 8585 10362
rect 8289 10308 8345 10310
rect 8369 10308 8425 10310
rect 8449 10308 8505 10310
rect 8529 10308 8585 10310
rect 8289 9274 8345 9276
rect 8369 9274 8425 9276
rect 8449 9274 8505 9276
rect 8529 9274 8585 9276
rect 8289 9222 8315 9274
rect 8315 9222 8345 9274
rect 8369 9222 8379 9274
rect 8379 9222 8425 9274
rect 8449 9222 8495 9274
rect 8495 9222 8505 9274
rect 8529 9222 8559 9274
rect 8559 9222 8585 9274
rect 8289 9220 8345 9222
rect 8369 9220 8425 9222
rect 8449 9220 8505 9222
rect 8529 9220 8585 9222
rect 8289 8186 8345 8188
rect 8369 8186 8425 8188
rect 8449 8186 8505 8188
rect 8529 8186 8585 8188
rect 8289 8134 8315 8186
rect 8315 8134 8345 8186
rect 8369 8134 8379 8186
rect 8379 8134 8425 8186
rect 8449 8134 8495 8186
rect 8495 8134 8505 8186
rect 8529 8134 8559 8186
rect 8559 8134 8585 8186
rect 8289 8132 8345 8134
rect 8369 8132 8425 8134
rect 8449 8132 8505 8134
rect 8529 8132 8585 8134
rect 8666 7928 8722 7984
rect 8289 7098 8345 7100
rect 8369 7098 8425 7100
rect 8449 7098 8505 7100
rect 8529 7098 8585 7100
rect 8289 7046 8315 7098
rect 8315 7046 8345 7098
rect 8369 7046 8379 7098
rect 8379 7046 8425 7098
rect 8449 7046 8495 7098
rect 8495 7046 8505 7098
rect 8529 7046 8559 7098
rect 8559 7046 8585 7098
rect 8289 7044 8345 7046
rect 8369 7044 8425 7046
rect 8449 7044 8505 7046
rect 8529 7044 8585 7046
rect 7194 3440 7250 3496
rect 7838 4936 7894 4992
rect 8289 6010 8345 6012
rect 8369 6010 8425 6012
rect 8449 6010 8505 6012
rect 8529 6010 8585 6012
rect 8289 5958 8315 6010
rect 8315 5958 8345 6010
rect 8369 5958 8379 6010
rect 8379 5958 8425 6010
rect 8449 5958 8495 6010
rect 8495 5958 8505 6010
rect 8529 5958 8559 6010
rect 8559 5958 8585 6010
rect 8289 5956 8345 5958
rect 8369 5956 8425 5958
rect 8449 5956 8505 5958
rect 8529 5956 8585 5958
rect 8206 5752 8262 5808
rect 8289 4922 8345 4924
rect 8369 4922 8425 4924
rect 8449 4922 8505 4924
rect 8529 4922 8585 4924
rect 8289 4870 8315 4922
rect 8315 4870 8345 4922
rect 8369 4870 8379 4922
rect 8379 4870 8425 4922
rect 8449 4870 8495 4922
rect 8495 4870 8505 4922
rect 8529 4870 8559 4922
rect 8559 4870 8585 4922
rect 8289 4868 8345 4870
rect 8369 4868 8425 4870
rect 8449 4868 8505 4870
rect 8529 4868 8585 4870
rect 9310 16768 9366 16824
rect 9402 15272 9458 15328
rect 9586 14456 9642 14512
rect 9862 14320 9918 14376
rect 9218 12144 9274 12200
rect 8758 4664 8814 4720
rect 8114 3984 8170 4040
rect 8574 3984 8630 4040
rect 8289 3834 8345 3836
rect 8369 3834 8425 3836
rect 8449 3834 8505 3836
rect 8529 3834 8585 3836
rect 8289 3782 8315 3834
rect 8315 3782 8345 3834
rect 8369 3782 8379 3834
rect 8379 3782 8425 3834
rect 8449 3782 8495 3834
rect 8495 3782 8505 3834
rect 8529 3782 8559 3834
rect 8559 3782 8585 3834
rect 8289 3780 8345 3782
rect 8369 3780 8425 3782
rect 8449 3780 8505 3782
rect 8529 3780 8585 3782
rect 9126 2896 9182 2952
rect 8289 2746 8345 2748
rect 8369 2746 8425 2748
rect 8449 2746 8505 2748
rect 8529 2746 8585 2748
rect 8289 2694 8315 2746
rect 8315 2694 8345 2746
rect 8369 2694 8379 2746
rect 8379 2694 8425 2746
rect 8449 2694 8495 2746
rect 8495 2694 8505 2746
rect 8529 2694 8559 2746
rect 8559 2694 8585 2746
rect 8289 2692 8345 2694
rect 8369 2692 8425 2694
rect 8449 2692 8505 2694
rect 8529 2692 8585 2694
rect 10506 16496 10562 16552
rect 9862 8880 9918 8936
rect 9770 4256 9826 4312
rect 10598 11600 10654 11656
rect 10782 16904 10838 16960
rect 10598 4528 10654 4584
rect 10874 5616 10930 5672
rect 11956 19610 12012 19612
rect 12036 19610 12092 19612
rect 12116 19610 12172 19612
rect 12196 19610 12252 19612
rect 11956 19558 11982 19610
rect 11982 19558 12012 19610
rect 12036 19558 12046 19610
rect 12046 19558 12092 19610
rect 12116 19558 12162 19610
rect 12162 19558 12172 19610
rect 12196 19558 12226 19610
rect 12226 19558 12252 19610
rect 11956 19556 12012 19558
rect 12036 19556 12092 19558
rect 12116 19556 12172 19558
rect 12196 19556 12252 19558
rect 11426 15816 11482 15872
rect 11334 14728 11390 14784
rect 11150 9560 11206 9616
rect 11956 18522 12012 18524
rect 12036 18522 12092 18524
rect 12116 18522 12172 18524
rect 12196 18522 12252 18524
rect 11956 18470 11982 18522
rect 11982 18470 12012 18522
rect 12036 18470 12046 18522
rect 12046 18470 12092 18522
rect 12116 18470 12162 18522
rect 12162 18470 12172 18522
rect 12196 18470 12226 18522
rect 12226 18470 12252 18522
rect 11956 18468 12012 18470
rect 12036 18468 12092 18470
rect 12116 18468 12172 18470
rect 12196 18468 12252 18470
rect 11702 17040 11758 17096
rect 11956 17434 12012 17436
rect 12036 17434 12092 17436
rect 12116 17434 12172 17436
rect 12196 17434 12252 17436
rect 11956 17382 11982 17434
rect 11982 17382 12012 17434
rect 12036 17382 12046 17434
rect 12046 17382 12092 17434
rect 12116 17382 12162 17434
rect 12162 17382 12172 17434
rect 12196 17382 12226 17434
rect 12226 17382 12252 17434
rect 11956 17380 12012 17382
rect 12036 17380 12092 17382
rect 12116 17380 12172 17382
rect 12196 17380 12252 17382
rect 11956 16346 12012 16348
rect 12036 16346 12092 16348
rect 12116 16346 12172 16348
rect 12196 16346 12252 16348
rect 11956 16294 11982 16346
rect 11982 16294 12012 16346
rect 12036 16294 12046 16346
rect 12046 16294 12092 16346
rect 12116 16294 12162 16346
rect 12162 16294 12172 16346
rect 12196 16294 12226 16346
rect 12226 16294 12252 16346
rect 11956 16292 12012 16294
rect 12036 16292 12092 16294
rect 12116 16292 12172 16294
rect 12196 16292 12252 16294
rect 11956 15258 12012 15260
rect 12036 15258 12092 15260
rect 12116 15258 12172 15260
rect 12196 15258 12252 15260
rect 11956 15206 11982 15258
rect 11982 15206 12012 15258
rect 12036 15206 12046 15258
rect 12046 15206 12092 15258
rect 12116 15206 12162 15258
rect 12162 15206 12172 15258
rect 12196 15206 12226 15258
rect 12226 15206 12252 15258
rect 11956 15204 12012 15206
rect 12036 15204 12092 15206
rect 12116 15204 12172 15206
rect 12196 15204 12252 15206
rect 11956 14170 12012 14172
rect 12036 14170 12092 14172
rect 12116 14170 12172 14172
rect 12196 14170 12252 14172
rect 11956 14118 11982 14170
rect 11982 14118 12012 14170
rect 12036 14118 12046 14170
rect 12046 14118 12092 14170
rect 12116 14118 12162 14170
rect 12162 14118 12172 14170
rect 12196 14118 12226 14170
rect 12226 14118 12252 14170
rect 11956 14116 12012 14118
rect 12036 14116 12092 14118
rect 12116 14116 12172 14118
rect 12196 14116 12252 14118
rect 12070 13912 12126 13968
rect 11956 13082 12012 13084
rect 12036 13082 12092 13084
rect 12116 13082 12172 13084
rect 12196 13082 12252 13084
rect 11956 13030 11982 13082
rect 11982 13030 12012 13082
rect 12036 13030 12046 13082
rect 12046 13030 12092 13082
rect 12116 13030 12162 13082
rect 12162 13030 12172 13082
rect 12196 13030 12226 13082
rect 12226 13030 12252 13082
rect 11956 13028 12012 13030
rect 12036 13028 12092 13030
rect 12116 13028 12172 13030
rect 12196 13028 12252 13030
rect 11956 11994 12012 11996
rect 12036 11994 12092 11996
rect 12116 11994 12172 11996
rect 12196 11994 12252 11996
rect 11956 11942 11982 11994
rect 11982 11942 12012 11994
rect 12036 11942 12046 11994
rect 12046 11942 12092 11994
rect 12116 11942 12162 11994
rect 12162 11942 12172 11994
rect 12196 11942 12226 11994
rect 12226 11942 12252 11994
rect 11956 11940 12012 11942
rect 12036 11940 12092 11942
rect 12116 11940 12172 11942
rect 12196 11940 12252 11942
rect 11956 10906 12012 10908
rect 12036 10906 12092 10908
rect 12116 10906 12172 10908
rect 12196 10906 12252 10908
rect 11956 10854 11982 10906
rect 11982 10854 12012 10906
rect 12036 10854 12046 10906
rect 12046 10854 12092 10906
rect 12116 10854 12162 10906
rect 12162 10854 12172 10906
rect 12196 10854 12226 10906
rect 12226 10854 12252 10906
rect 11956 10852 12012 10854
rect 12036 10852 12092 10854
rect 12116 10852 12172 10854
rect 12196 10852 12252 10854
rect 11956 9818 12012 9820
rect 12036 9818 12092 9820
rect 12116 9818 12172 9820
rect 12196 9818 12252 9820
rect 11956 9766 11982 9818
rect 11982 9766 12012 9818
rect 12036 9766 12046 9818
rect 12046 9766 12092 9818
rect 12116 9766 12162 9818
rect 12162 9766 12172 9818
rect 12196 9766 12226 9818
rect 12226 9766 12252 9818
rect 11956 9764 12012 9766
rect 12036 9764 12092 9766
rect 12116 9764 12172 9766
rect 12196 9764 12252 9766
rect 11956 8730 12012 8732
rect 12036 8730 12092 8732
rect 12116 8730 12172 8732
rect 12196 8730 12252 8732
rect 11956 8678 11982 8730
rect 11982 8678 12012 8730
rect 12036 8678 12046 8730
rect 12046 8678 12092 8730
rect 12116 8678 12162 8730
rect 12162 8678 12172 8730
rect 12196 8678 12226 8730
rect 12226 8678 12252 8730
rect 11956 8676 12012 8678
rect 12036 8676 12092 8678
rect 12116 8676 12172 8678
rect 12196 8676 12252 8678
rect 11956 7642 12012 7644
rect 12036 7642 12092 7644
rect 12116 7642 12172 7644
rect 12196 7642 12252 7644
rect 11956 7590 11982 7642
rect 11982 7590 12012 7642
rect 12036 7590 12046 7642
rect 12046 7590 12092 7642
rect 12116 7590 12162 7642
rect 12162 7590 12172 7642
rect 12196 7590 12226 7642
rect 12226 7590 12252 7642
rect 11956 7588 12012 7590
rect 12036 7588 12092 7590
rect 12116 7588 12172 7590
rect 12196 7588 12252 7590
rect 11956 6554 12012 6556
rect 12036 6554 12092 6556
rect 12116 6554 12172 6556
rect 12196 6554 12252 6556
rect 11956 6502 11982 6554
rect 11982 6502 12012 6554
rect 12036 6502 12046 6554
rect 12046 6502 12092 6554
rect 12116 6502 12162 6554
rect 12162 6502 12172 6554
rect 12196 6502 12226 6554
rect 12226 6502 12252 6554
rect 11956 6500 12012 6502
rect 12036 6500 12092 6502
rect 12116 6500 12172 6502
rect 12196 6500 12252 6502
rect 11956 5466 12012 5468
rect 12036 5466 12092 5468
rect 12116 5466 12172 5468
rect 12196 5466 12252 5468
rect 11956 5414 11982 5466
rect 11982 5414 12012 5466
rect 12036 5414 12046 5466
rect 12046 5414 12092 5466
rect 12116 5414 12162 5466
rect 12162 5414 12172 5466
rect 12196 5414 12226 5466
rect 12226 5414 12252 5466
rect 11956 5412 12012 5414
rect 12036 5412 12092 5414
rect 12116 5412 12172 5414
rect 12196 5412 12252 5414
rect 11702 5072 11758 5128
rect 12622 14184 12678 14240
rect 12806 10104 12862 10160
rect 12990 10512 13046 10568
rect 11956 4378 12012 4380
rect 12036 4378 12092 4380
rect 12116 4378 12172 4380
rect 12196 4378 12252 4380
rect 11956 4326 11982 4378
rect 11982 4326 12012 4378
rect 12036 4326 12046 4378
rect 12046 4326 12092 4378
rect 12116 4326 12162 4378
rect 12162 4326 12172 4378
rect 12196 4326 12226 4378
rect 12226 4326 12252 4378
rect 11956 4324 12012 4326
rect 12036 4324 12092 4326
rect 12116 4324 12172 4326
rect 12196 4324 12252 4326
rect 12622 4528 12678 4584
rect 11956 3290 12012 3292
rect 12036 3290 12092 3292
rect 12116 3290 12172 3292
rect 12196 3290 12252 3292
rect 11956 3238 11982 3290
rect 11982 3238 12012 3290
rect 12036 3238 12046 3290
rect 12046 3238 12092 3290
rect 12116 3238 12162 3290
rect 12162 3238 12172 3290
rect 12196 3238 12226 3290
rect 12226 3238 12252 3290
rect 11956 3236 12012 3238
rect 12036 3236 12092 3238
rect 12116 3236 12172 3238
rect 12196 3236 12252 3238
rect 11242 2352 11298 2408
rect 11956 2202 12012 2204
rect 12036 2202 12092 2204
rect 12116 2202 12172 2204
rect 12196 2202 12252 2204
rect 11956 2150 11982 2202
rect 11982 2150 12012 2202
rect 12036 2150 12046 2202
rect 12046 2150 12092 2202
rect 12116 2150 12162 2202
rect 12162 2150 12172 2202
rect 12196 2150 12226 2202
rect 12226 2150 12252 2202
rect 11956 2148 12012 2150
rect 12036 2148 12092 2150
rect 12116 2148 12172 2150
rect 12196 2148 12252 2150
rect 13266 14184 13322 14240
rect 13542 14864 13598 14920
rect 13450 14320 13506 14376
rect 13358 10784 13414 10840
rect 13818 17176 13874 17232
rect 13726 14864 13782 14920
rect 13818 13232 13874 13288
rect 14094 13368 14150 13424
rect 13726 10104 13782 10160
rect 13358 2488 13414 2544
rect 14646 17584 14702 17640
rect 15622 19066 15678 19068
rect 15702 19066 15758 19068
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15622 19014 15648 19066
rect 15648 19014 15678 19066
rect 15702 19014 15712 19066
rect 15712 19014 15758 19066
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15918 19066
rect 15622 19012 15678 19014
rect 15702 19012 15758 19014
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 15622 17978 15678 17980
rect 15702 17978 15758 17980
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15622 17926 15648 17978
rect 15648 17926 15678 17978
rect 15702 17926 15712 17978
rect 15712 17926 15758 17978
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15918 17978
rect 15622 17924 15678 17926
rect 15702 17924 15758 17926
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 16026 17720 16082 17776
rect 15622 16890 15678 16892
rect 15702 16890 15758 16892
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15622 16838 15648 16890
rect 15648 16838 15678 16890
rect 15702 16838 15712 16890
rect 15712 16838 15758 16890
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15918 16890
rect 15622 16836 15678 16838
rect 15702 16836 15758 16838
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15622 15802 15678 15804
rect 15702 15802 15758 15804
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15622 15750 15648 15802
rect 15648 15750 15678 15802
rect 15702 15750 15712 15802
rect 15712 15750 15758 15802
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15918 15802
rect 15622 15748 15678 15750
rect 15702 15748 15758 15750
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15622 14714 15678 14716
rect 15702 14714 15758 14716
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15622 14662 15648 14714
rect 15648 14662 15678 14714
rect 15702 14662 15712 14714
rect 15712 14662 15758 14714
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15918 14714
rect 15622 14660 15678 14662
rect 15702 14660 15758 14662
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15290 10104 15346 10160
rect 15622 13626 15678 13628
rect 15702 13626 15758 13628
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15622 13574 15648 13626
rect 15648 13574 15678 13626
rect 15702 13574 15712 13626
rect 15712 13574 15758 13626
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15918 13626
rect 15622 13572 15678 13574
rect 15702 13572 15758 13574
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15622 12538 15678 12540
rect 15702 12538 15758 12540
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15622 12486 15648 12538
rect 15648 12486 15678 12538
rect 15702 12486 15712 12538
rect 15712 12486 15758 12538
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15918 12538
rect 15622 12484 15678 12486
rect 15702 12484 15758 12486
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15622 11450 15678 11452
rect 15702 11450 15758 11452
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15622 11398 15648 11450
rect 15648 11398 15678 11450
rect 15702 11398 15712 11450
rect 15712 11398 15758 11450
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15918 11450
rect 15622 11396 15678 11398
rect 15702 11396 15758 11398
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15622 10362 15678 10364
rect 15702 10362 15758 10364
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15622 10310 15648 10362
rect 15648 10310 15678 10362
rect 15702 10310 15712 10362
rect 15712 10310 15758 10362
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15918 10362
rect 15622 10308 15678 10310
rect 15702 10308 15758 10310
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 15750 9424 15806 9480
rect 15622 9274 15678 9276
rect 15702 9274 15758 9276
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15622 9222 15648 9274
rect 15648 9222 15678 9274
rect 15702 9222 15712 9274
rect 15712 9222 15758 9274
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15918 9274
rect 15622 9220 15678 9222
rect 15702 9220 15758 9222
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 16118 11328 16174 11384
rect 15622 8186 15678 8188
rect 15702 8186 15758 8188
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15622 8134 15648 8186
rect 15648 8134 15678 8186
rect 15702 8134 15712 8186
rect 15712 8134 15758 8186
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15918 8186
rect 15622 8132 15678 8134
rect 15702 8132 15758 8134
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15622 7098 15678 7100
rect 15702 7098 15758 7100
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15622 7046 15648 7098
rect 15648 7046 15678 7098
rect 15702 7046 15712 7098
rect 15712 7046 15758 7098
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15918 7098
rect 15622 7044 15678 7046
rect 15702 7044 15758 7046
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 16026 6296 16082 6352
rect 15198 5208 15254 5264
rect 14830 4664 14886 4720
rect 15622 6010 15678 6012
rect 15702 6010 15758 6012
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15622 5958 15648 6010
rect 15648 5958 15678 6010
rect 15702 5958 15712 6010
rect 15712 5958 15758 6010
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15918 6010
rect 15622 5956 15678 5958
rect 15702 5956 15758 5958
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 17498 18672 17554 18728
rect 16762 17992 16818 18048
rect 16670 8880 16726 8936
rect 15622 4922 15678 4924
rect 15702 4922 15758 4924
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15622 4870 15648 4922
rect 15648 4870 15678 4922
rect 15702 4870 15712 4922
rect 15712 4870 15758 4922
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15918 4922
rect 15622 4868 15678 4870
rect 15702 4868 15758 4870
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15622 3834 15678 3836
rect 15702 3834 15758 3836
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15622 3782 15648 3834
rect 15648 3782 15678 3834
rect 15702 3782 15712 3834
rect 15712 3782 15758 3834
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15918 3834
rect 15622 3780 15678 3782
rect 15702 3780 15758 3782
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 15622 2746 15678 2748
rect 15702 2746 15758 2748
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15622 2694 15648 2746
rect 15648 2694 15678 2746
rect 15702 2694 15712 2746
rect 15712 2694 15758 2746
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15918 2746
rect 15622 2692 15678 2694
rect 15702 2692 15758 2694
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 16026 3032 16082 3088
rect 17406 15952 17462 16008
rect 18510 17992 18566 18048
rect 18694 17584 18750 17640
rect 17406 13640 17462 13696
rect 17130 4528 17186 4584
rect 17774 15408 17830 15464
rect 17682 13504 17738 13560
rect 18142 13776 18198 13832
rect 17774 4120 17830 4176
rect 19614 20440 19670 20496
rect 19289 19610 19345 19612
rect 19369 19610 19425 19612
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19289 19558 19315 19610
rect 19315 19558 19345 19610
rect 19369 19558 19379 19610
rect 19379 19558 19425 19610
rect 19449 19558 19495 19610
rect 19495 19558 19505 19610
rect 19529 19558 19559 19610
rect 19559 19558 19585 19610
rect 19289 19556 19345 19558
rect 19369 19556 19425 19558
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19289 18522 19345 18524
rect 19369 18522 19425 18524
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19289 18470 19315 18522
rect 19315 18470 19345 18522
rect 19369 18470 19379 18522
rect 19379 18470 19425 18522
rect 19449 18470 19495 18522
rect 19495 18470 19505 18522
rect 19529 18470 19559 18522
rect 19559 18470 19585 18522
rect 19289 18468 19345 18470
rect 19369 18468 19425 18470
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19289 17434 19345 17436
rect 19369 17434 19425 17436
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19289 17382 19315 17434
rect 19315 17382 19345 17434
rect 19369 17382 19379 17434
rect 19379 17382 19425 17434
rect 19449 17382 19495 17434
rect 19495 17382 19505 17434
rect 19529 17382 19559 17434
rect 19559 17382 19585 17434
rect 19289 17380 19345 17382
rect 19369 17380 19425 17382
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19522 16904 19578 16960
rect 19289 16346 19345 16348
rect 19369 16346 19425 16348
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19289 16294 19315 16346
rect 19315 16294 19345 16346
rect 19369 16294 19379 16346
rect 19379 16294 19425 16346
rect 19449 16294 19495 16346
rect 19495 16294 19505 16346
rect 19529 16294 19559 16346
rect 19559 16294 19585 16346
rect 19289 16292 19345 16294
rect 19369 16292 19425 16294
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19289 15258 19345 15260
rect 19369 15258 19425 15260
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19289 15206 19315 15258
rect 19315 15206 19345 15258
rect 19369 15206 19379 15258
rect 19379 15206 19425 15258
rect 19449 15206 19495 15258
rect 19495 15206 19505 15258
rect 19529 15206 19559 15258
rect 19559 15206 19585 15258
rect 19289 15204 19345 15206
rect 19369 15204 19425 15206
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19154 15000 19210 15056
rect 19154 14456 19210 14512
rect 19289 14170 19345 14172
rect 19369 14170 19425 14172
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19289 14118 19315 14170
rect 19315 14118 19345 14170
rect 19369 14118 19379 14170
rect 19379 14118 19425 14170
rect 19449 14118 19495 14170
rect 19495 14118 19505 14170
rect 19529 14118 19559 14170
rect 19559 14118 19585 14170
rect 19289 14116 19345 14118
rect 19369 14116 19425 14118
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19289 13082 19345 13084
rect 19369 13082 19425 13084
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19289 13030 19315 13082
rect 19315 13030 19345 13082
rect 19369 13030 19379 13082
rect 19379 13030 19425 13082
rect 19449 13030 19495 13082
rect 19495 13030 19505 13082
rect 19529 13030 19559 13082
rect 19559 13030 19585 13082
rect 19289 13028 19345 13030
rect 19369 13028 19425 13030
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19289 11994 19345 11996
rect 19369 11994 19425 11996
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19289 11942 19315 11994
rect 19315 11942 19345 11994
rect 19369 11942 19379 11994
rect 19379 11942 19425 11994
rect 19449 11942 19495 11994
rect 19495 11942 19505 11994
rect 19529 11942 19559 11994
rect 19559 11942 19585 11994
rect 19289 11940 19345 11942
rect 19369 11940 19425 11942
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19289 10906 19345 10908
rect 19369 10906 19425 10908
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19289 10854 19315 10906
rect 19315 10854 19345 10906
rect 19369 10854 19379 10906
rect 19379 10854 19425 10906
rect 19449 10854 19495 10906
rect 19495 10854 19505 10906
rect 19529 10854 19559 10906
rect 19559 10854 19585 10906
rect 19289 10852 19345 10854
rect 19369 10852 19425 10854
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19289 9818 19345 9820
rect 19369 9818 19425 9820
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19289 9766 19315 9818
rect 19315 9766 19345 9818
rect 19369 9766 19379 9818
rect 19379 9766 19425 9818
rect 19449 9766 19495 9818
rect 19495 9766 19505 9818
rect 19529 9766 19559 9818
rect 19559 9766 19585 9818
rect 19289 9764 19345 9766
rect 19369 9764 19425 9766
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19289 8730 19345 8732
rect 19369 8730 19425 8732
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19289 8678 19315 8730
rect 19315 8678 19345 8730
rect 19369 8678 19379 8730
rect 19379 8678 19425 8730
rect 19449 8678 19495 8730
rect 19495 8678 19505 8730
rect 19529 8678 19559 8730
rect 19559 8678 19585 8730
rect 19289 8676 19345 8678
rect 19369 8676 19425 8678
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 21546 15544 21602 15600
rect 20074 9560 20130 9616
rect 19289 7642 19345 7644
rect 19369 7642 19425 7644
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19289 7590 19315 7642
rect 19315 7590 19345 7642
rect 19369 7590 19379 7642
rect 19379 7590 19425 7642
rect 19449 7590 19495 7642
rect 19495 7590 19505 7642
rect 19529 7590 19559 7642
rect 19559 7590 19585 7642
rect 19289 7588 19345 7590
rect 19369 7588 19425 7590
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19289 6554 19345 6556
rect 19369 6554 19425 6556
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19289 6502 19315 6554
rect 19315 6502 19345 6554
rect 19369 6502 19379 6554
rect 19379 6502 19425 6554
rect 19449 6502 19495 6554
rect 19495 6502 19505 6554
rect 19529 6502 19559 6554
rect 19559 6502 19585 6554
rect 19289 6500 19345 6502
rect 19369 6500 19425 6502
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19289 5466 19345 5468
rect 19369 5466 19425 5468
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19289 5414 19315 5466
rect 19315 5414 19345 5466
rect 19369 5414 19379 5466
rect 19379 5414 19425 5466
rect 19449 5414 19495 5466
rect 19495 5414 19505 5466
rect 19529 5414 19559 5466
rect 19559 5414 19585 5466
rect 19289 5412 19345 5414
rect 19369 5412 19425 5414
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 19154 4528 19210 4584
rect 19430 4528 19486 4584
rect 19289 4378 19345 4380
rect 19369 4378 19425 4380
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19289 4326 19315 4378
rect 19315 4326 19345 4378
rect 19369 4326 19379 4378
rect 19379 4326 19425 4378
rect 19449 4326 19495 4378
rect 19495 4326 19505 4378
rect 19529 4326 19559 4378
rect 19559 4326 19585 4378
rect 19289 4324 19345 4326
rect 19369 4324 19425 4326
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 18878 3440 18934 3496
rect 19289 3290 19345 3292
rect 19369 3290 19425 3292
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19289 3238 19315 3290
rect 19315 3238 19345 3290
rect 19369 3238 19379 3290
rect 19379 3238 19425 3290
rect 19449 3238 19495 3290
rect 19495 3238 19505 3290
rect 19529 3238 19559 3290
rect 19559 3238 19585 3290
rect 19289 3236 19345 3238
rect 19369 3236 19425 3238
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19289 2202 19345 2204
rect 19369 2202 19425 2204
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19289 2150 19315 2202
rect 19315 2150 19345 2202
rect 19369 2150 19379 2202
rect 19379 2150 19425 2202
rect 19449 2150 19495 2202
rect 19495 2150 19505 2202
rect 19529 2150 19559 2202
rect 19559 2150 19585 2202
rect 19289 2148 19345 2150
rect 19369 2148 19425 2150
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 17958 1264 18014 1320
rect 20350 1400 20406 1456
rect 21546 8200 21602 8256
rect 21546 6296 21602 6352
<< metal3 >>
rect 0 20952 480 21072
rect 21520 20952 22000 21072
rect 62 20498 122 20952
rect 1485 20498 1551 20501
rect 62 20496 1551 20498
rect 62 20440 1490 20496
rect 1546 20440 1551 20496
rect 62 20438 1551 20440
rect 1485 20435 1551 20438
rect 19609 20498 19675 20501
rect 21590 20498 21650 20952
rect 19609 20496 21650 20498
rect 19609 20440 19614 20496
rect 19670 20440 21650 20496
rect 19609 20438 21650 20440
rect 19609 20435 19675 20438
rect 4610 19616 4930 19617
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4930 19616
rect 4610 19551 4930 19552
rect 11944 19616 12264 19617
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 19551 12264 19552
rect 19277 19616 19597 19617
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 19551 19597 19552
rect 0 19184 480 19304
rect 21520 19184 22000 19304
rect 62 18730 122 19184
rect 8277 19072 8597 19073
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 19007 8597 19008
rect 15610 19072 15930 19073
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 19007 15930 19008
rect 1301 18730 1367 18733
rect 62 18728 1367 18730
rect 62 18672 1306 18728
rect 1362 18672 1367 18728
rect 62 18670 1367 18672
rect 1301 18667 1367 18670
rect 17493 18730 17559 18733
rect 21590 18730 21650 19184
rect 17493 18728 21650 18730
rect 17493 18672 17498 18728
rect 17554 18672 21650 18728
rect 17493 18670 21650 18672
rect 17493 18667 17559 18670
rect 4610 18528 4930 18529
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4930 18528
rect 4610 18463 4930 18464
rect 11944 18528 12264 18529
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 18463 12264 18464
rect 19277 18528 19597 18529
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 18463 19597 18464
rect 16757 18052 16823 18053
rect 16757 18050 16804 18052
rect 16676 18048 16804 18050
rect 16868 18050 16874 18052
rect 18505 18050 18571 18053
rect 16868 18048 18571 18050
rect 16676 17992 16762 18048
rect 16868 17992 18510 18048
rect 18566 17992 18571 18048
rect 16676 17990 16804 17992
rect 16757 17988 16804 17990
rect 16868 17990 18571 17992
rect 16868 17988 16874 17990
rect 16757 17987 16823 17988
rect 18505 17987 18571 17990
rect 8277 17984 8597 17985
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 17919 8597 17920
rect 15610 17984 15930 17985
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 17919 15930 17920
rect 6361 17778 6427 17781
rect 16021 17778 16087 17781
rect 6361 17776 16087 17778
rect 6361 17720 6366 17776
rect 6422 17720 16026 17776
rect 16082 17720 16087 17776
rect 6361 17718 16087 17720
rect 6361 17715 6427 17718
rect 16021 17715 16087 17718
rect 4521 17642 4587 17645
rect 6637 17642 6703 17645
rect 14641 17642 14707 17645
rect 18689 17642 18755 17645
rect 4521 17640 18755 17642
rect 4521 17584 4526 17640
rect 4582 17584 6642 17640
rect 6698 17584 14646 17640
rect 14702 17584 18694 17640
rect 18750 17584 18755 17640
rect 4521 17582 18755 17584
rect 4521 17579 4587 17582
rect 6637 17579 6703 17582
rect 14641 17579 14707 17582
rect 18689 17579 18755 17582
rect 4610 17440 4930 17441
rect 0 17368 480 17400
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4930 17440
rect 4610 17375 4930 17376
rect 11944 17440 12264 17441
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 17375 12264 17376
rect 19277 17440 19597 17441
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 17375 19597 17376
rect 0 17312 110 17368
rect 166 17312 480 17368
rect 0 17280 480 17312
rect 21520 17280 22000 17400
rect 13486 17172 13492 17236
rect 13556 17234 13562 17236
rect 13813 17234 13879 17237
rect 13556 17232 13879 17234
rect 13556 17176 13818 17232
rect 13874 17176 13879 17232
rect 13556 17174 13879 17176
rect 13556 17172 13562 17174
rect 13813 17171 13879 17174
rect 749 17098 815 17101
rect 11697 17098 11763 17101
rect 749 17096 11763 17098
rect 749 17040 754 17096
rect 810 17040 11702 17096
rect 11758 17040 11763 17096
rect 749 17038 11763 17040
rect 749 17035 815 17038
rect 11697 17035 11763 17038
rect 7598 16900 7604 16964
rect 7668 16962 7674 16964
rect 7741 16962 7807 16965
rect 7668 16960 7807 16962
rect 7668 16904 7746 16960
rect 7802 16904 7807 16960
rect 7668 16902 7807 16904
rect 7668 16900 7674 16902
rect 7741 16899 7807 16902
rect 8753 16962 8819 16965
rect 9990 16962 9996 16964
rect 8753 16960 9996 16962
rect 8753 16904 8758 16960
rect 8814 16904 9996 16960
rect 8753 16902 9996 16904
rect 8753 16899 8819 16902
rect 9990 16900 9996 16902
rect 10060 16962 10066 16964
rect 10777 16962 10843 16965
rect 10060 16960 10843 16962
rect 10060 16904 10782 16960
rect 10838 16904 10843 16960
rect 10060 16902 10843 16904
rect 10060 16900 10066 16902
rect 10777 16899 10843 16902
rect 19517 16962 19583 16965
rect 21590 16962 21650 17280
rect 19517 16960 21650 16962
rect 19517 16904 19522 16960
rect 19578 16904 21650 16960
rect 19517 16902 21650 16904
rect 19517 16899 19583 16902
rect 8277 16896 8597 16897
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 16831 8597 16832
rect 15610 16896 15930 16897
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 16831 15930 16832
rect 9305 16826 9371 16829
rect 9438 16826 9444 16828
rect 9305 16824 9444 16826
rect 9305 16768 9310 16824
rect 9366 16768 9444 16824
rect 9305 16766 9444 16768
rect 9305 16763 9371 16766
rect 9438 16764 9444 16766
rect 9508 16764 9514 16828
rect 9070 16492 9076 16556
rect 9140 16554 9146 16556
rect 10501 16554 10567 16557
rect 9140 16552 10567 16554
rect 9140 16496 10506 16552
rect 10562 16496 10567 16552
rect 9140 16494 10567 16496
rect 9140 16492 9146 16494
rect 10501 16491 10567 16494
rect 4610 16352 4930 16353
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4930 16352
rect 4610 16287 4930 16288
rect 11944 16352 12264 16353
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 16287 12264 16288
rect 19277 16352 19597 16353
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 16287 19597 16288
rect 8702 16220 8708 16284
rect 8772 16282 8778 16284
rect 8845 16282 8911 16285
rect 8772 16280 8911 16282
rect 8772 16224 8850 16280
rect 8906 16224 8911 16280
rect 8772 16222 8911 16224
rect 8772 16220 8778 16222
rect 8845 16219 8911 16222
rect 6637 16012 6703 16013
rect 6637 16010 6684 16012
rect 6556 16008 6684 16010
rect 6748 16010 6754 16012
rect 17401 16010 17467 16013
rect 6748 16008 17467 16010
rect 6556 15952 6642 16008
rect 6748 15952 17406 16008
rect 17462 15952 17467 16008
rect 6556 15950 6684 15952
rect 6637 15948 6684 15950
rect 6748 15950 17467 15952
rect 6748 15948 6754 15950
rect 6637 15947 6703 15948
rect 17401 15947 17467 15950
rect 11278 15812 11284 15876
rect 11348 15874 11354 15876
rect 11421 15874 11487 15877
rect 11348 15872 11487 15874
rect 11348 15816 11426 15872
rect 11482 15816 11487 15872
rect 11348 15814 11487 15816
rect 11348 15812 11354 15814
rect 11421 15811 11487 15814
rect 8277 15808 8597 15809
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 15743 8597 15744
rect 15610 15808 15930 15809
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 15743 15930 15744
rect 0 15600 480 15632
rect 21520 15602 22000 15632
rect 0 15544 110 15600
rect 166 15544 480 15600
rect 0 15512 480 15544
rect 21460 15600 22000 15602
rect 21460 15544 21546 15600
rect 21602 15544 22000 15600
rect 21460 15542 22000 15544
rect 21520 15512 22000 15542
rect 8845 15466 8911 15469
rect 17769 15466 17835 15469
rect 8845 15464 17835 15466
rect 8845 15408 8850 15464
rect 8906 15408 17774 15464
rect 17830 15408 17835 15464
rect 8845 15406 17835 15408
rect 8845 15403 8911 15406
rect 17769 15403 17835 15406
rect 3233 15330 3299 15333
rect 4102 15330 4108 15332
rect 3233 15328 4108 15330
rect 3233 15272 3238 15328
rect 3294 15272 4108 15328
rect 3233 15270 4108 15272
rect 3233 15267 3299 15270
rect 4102 15268 4108 15270
rect 4172 15330 4178 15332
rect 4429 15330 4495 15333
rect 4172 15328 4495 15330
rect 4172 15272 4434 15328
rect 4490 15272 4495 15328
rect 4172 15270 4495 15272
rect 4172 15268 4178 15270
rect 4429 15267 4495 15270
rect 9254 15268 9260 15332
rect 9324 15330 9330 15332
rect 9397 15330 9463 15333
rect 9324 15328 9463 15330
rect 9324 15272 9402 15328
rect 9458 15272 9463 15328
rect 9324 15270 9463 15272
rect 9324 15268 9330 15270
rect 9397 15267 9463 15270
rect 4610 15264 4930 15265
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4930 15264
rect 4610 15199 4930 15200
rect 11944 15264 12264 15265
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 15199 12264 15200
rect 19277 15264 19597 15265
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 15199 19597 15200
rect 18822 14996 18828 15060
rect 18892 15058 18898 15060
rect 19149 15058 19215 15061
rect 18892 15056 19215 15058
rect 18892 15000 19154 15056
rect 19210 15000 19215 15056
rect 18892 14998 19215 15000
rect 18892 14996 18898 14998
rect 19149 14995 19215 14998
rect 13537 14922 13603 14925
rect 13721 14922 13787 14925
rect 13537 14920 13787 14922
rect 13537 14864 13542 14920
rect 13598 14864 13726 14920
rect 13782 14864 13787 14920
rect 13537 14862 13787 14864
rect 13537 14859 13603 14862
rect 13721 14859 13787 14862
rect 11329 14786 11395 14789
rect 11646 14786 11652 14788
rect 11329 14784 11652 14786
rect 11329 14728 11334 14784
rect 11390 14728 11652 14784
rect 11329 14726 11652 14728
rect 11329 14723 11395 14726
rect 11646 14724 11652 14726
rect 11716 14724 11722 14788
rect 8277 14720 8597 14721
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 14655 8597 14656
rect 15610 14720 15930 14721
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 14655 15930 14656
rect 5257 14514 5323 14517
rect 7782 14514 7788 14516
rect 5257 14512 7788 14514
rect 5257 14456 5262 14512
rect 5318 14456 7788 14512
rect 5257 14454 7788 14456
rect 5257 14451 5323 14454
rect 7782 14452 7788 14454
rect 7852 14514 7858 14516
rect 7925 14514 7991 14517
rect 9581 14516 9647 14517
rect 9581 14514 9628 14516
rect 7852 14512 7991 14514
rect 7852 14456 7930 14512
rect 7986 14456 7991 14512
rect 7852 14454 7991 14456
rect 9500 14512 9628 14514
rect 9692 14514 9698 14516
rect 19149 14514 19215 14517
rect 9692 14512 19215 14514
rect 9500 14456 9586 14512
rect 9692 14456 19154 14512
rect 19210 14456 19215 14512
rect 9500 14454 9628 14456
rect 7852 14452 7858 14454
rect 7925 14451 7991 14454
rect 9581 14452 9628 14454
rect 9692 14454 19215 14456
rect 9692 14452 9698 14454
rect 9581 14451 9647 14452
rect 19149 14451 19215 14454
rect 9857 14378 9923 14381
rect 13445 14378 13511 14381
rect 9857 14376 13511 14378
rect 9857 14320 9862 14376
rect 9918 14320 13450 14376
rect 13506 14320 13511 14376
rect 9857 14318 13511 14320
rect 9857 14315 9923 14318
rect 13445 14315 13511 14318
rect 12617 14242 12683 14245
rect 13261 14242 13327 14245
rect 12617 14240 13327 14242
rect 12617 14184 12622 14240
rect 12678 14184 13266 14240
rect 13322 14184 13327 14240
rect 12617 14182 13327 14184
rect 12617 14179 12683 14182
rect 13261 14179 13327 14182
rect 4610 14176 4930 14177
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4930 14176
rect 4610 14111 4930 14112
rect 11944 14176 12264 14177
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 14111 12264 14112
rect 19277 14176 19597 14177
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 14111 19597 14112
rect 11646 13908 11652 13972
rect 11716 13970 11722 13972
rect 12065 13970 12131 13973
rect 11716 13968 12131 13970
rect 11716 13912 12070 13968
rect 12126 13912 12131 13968
rect 11716 13910 12131 13912
rect 11716 13908 11722 13910
rect 12065 13907 12131 13910
rect 18137 13834 18203 13837
rect 17772 13832 18203 13834
rect 17772 13776 18142 13832
rect 18198 13776 18203 13832
rect 17772 13774 18203 13776
rect 0 13700 480 13728
rect 0 13636 60 13700
rect 124 13636 480 13700
rect 0 13608 480 13636
rect 17401 13698 17467 13701
rect 17772 13698 17832 13774
rect 18137 13771 18203 13774
rect 21520 13700 22000 13728
rect 21520 13698 21588 13700
rect 17401 13696 17832 13698
rect 17401 13640 17406 13696
rect 17462 13640 17832 13696
rect 17401 13638 17832 13640
rect 21460 13638 21588 13698
rect 17401 13635 17467 13638
rect 21520 13636 21588 13638
rect 21652 13636 22000 13700
rect 8277 13632 8597 13633
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 13567 8597 13568
rect 15610 13632 15930 13633
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 21520 13608 22000 13636
rect 15610 13567 15930 13568
rect 7833 13562 7899 13565
rect 7966 13562 7972 13564
rect 7833 13560 7972 13562
rect 7833 13504 7838 13560
rect 7894 13504 7972 13560
rect 7833 13502 7972 13504
rect 7833 13499 7899 13502
rect 7966 13500 7972 13502
rect 8036 13500 8042 13564
rect 17677 13562 17743 13565
rect 17677 13560 19350 13562
rect 17677 13504 17682 13560
rect 17738 13504 19350 13560
rect 17677 13502 19350 13504
rect 17677 13499 17743 13502
rect 54 13364 60 13428
rect 124 13426 130 13428
rect 1577 13426 1643 13429
rect 124 13424 1643 13426
rect 124 13368 1582 13424
rect 1638 13368 1643 13424
rect 124 13366 1643 13368
rect 124 13364 130 13366
rect 1577 13363 1643 13366
rect 4521 13426 4587 13429
rect 5206 13426 5212 13428
rect 4521 13424 5212 13426
rect 4521 13368 4526 13424
rect 4582 13368 5212 13424
rect 4521 13366 5212 13368
rect 4521 13363 4587 13366
rect 5206 13364 5212 13366
rect 5276 13364 5282 13428
rect 8017 13426 8083 13429
rect 14089 13426 14155 13429
rect 8017 13424 14155 13426
rect 8017 13368 8022 13424
rect 8078 13368 14094 13424
rect 14150 13368 14155 13424
rect 8017 13366 14155 13368
rect 19290 13426 19350 13502
rect 21582 13426 21588 13428
rect 19290 13366 21588 13426
rect 8017 13363 8083 13366
rect 14089 13363 14155 13366
rect 21582 13364 21588 13366
rect 21652 13364 21658 13428
rect 7782 13228 7788 13292
rect 7852 13290 7858 13292
rect 13813 13290 13879 13293
rect 7852 13288 13879 13290
rect 7852 13232 13818 13288
rect 13874 13232 13879 13288
rect 7852 13230 13879 13232
rect 7852 13228 7858 13230
rect 13813 13227 13879 13230
rect 4610 13088 4930 13089
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4930 13088
rect 4610 13023 4930 13024
rect 11944 13088 12264 13089
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 13023 12264 13024
rect 19277 13088 19597 13089
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 13023 19597 13024
rect 8277 12544 8597 12545
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 12479 8597 12480
rect 15610 12544 15930 12545
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 12479 15930 12480
rect 9213 12202 9279 12205
rect 9438 12202 9444 12204
rect 9213 12200 9444 12202
rect 9213 12144 9218 12200
rect 9274 12144 9444 12200
rect 9213 12142 9444 12144
rect 9213 12139 9279 12142
rect 9438 12140 9444 12142
rect 9508 12140 9514 12204
rect 4610 12000 4930 12001
rect 0 11928 480 11960
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4930 12000
rect 4610 11935 4930 11936
rect 11944 12000 12264 12001
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 11935 12264 11936
rect 19277 12000 19597 12001
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 11935 19597 11936
rect 0 11872 110 11928
rect 166 11872 480 11928
rect 0 11840 480 11872
rect 21520 11840 22000 11960
rect 4061 11658 4127 11661
rect 10593 11658 10659 11661
rect 4061 11656 10659 11658
rect 4061 11600 4066 11656
rect 4122 11600 10598 11656
rect 10654 11600 10659 11656
rect 4061 11598 10659 11600
rect 4061 11595 4127 11598
rect 10593 11595 10659 11598
rect 8277 11456 8597 11457
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 11391 8597 11392
rect 15610 11456 15930 11457
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 11391 15930 11392
rect 16113 11386 16179 11389
rect 21590 11386 21650 11840
rect 16113 11384 21650 11386
rect 16113 11328 16118 11384
rect 16174 11328 21650 11384
rect 16113 11326 21650 11328
rect 16113 11323 16179 11326
rect 4610 10912 4930 10913
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4930 10912
rect 4610 10847 4930 10848
rect 11944 10912 12264 10913
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 10847 12264 10848
rect 19277 10912 19597 10913
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 10847 19597 10848
rect 13353 10842 13419 10845
rect 13486 10842 13492 10844
rect 13353 10840 13492 10842
rect 13353 10784 13358 10840
rect 13414 10784 13492 10840
rect 13353 10782 13492 10784
rect 13353 10779 13419 10782
rect 13486 10780 13492 10782
rect 13556 10780 13562 10844
rect 1669 10706 1735 10709
rect 3417 10706 3483 10709
rect 1669 10704 3483 10706
rect 1669 10648 1674 10704
rect 1730 10648 3422 10704
rect 3478 10648 3483 10704
rect 1669 10646 3483 10648
rect 1669 10643 1735 10646
rect 3417 10643 3483 10646
rect 12985 10570 13051 10573
rect 12985 10568 21650 10570
rect 12985 10512 12990 10568
rect 13046 10512 21650 10568
rect 12985 10510 21650 10512
rect 12985 10507 13051 10510
rect 8277 10368 8597 10369
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 10303 8597 10304
rect 15610 10368 15930 10369
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 10303 15930 10304
rect 11278 10100 11284 10164
rect 11348 10162 11354 10164
rect 12801 10162 12867 10165
rect 11348 10160 12867 10162
rect 11348 10104 12806 10160
rect 12862 10104 12867 10160
rect 11348 10102 12867 10104
rect 11348 10100 11354 10102
rect 12801 10099 12867 10102
rect 13721 10162 13787 10165
rect 15285 10162 15351 10165
rect 13721 10160 15351 10162
rect 13721 10104 13726 10160
rect 13782 10104 15290 10160
rect 15346 10104 15351 10160
rect 13721 10102 15351 10104
rect 13721 10099 13787 10102
rect 15285 10099 15351 10102
rect 21590 10056 21650 10510
rect 0 9936 480 10056
rect 3877 10026 3943 10029
rect 5441 10026 5507 10029
rect 3877 10024 5507 10026
rect 3877 9968 3882 10024
rect 3938 9968 5446 10024
rect 5502 9968 5507 10024
rect 3877 9966 5507 9968
rect 3877 9963 3943 9966
rect 5441 9963 5507 9966
rect 21520 9936 22000 10056
rect 62 9482 122 9936
rect 4610 9824 4930 9825
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4930 9824
rect 4610 9759 4930 9760
rect 11944 9824 12264 9825
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 9759 12264 9760
rect 19277 9824 19597 9825
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 9759 19597 9760
rect 7598 9754 7604 9756
rect 5260 9694 7604 9754
rect 5260 9621 5320 9694
rect 7598 9692 7604 9694
rect 7668 9692 7674 9756
rect 2957 9618 3023 9621
rect 5257 9618 5323 9621
rect 2957 9616 5323 9618
rect 2957 9560 2962 9616
rect 3018 9560 5262 9616
rect 5318 9560 5323 9616
rect 2957 9558 5323 9560
rect 2957 9555 3023 9558
rect 5257 9555 5323 9558
rect 6729 9618 6795 9621
rect 9622 9618 9628 9620
rect 6729 9616 9628 9618
rect 6729 9560 6734 9616
rect 6790 9560 9628 9616
rect 6729 9558 9628 9560
rect 6729 9555 6795 9558
rect 9622 9556 9628 9558
rect 9692 9618 9698 9620
rect 11145 9618 11211 9621
rect 9692 9616 11211 9618
rect 9692 9560 11150 9616
rect 11206 9560 11211 9616
rect 9692 9558 11211 9560
rect 9692 9556 9698 9558
rect 11145 9555 11211 9558
rect 18822 9556 18828 9620
rect 18892 9618 18898 9620
rect 20069 9618 20135 9621
rect 18892 9616 20135 9618
rect 18892 9560 20074 9616
rect 20130 9560 20135 9616
rect 18892 9558 20135 9560
rect 18892 9556 18898 9558
rect 20069 9555 20135 9558
rect 1577 9482 1643 9485
rect 62 9480 1643 9482
rect 62 9424 1582 9480
rect 1638 9424 1643 9480
rect 62 9422 1643 9424
rect 1577 9419 1643 9422
rect 7833 9482 7899 9485
rect 15745 9482 15811 9485
rect 7833 9480 15811 9482
rect 7833 9424 7838 9480
rect 7894 9424 15750 9480
rect 15806 9424 15811 9480
rect 7833 9422 15811 9424
rect 7833 9419 7899 9422
rect 15745 9419 15811 9422
rect 8277 9280 8597 9281
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 9215 8597 9216
rect 15610 9280 15930 9281
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 9215 15930 9216
rect 381 9210 447 9213
rect 4429 9210 4495 9213
rect 381 9208 4495 9210
rect 381 9152 386 9208
rect 442 9152 4434 9208
rect 4490 9152 4495 9208
rect 381 9150 4495 9152
rect 381 9147 447 9150
rect 4429 9147 4495 9150
rect 9857 8938 9923 8941
rect 9990 8938 9996 8940
rect 9857 8936 9996 8938
rect 9857 8880 9862 8936
rect 9918 8880 9996 8936
rect 9857 8878 9996 8880
rect 9857 8875 9923 8878
rect 9990 8876 9996 8878
rect 10060 8876 10066 8940
rect 16665 8938 16731 8941
rect 16798 8938 16804 8940
rect 16665 8936 16804 8938
rect 16665 8880 16670 8936
rect 16726 8880 16804 8936
rect 16665 8878 16804 8880
rect 16665 8875 16731 8878
rect 16798 8876 16804 8878
rect 16868 8876 16874 8940
rect 4610 8736 4930 8737
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4930 8736
rect 4610 8671 4930 8672
rect 11944 8736 12264 8737
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 8671 12264 8672
rect 19277 8736 19597 8737
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 8671 19597 8672
rect 105 8530 171 8533
rect 5625 8530 5691 8533
rect 105 8528 5691 8530
rect 105 8472 110 8528
rect 166 8472 5630 8528
rect 5686 8472 5691 8528
rect 105 8470 5691 8472
rect 105 8467 171 8470
rect 5625 8467 5691 8470
rect 0 8256 480 8288
rect 21520 8258 22000 8288
rect 0 8200 110 8256
rect 166 8200 480 8256
rect 0 8168 480 8200
rect 21460 8256 22000 8258
rect 21460 8200 21546 8256
rect 21602 8200 22000 8256
rect 21460 8198 22000 8200
rect 8277 8192 8597 8193
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 8127 8597 8128
rect 15610 8192 15930 8193
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 21520 8168 22000 8198
rect 15610 8127 15930 8128
rect 8661 7986 8727 7989
rect 9070 7986 9076 7988
rect 8661 7984 9076 7986
rect 8661 7928 8666 7984
rect 8722 7928 9076 7984
rect 8661 7926 9076 7928
rect 8661 7923 8727 7926
rect 9070 7924 9076 7926
rect 9140 7924 9146 7988
rect 4610 7648 4930 7649
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4930 7648
rect 4610 7583 4930 7584
rect 11944 7648 12264 7649
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 7583 12264 7584
rect 19277 7648 19597 7649
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 7583 19597 7584
rect 8277 7104 8597 7105
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 7039 8597 7040
rect 15610 7104 15930 7105
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 7039 15930 7040
rect 54 6700 60 6764
rect 124 6762 130 6764
rect 4245 6762 4311 6765
rect 124 6760 4311 6762
rect 124 6704 4250 6760
rect 4306 6704 4311 6760
rect 124 6702 4311 6704
rect 124 6700 130 6702
rect 4245 6699 4311 6702
rect 4610 6560 4930 6561
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4930 6560
rect 4610 6495 4930 6496
rect 11944 6560 12264 6561
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 6495 12264 6496
rect 19277 6560 19597 6561
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 6495 19597 6496
rect 0 6356 480 6384
rect 0 6292 60 6356
rect 124 6292 480 6356
rect 0 6264 480 6292
rect 2865 6354 2931 6357
rect 7966 6354 7972 6356
rect 2865 6352 7972 6354
rect 2865 6296 2870 6352
rect 2926 6296 7972 6352
rect 2865 6294 7972 6296
rect 2865 6291 2931 6294
rect 7966 6292 7972 6294
rect 8036 6354 8042 6356
rect 16021 6354 16087 6357
rect 21520 6354 22000 6384
rect 8036 6352 16087 6354
rect 8036 6296 16026 6352
rect 16082 6296 16087 6352
rect 8036 6294 16087 6296
rect 21460 6352 22000 6354
rect 21460 6296 21546 6352
rect 21602 6296 22000 6352
rect 21460 6294 22000 6296
rect 8036 6292 8042 6294
rect 16021 6291 16087 6294
rect 21520 6264 22000 6294
rect 8277 6016 8597 6017
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 5951 8597 5952
rect 15610 6016 15930 6017
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 5951 15930 5952
rect 5206 5748 5212 5812
rect 5276 5810 5282 5812
rect 8201 5810 8267 5813
rect 5276 5808 8267 5810
rect 5276 5752 8206 5808
rect 8262 5752 8267 5808
rect 5276 5750 8267 5752
rect 5276 5748 5282 5750
rect 8201 5747 8267 5750
rect 5257 5674 5323 5677
rect 10869 5674 10935 5677
rect 5257 5672 10935 5674
rect 5257 5616 5262 5672
rect 5318 5616 10874 5672
rect 10930 5616 10935 5672
rect 5257 5614 10935 5616
rect 5257 5611 5323 5614
rect 10869 5611 10935 5614
rect 4610 5472 4930 5473
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4930 5472
rect 4610 5407 4930 5408
rect 11944 5472 12264 5473
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 5407 12264 5408
rect 19277 5472 19597 5473
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 5407 19597 5408
rect 2313 5266 2379 5269
rect 2957 5266 3023 5269
rect 5257 5266 5323 5269
rect 9254 5266 9260 5268
rect 2313 5264 9260 5266
rect 2313 5208 2318 5264
rect 2374 5208 2962 5264
rect 3018 5208 5262 5264
rect 5318 5208 9260 5264
rect 2313 5206 9260 5208
rect 2313 5203 2379 5206
rect 2957 5203 3023 5206
rect 5257 5203 5323 5206
rect 9254 5204 9260 5206
rect 9324 5266 9330 5268
rect 15193 5266 15259 5269
rect 9324 5264 15259 5266
rect 9324 5208 15198 5264
rect 15254 5208 15259 5264
rect 9324 5206 15259 5208
rect 9324 5204 9330 5206
rect 15193 5203 15259 5206
rect 3601 5130 3667 5133
rect 11697 5130 11763 5133
rect 3601 5128 11763 5130
rect 3601 5072 3606 5128
rect 3662 5072 11702 5128
rect 11758 5072 11763 5128
rect 3601 5070 11763 5072
rect 3601 5067 3667 5070
rect 11697 5067 11763 5070
rect 5073 4994 5139 4997
rect 7833 4994 7899 4997
rect 5073 4992 7899 4994
rect 5073 4936 5078 4992
rect 5134 4936 7838 4992
rect 7894 4936 7899 4992
rect 5073 4934 7899 4936
rect 5073 4931 5139 4934
rect 7833 4931 7899 4934
rect 8277 4928 8597 4929
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 4863 8597 4864
rect 15610 4928 15930 4929
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 4863 15930 4864
rect 2773 4722 2839 4725
rect 8753 4722 8819 4725
rect 14825 4722 14891 4725
rect 2773 4720 14891 4722
rect 2773 4664 2778 4720
rect 2834 4664 8758 4720
rect 8814 4664 14830 4720
rect 14886 4664 14891 4720
rect 2773 4662 14891 4664
rect 2773 4659 2839 4662
rect 8753 4659 8819 4662
rect 14825 4659 14891 4662
rect 0 4496 480 4616
rect 4061 4586 4127 4589
rect 10593 4586 10659 4589
rect 4061 4584 10659 4586
rect 4061 4528 4066 4584
rect 4122 4528 10598 4584
rect 10654 4528 10659 4584
rect 4061 4526 10659 4528
rect 4061 4523 4127 4526
rect 10593 4523 10659 4526
rect 12617 4586 12683 4589
rect 17125 4586 17191 4589
rect 12617 4584 17191 4586
rect 12617 4528 12622 4584
rect 12678 4528 17130 4584
rect 17186 4528 17191 4584
rect 12617 4526 17191 4528
rect 12617 4523 12683 4526
rect 17125 4523 17191 4526
rect 19149 4586 19215 4589
rect 19425 4586 19491 4589
rect 21520 4586 22000 4616
rect 19149 4584 22000 4586
rect 19149 4528 19154 4584
rect 19210 4528 19430 4584
rect 19486 4528 22000 4584
rect 19149 4526 22000 4528
rect 19149 4523 19215 4526
rect 19425 4523 19491 4526
rect 21520 4496 22000 4526
rect 62 4042 122 4496
rect 5206 4388 5212 4452
rect 5276 4450 5282 4452
rect 5349 4450 5415 4453
rect 5276 4448 5415 4450
rect 5276 4392 5354 4448
rect 5410 4392 5415 4448
rect 5276 4390 5415 4392
rect 5276 4388 5282 4390
rect 5349 4387 5415 4390
rect 4610 4384 4930 4385
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4930 4384
rect 4610 4319 4930 4320
rect 11944 4384 12264 4385
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 4319 12264 4320
rect 19277 4384 19597 4385
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 4319 19597 4320
rect 1761 4314 1827 4317
rect 4245 4314 4311 4317
rect 9765 4314 9831 4317
rect 1761 4312 4311 4314
rect 1761 4256 1766 4312
rect 1822 4256 4250 4312
rect 4306 4256 4311 4312
rect 1761 4254 4311 4256
rect 1761 4251 1827 4254
rect 4245 4251 4311 4254
rect 9630 4312 9831 4314
rect 9630 4256 9770 4312
rect 9826 4256 9831 4312
rect 9630 4254 9831 4256
rect 2313 4178 2379 4181
rect 9630 4178 9690 4254
rect 9765 4251 9831 4254
rect 2313 4176 9690 4178
rect 2313 4120 2318 4176
rect 2374 4120 9690 4176
rect 2313 4118 9690 4120
rect 9768 4178 9828 4251
rect 17769 4178 17835 4181
rect 9768 4176 17835 4178
rect 9768 4120 17774 4176
rect 17830 4120 17835 4176
rect 9768 4118 17835 4120
rect 2313 4115 2379 4118
rect 17769 4115 17835 4118
rect 4245 4042 4311 4045
rect 62 4040 4311 4042
rect 62 3984 4250 4040
rect 4306 3984 4311 4040
rect 62 3982 4311 3984
rect 4245 3979 4311 3982
rect 8109 4042 8175 4045
rect 8569 4042 8635 4045
rect 8109 4040 8635 4042
rect 8109 3984 8114 4040
rect 8170 3984 8574 4040
rect 8630 3984 8635 4040
rect 8109 3982 8635 3984
rect 8109 3979 8175 3982
rect 8569 3979 8635 3982
rect 8277 3840 8597 3841
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 3775 8597 3776
rect 15610 3840 15930 3841
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 3775 15930 3776
rect 6678 3436 6684 3500
rect 6748 3498 6754 3500
rect 7189 3498 7255 3501
rect 18873 3498 18939 3501
rect 6748 3496 18939 3498
rect 6748 3440 7194 3496
rect 7250 3440 18878 3496
rect 18934 3440 18939 3496
rect 6748 3438 18939 3440
rect 6748 3436 6754 3438
rect 7189 3435 7255 3438
rect 18873 3435 18939 3438
rect 4610 3296 4930 3297
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4930 3296
rect 4610 3231 4930 3232
rect 11944 3296 12264 3297
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 3231 12264 3232
rect 19277 3296 19597 3297
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 3231 19597 3232
rect 1577 3226 1643 3229
rect 62 3224 1643 3226
rect 62 3168 1582 3224
rect 1638 3168 1643 3224
rect 62 3166 1643 3168
rect 62 2712 122 3166
rect 1577 3163 1643 3166
rect 16021 3090 16087 3093
rect 16021 3088 21650 3090
rect 16021 3032 16026 3088
rect 16082 3032 21650 3088
rect 16021 3030 21650 3032
rect 16021 3027 16087 3030
rect 2037 2954 2103 2957
rect 9121 2954 9187 2957
rect 2037 2952 9187 2954
rect 2037 2896 2042 2952
rect 2098 2896 9126 2952
rect 9182 2896 9187 2952
rect 2037 2894 9187 2896
rect 2037 2891 2103 2894
rect 9121 2891 9187 2894
rect 8277 2752 8597 2753
rect 0 2592 480 2712
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2687 8597 2688
rect 15610 2752 15930 2753
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 21590 2712 21650 3030
rect 15610 2687 15930 2688
rect 21520 2592 22000 2712
rect 4102 2484 4108 2548
rect 4172 2546 4178 2548
rect 4613 2546 4679 2549
rect 13353 2546 13419 2549
rect 4172 2544 13419 2546
rect 4172 2488 4618 2544
rect 4674 2488 13358 2544
rect 13414 2488 13419 2544
rect 4172 2486 13419 2488
rect 4172 2484 4178 2486
rect 4613 2483 4679 2486
rect 13353 2483 13419 2486
rect 1945 2410 2011 2413
rect 11237 2410 11303 2413
rect 1945 2408 11303 2410
rect 1945 2352 1950 2408
rect 2006 2352 11242 2408
rect 11298 2352 11303 2408
rect 1945 2350 11303 2352
rect 1945 2347 2011 2350
rect 11237 2347 11303 2350
rect 4610 2208 4930 2209
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4930 2208
rect 4610 2143 4930 2144
rect 11944 2208 12264 2209
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2143 12264 2144
rect 19277 2208 19597 2209
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2143 19597 2144
rect 2773 1458 2839 1461
rect 62 1456 2839 1458
rect 62 1400 2778 1456
rect 2834 1400 2839 1456
rect 62 1398 2839 1400
rect 62 944 122 1398
rect 2773 1395 2839 1398
rect 8702 1396 8708 1460
rect 8772 1458 8778 1460
rect 20345 1458 20411 1461
rect 8772 1456 20411 1458
rect 8772 1400 20350 1456
rect 20406 1400 20411 1456
rect 8772 1398 20411 1400
rect 8772 1396 8778 1398
rect 20345 1395 20411 1398
rect 17953 1322 18019 1325
rect 17953 1320 21650 1322
rect 17953 1264 17958 1320
rect 18014 1264 21650 1320
rect 17953 1262 21650 1264
rect 17953 1259 18019 1262
rect 21590 944 21650 1262
rect 0 824 480 944
rect 21520 824 22000 944
<< via3 >>
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 4698 19612 4762 19616
rect 4698 19556 4702 19612
rect 4702 19556 4758 19612
rect 4758 19556 4762 19612
rect 4698 19552 4762 19556
rect 4778 19612 4842 19616
rect 4778 19556 4782 19612
rect 4782 19556 4838 19612
rect 4838 19556 4842 19612
rect 4778 19552 4842 19556
rect 4858 19612 4922 19616
rect 4858 19556 4862 19612
rect 4862 19556 4918 19612
rect 4918 19556 4922 19612
rect 4858 19552 4922 19556
rect 11952 19612 12016 19616
rect 11952 19556 11956 19612
rect 11956 19556 12012 19612
rect 12012 19556 12016 19612
rect 11952 19552 12016 19556
rect 12032 19612 12096 19616
rect 12032 19556 12036 19612
rect 12036 19556 12092 19612
rect 12092 19556 12096 19612
rect 12032 19552 12096 19556
rect 12112 19612 12176 19616
rect 12112 19556 12116 19612
rect 12116 19556 12172 19612
rect 12172 19556 12176 19612
rect 12112 19552 12176 19556
rect 12192 19612 12256 19616
rect 12192 19556 12196 19612
rect 12196 19556 12252 19612
rect 12252 19556 12256 19612
rect 12192 19552 12256 19556
rect 19285 19612 19349 19616
rect 19285 19556 19289 19612
rect 19289 19556 19345 19612
rect 19345 19556 19349 19612
rect 19285 19552 19349 19556
rect 19365 19612 19429 19616
rect 19365 19556 19369 19612
rect 19369 19556 19425 19612
rect 19425 19556 19429 19612
rect 19365 19552 19429 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 8285 19068 8349 19072
rect 8285 19012 8289 19068
rect 8289 19012 8345 19068
rect 8345 19012 8349 19068
rect 8285 19008 8349 19012
rect 8365 19068 8429 19072
rect 8365 19012 8369 19068
rect 8369 19012 8425 19068
rect 8425 19012 8429 19068
rect 8365 19008 8429 19012
rect 8445 19068 8509 19072
rect 8445 19012 8449 19068
rect 8449 19012 8505 19068
rect 8505 19012 8509 19068
rect 8445 19008 8509 19012
rect 8525 19068 8589 19072
rect 8525 19012 8529 19068
rect 8529 19012 8585 19068
rect 8585 19012 8589 19068
rect 8525 19008 8589 19012
rect 15618 19068 15682 19072
rect 15618 19012 15622 19068
rect 15622 19012 15678 19068
rect 15678 19012 15682 19068
rect 15618 19008 15682 19012
rect 15698 19068 15762 19072
rect 15698 19012 15702 19068
rect 15702 19012 15758 19068
rect 15758 19012 15762 19068
rect 15698 19008 15762 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 4698 18524 4762 18528
rect 4698 18468 4702 18524
rect 4702 18468 4758 18524
rect 4758 18468 4762 18524
rect 4698 18464 4762 18468
rect 4778 18524 4842 18528
rect 4778 18468 4782 18524
rect 4782 18468 4838 18524
rect 4838 18468 4842 18524
rect 4778 18464 4842 18468
rect 4858 18524 4922 18528
rect 4858 18468 4862 18524
rect 4862 18468 4918 18524
rect 4918 18468 4922 18524
rect 4858 18464 4922 18468
rect 11952 18524 12016 18528
rect 11952 18468 11956 18524
rect 11956 18468 12012 18524
rect 12012 18468 12016 18524
rect 11952 18464 12016 18468
rect 12032 18524 12096 18528
rect 12032 18468 12036 18524
rect 12036 18468 12092 18524
rect 12092 18468 12096 18524
rect 12032 18464 12096 18468
rect 12112 18524 12176 18528
rect 12112 18468 12116 18524
rect 12116 18468 12172 18524
rect 12172 18468 12176 18524
rect 12112 18464 12176 18468
rect 12192 18524 12256 18528
rect 12192 18468 12196 18524
rect 12196 18468 12252 18524
rect 12252 18468 12256 18524
rect 12192 18464 12256 18468
rect 19285 18524 19349 18528
rect 19285 18468 19289 18524
rect 19289 18468 19345 18524
rect 19345 18468 19349 18524
rect 19285 18464 19349 18468
rect 19365 18524 19429 18528
rect 19365 18468 19369 18524
rect 19369 18468 19425 18524
rect 19425 18468 19429 18524
rect 19365 18464 19429 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 16804 18048 16868 18052
rect 16804 17992 16818 18048
rect 16818 17992 16868 18048
rect 16804 17988 16868 17992
rect 8285 17980 8349 17984
rect 8285 17924 8289 17980
rect 8289 17924 8345 17980
rect 8345 17924 8349 17980
rect 8285 17920 8349 17924
rect 8365 17980 8429 17984
rect 8365 17924 8369 17980
rect 8369 17924 8425 17980
rect 8425 17924 8429 17980
rect 8365 17920 8429 17924
rect 8445 17980 8509 17984
rect 8445 17924 8449 17980
rect 8449 17924 8505 17980
rect 8505 17924 8509 17980
rect 8445 17920 8509 17924
rect 8525 17980 8589 17984
rect 8525 17924 8529 17980
rect 8529 17924 8585 17980
rect 8585 17924 8589 17980
rect 8525 17920 8589 17924
rect 15618 17980 15682 17984
rect 15618 17924 15622 17980
rect 15622 17924 15678 17980
rect 15678 17924 15682 17980
rect 15618 17920 15682 17924
rect 15698 17980 15762 17984
rect 15698 17924 15702 17980
rect 15702 17924 15758 17980
rect 15758 17924 15762 17980
rect 15698 17920 15762 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 4698 17436 4762 17440
rect 4698 17380 4702 17436
rect 4702 17380 4758 17436
rect 4758 17380 4762 17436
rect 4698 17376 4762 17380
rect 4778 17436 4842 17440
rect 4778 17380 4782 17436
rect 4782 17380 4838 17436
rect 4838 17380 4842 17436
rect 4778 17376 4842 17380
rect 4858 17436 4922 17440
rect 4858 17380 4862 17436
rect 4862 17380 4918 17436
rect 4918 17380 4922 17436
rect 4858 17376 4922 17380
rect 11952 17436 12016 17440
rect 11952 17380 11956 17436
rect 11956 17380 12012 17436
rect 12012 17380 12016 17436
rect 11952 17376 12016 17380
rect 12032 17436 12096 17440
rect 12032 17380 12036 17436
rect 12036 17380 12092 17436
rect 12092 17380 12096 17436
rect 12032 17376 12096 17380
rect 12112 17436 12176 17440
rect 12112 17380 12116 17436
rect 12116 17380 12172 17436
rect 12172 17380 12176 17436
rect 12112 17376 12176 17380
rect 12192 17436 12256 17440
rect 12192 17380 12196 17436
rect 12196 17380 12252 17436
rect 12252 17380 12256 17436
rect 12192 17376 12256 17380
rect 19285 17436 19349 17440
rect 19285 17380 19289 17436
rect 19289 17380 19345 17436
rect 19345 17380 19349 17436
rect 19285 17376 19349 17380
rect 19365 17436 19429 17440
rect 19365 17380 19369 17436
rect 19369 17380 19425 17436
rect 19425 17380 19429 17436
rect 19365 17376 19429 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 13492 17172 13556 17236
rect 7604 16900 7668 16964
rect 9996 16900 10060 16964
rect 8285 16892 8349 16896
rect 8285 16836 8289 16892
rect 8289 16836 8345 16892
rect 8345 16836 8349 16892
rect 8285 16832 8349 16836
rect 8365 16892 8429 16896
rect 8365 16836 8369 16892
rect 8369 16836 8425 16892
rect 8425 16836 8429 16892
rect 8365 16832 8429 16836
rect 8445 16892 8509 16896
rect 8445 16836 8449 16892
rect 8449 16836 8505 16892
rect 8505 16836 8509 16892
rect 8445 16832 8509 16836
rect 8525 16892 8589 16896
rect 8525 16836 8529 16892
rect 8529 16836 8585 16892
rect 8585 16836 8589 16892
rect 8525 16832 8589 16836
rect 15618 16892 15682 16896
rect 15618 16836 15622 16892
rect 15622 16836 15678 16892
rect 15678 16836 15682 16892
rect 15618 16832 15682 16836
rect 15698 16892 15762 16896
rect 15698 16836 15702 16892
rect 15702 16836 15758 16892
rect 15758 16836 15762 16892
rect 15698 16832 15762 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 9444 16764 9508 16828
rect 9076 16492 9140 16556
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 4698 16348 4762 16352
rect 4698 16292 4702 16348
rect 4702 16292 4758 16348
rect 4758 16292 4762 16348
rect 4698 16288 4762 16292
rect 4778 16348 4842 16352
rect 4778 16292 4782 16348
rect 4782 16292 4838 16348
rect 4838 16292 4842 16348
rect 4778 16288 4842 16292
rect 4858 16348 4922 16352
rect 4858 16292 4862 16348
rect 4862 16292 4918 16348
rect 4918 16292 4922 16348
rect 4858 16288 4922 16292
rect 11952 16348 12016 16352
rect 11952 16292 11956 16348
rect 11956 16292 12012 16348
rect 12012 16292 12016 16348
rect 11952 16288 12016 16292
rect 12032 16348 12096 16352
rect 12032 16292 12036 16348
rect 12036 16292 12092 16348
rect 12092 16292 12096 16348
rect 12032 16288 12096 16292
rect 12112 16348 12176 16352
rect 12112 16292 12116 16348
rect 12116 16292 12172 16348
rect 12172 16292 12176 16348
rect 12112 16288 12176 16292
rect 12192 16348 12256 16352
rect 12192 16292 12196 16348
rect 12196 16292 12252 16348
rect 12252 16292 12256 16348
rect 12192 16288 12256 16292
rect 19285 16348 19349 16352
rect 19285 16292 19289 16348
rect 19289 16292 19345 16348
rect 19345 16292 19349 16348
rect 19285 16288 19349 16292
rect 19365 16348 19429 16352
rect 19365 16292 19369 16348
rect 19369 16292 19425 16348
rect 19425 16292 19429 16348
rect 19365 16288 19429 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 8708 16220 8772 16284
rect 6684 16008 6748 16012
rect 6684 15952 6698 16008
rect 6698 15952 6748 16008
rect 6684 15948 6748 15952
rect 11284 15812 11348 15876
rect 8285 15804 8349 15808
rect 8285 15748 8289 15804
rect 8289 15748 8345 15804
rect 8345 15748 8349 15804
rect 8285 15744 8349 15748
rect 8365 15804 8429 15808
rect 8365 15748 8369 15804
rect 8369 15748 8425 15804
rect 8425 15748 8429 15804
rect 8365 15744 8429 15748
rect 8445 15804 8509 15808
rect 8445 15748 8449 15804
rect 8449 15748 8505 15804
rect 8505 15748 8509 15804
rect 8445 15744 8509 15748
rect 8525 15804 8589 15808
rect 8525 15748 8529 15804
rect 8529 15748 8585 15804
rect 8585 15748 8589 15804
rect 8525 15744 8589 15748
rect 15618 15804 15682 15808
rect 15618 15748 15622 15804
rect 15622 15748 15678 15804
rect 15678 15748 15682 15804
rect 15618 15744 15682 15748
rect 15698 15804 15762 15808
rect 15698 15748 15702 15804
rect 15702 15748 15758 15804
rect 15758 15748 15762 15804
rect 15698 15744 15762 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 4108 15268 4172 15332
rect 9260 15268 9324 15332
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 4698 15260 4762 15264
rect 4698 15204 4702 15260
rect 4702 15204 4758 15260
rect 4758 15204 4762 15260
rect 4698 15200 4762 15204
rect 4778 15260 4842 15264
rect 4778 15204 4782 15260
rect 4782 15204 4838 15260
rect 4838 15204 4842 15260
rect 4778 15200 4842 15204
rect 4858 15260 4922 15264
rect 4858 15204 4862 15260
rect 4862 15204 4918 15260
rect 4918 15204 4922 15260
rect 4858 15200 4922 15204
rect 11952 15260 12016 15264
rect 11952 15204 11956 15260
rect 11956 15204 12012 15260
rect 12012 15204 12016 15260
rect 11952 15200 12016 15204
rect 12032 15260 12096 15264
rect 12032 15204 12036 15260
rect 12036 15204 12092 15260
rect 12092 15204 12096 15260
rect 12032 15200 12096 15204
rect 12112 15260 12176 15264
rect 12112 15204 12116 15260
rect 12116 15204 12172 15260
rect 12172 15204 12176 15260
rect 12112 15200 12176 15204
rect 12192 15260 12256 15264
rect 12192 15204 12196 15260
rect 12196 15204 12252 15260
rect 12252 15204 12256 15260
rect 12192 15200 12256 15204
rect 19285 15260 19349 15264
rect 19285 15204 19289 15260
rect 19289 15204 19345 15260
rect 19345 15204 19349 15260
rect 19285 15200 19349 15204
rect 19365 15260 19429 15264
rect 19365 15204 19369 15260
rect 19369 15204 19425 15260
rect 19425 15204 19429 15260
rect 19365 15200 19429 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 18828 14996 18892 15060
rect 11652 14724 11716 14788
rect 8285 14716 8349 14720
rect 8285 14660 8289 14716
rect 8289 14660 8345 14716
rect 8345 14660 8349 14716
rect 8285 14656 8349 14660
rect 8365 14716 8429 14720
rect 8365 14660 8369 14716
rect 8369 14660 8425 14716
rect 8425 14660 8429 14716
rect 8365 14656 8429 14660
rect 8445 14716 8509 14720
rect 8445 14660 8449 14716
rect 8449 14660 8505 14716
rect 8505 14660 8509 14716
rect 8445 14656 8509 14660
rect 8525 14716 8589 14720
rect 8525 14660 8529 14716
rect 8529 14660 8585 14716
rect 8585 14660 8589 14716
rect 8525 14656 8589 14660
rect 15618 14716 15682 14720
rect 15618 14660 15622 14716
rect 15622 14660 15678 14716
rect 15678 14660 15682 14716
rect 15618 14656 15682 14660
rect 15698 14716 15762 14720
rect 15698 14660 15702 14716
rect 15702 14660 15758 14716
rect 15758 14660 15762 14716
rect 15698 14656 15762 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 7788 14452 7852 14516
rect 9628 14512 9692 14516
rect 9628 14456 9642 14512
rect 9642 14456 9692 14512
rect 9628 14452 9692 14456
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 4698 14172 4762 14176
rect 4698 14116 4702 14172
rect 4702 14116 4758 14172
rect 4758 14116 4762 14172
rect 4698 14112 4762 14116
rect 4778 14172 4842 14176
rect 4778 14116 4782 14172
rect 4782 14116 4838 14172
rect 4838 14116 4842 14172
rect 4778 14112 4842 14116
rect 4858 14172 4922 14176
rect 4858 14116 4862 14172
rect 4862 14116 4918 14172
rect 4918 14116 4922 14172
rect 4858 14112 4922 14116
rect 11952 14172 12016 14176
rect 11952 14116 11956 14172
rect 11956 14116 12012 14172
rect 12012 14116 12016 14172
rect 11952 14112 12016 14116
rect 12032 14172 12096 14176
rect 12032 14116 12036 14172
rect 12036 14116 12092 14172
rect 12092 14116 12096 14172
rect 12032 14112 12096 14116
rect 12112 14172 12176 14176
rect 12112 14116 12116 14172
rect 12116 14116 12172 14172
rect 12172 14116 12176 14172
rect 12112 14112 12176 14116
rect 12192 14172 12256 14176
rect 12192 14116 12196 14172
rect 12196 14116 12252 14172
rect 12252 14116 12256 14172
rect 12192 14112 12256 14116
rect 19285 14172 19349 14176
rect 19285 14116 19289 14172
rect 19289 14116 19345 14172
rect 19345 14116 19349 14172
rect 19285 14112 19349 14116
rect 19365 14172 19429 14176
rect 19365 14116 19369 14172
rect 19369 14116 19425 14172
rect 19425 14116 19429 14172
rect 19365 14112 19429 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 11652 13908 11716 13972
rect 60 13636 124 13700
rect 21588 13636 21652 13700
rect 8285 13628 8349 13632
rect 8285 13572 8289 13628
rect 8289 13572 8345 13628
rect 8345 13572 8349 13628
rect 8285 13568 8349 13572
rect 8365 13628 8429 13632
rect 8365 13572 8369 13628
rect 8369 13572 8425 13628
rect 8425 13572 8429 13628
rect 8365 13568 8429 13572
rect 8445 13628 8509 13632
rect 8445 13572 8449 13628
rect 8449 13572 8505 13628
rect 8505 13572 8509 13628
rect 8445 13568 8509 13572
rect 8525 13628 8589 13632
rect 8525 13572 8529 13628
rect 8529 13572 8585 13628
rect 8585 13572 8589 13628
rect 8525 13568 8589 13572
rect 15618 13628 15682 13632
rect 15618 13572 15622 13628
rect 15622 13572 15678 13628
rect 15678 13572 15682 13628
rect 15618 13568 15682 13572
rect 15698 13628 15762 13632
rect 15698 13572 15702 13628
rect 15702 13572 15758 13628
rect 15758 13572 15762 13628
rect 15698 13568 15762 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 7972 13500 8036 13564
rect 60 13364 124 13428
rect 5212 13364 5276 13428
rect 21588 13364 21652 13428
rect 7788 13228 7852 13292
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 4698 13084 4762 13088
rect 4698 13028 4702 13084
rect 4702 13028 4758 13084
rect 4758 13028 4762 13084
rect 4698 13024 4762 13028
rect 4778 13084 4842 13088
rect 4778 13028 4782 13084
rect 4782 13028 4838 13084
rect 4838 13028 4842 13084
rect 4778 13024 4842 13028
rect 4858 13084 4922 13088
rect 4858 13028 4862 13084
rect 4862 13028 4918 13084
rect 4918 13028 4922 13084
rect 4858 13024 4922 13028
rect 11952 13084 12016 13088
rect 11952 13028 11956 13084
rect 11956 13028 12012 13084
rect 12012 13028 12016 13084
rect 11952 13024 12016 13028
rect 12032 13084 12096 13088
rect 12032 13028 12036 13084
rect 12036 13028 12092 13084
rect 12092 13028 12096 13084
rect 12032 13024 12096 13028
rect 12112 13084 12176 13088
rect 12112 13028 12116 13084
rect 12116 13028 12172 13084
rect 12172 13028 12176 13084
rect 12112 13024 12176 13028
rect 12192 13084 12256 13088
rect 12192 13028 12196 13084
rect 12196 13028 12252 13084
rect 12252 13028 12256 13084
rect 12192 13024 12256 13028
rect 19285 13084 19349 13088
rect 19285 13028 19289 13084
rect 19289 13028 19345 13084
rect 19345 13028 19349 13084
rect 19285 13024 19349 13028
rect 19365 13084 19429 13088
rect 19365 13028 19369 13084
rect 19369 13028 19425 13084
rect 19425 13028 19429 13084
rect 19365 13024 19429 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 8285 12540 8349 12544
rect 8285 12484 8289 12540
rect 8289 12484 8345 12540
rect 8345 12484 8349 12540
rect 8285 12480 8349 12484
rect 8365 12540 8429 12544
rect 8365 12484 8369 12540
rect 8369 12484 8425 12540
rect 8425 12484 8429 12540
rect 8365 12480 8429 12484
rect 8445 12540 8509 12544
rect 8445 12484 8449 12540
rect 8449 12484 8505 12540
rect 8505 12484 8509 12540
rect 8445 12480 8509 12484
rect 8525 12540 8589 12544
rect 8525 12484 8529 12540
rect 8529 12484 8585 12540
rect 8585 12484 8589 12540
rect 8525 12480 8589 12484
rect 15618 12540 15682 12544
rect 15618 12484 15622 12540
rect 15622 12484 15678 12540
rect 15678 12484 15682 12540
rect 15618 12480 15682 12484
rect 15698 12540 15762 12544
rect 15698 12484 15702 12540
rect 15702 12484 15758 12540
rect 15758 12484 15762 12540
rect 15698 12480 15762 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 9444 12140 9508 12204
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 4698 11996 4762 12000
rect 4698 11940 4702 11996
rect 4702 11940 4758 11996
rect 4758 11940 4762 11996
rect 4698 11936 4762 11940
rect 4778 11996 4842 12000
rect 4778 11940 4782 11996
rect 4782 11940 4838 11996
rect 4838 11940 4842 11996
rect 4778 11936 4842 11940
rect 4858 11996 4922 12000
rect 4858 11940 4862 11996
rect 4862 11940 4918 11996
rect 4918 11940 4922 11996
rect 4858 11936 4922 11940
rect 11952 11996 12016 12000
rect 11952 11940 11956 11996
rect 11956 11940 12012 11996
rect 12012 11940 12016 11996
rect 11952 11936 12016 11940
rect 12032 11996 12096 12000
rect 12032 11940 12036 11996
rect 12036 11940 12092 11996
rect 12092 11940 12096 11996
rect 12032 11936 12096 11940
rect 12112 11996 12176 12000
rect 12112 11940 12116 11996
rect 12116 11940 12172 11996
rect 12172 11940 12176 11996
rect 12112 11936 12176 11940
rect 12192 11996 12256 12000
rect 12192 11940 12196 11996
rect 12196 11940 12252 11996
rect 12252 11940 12256 11996
rect 12192 11936 12256 11940
rect 19285 11996 19349 12000
rect 19285 11940 19289 11996
rect 19289 11940 19345 11996
rect 19345 11940 19349 11996
rect 19285 11936 19349 11940
rect 19365 11996 19429 12000
rect 19365 11940 19369 11996
rect 19369 11940 19425 11996
rect 19425 11940 19429 11996
rect 19365 11936 19429 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 8285 11452 8349 11456
rect 8285 11396 8289 11452
rect 8289 11396 8345 11452
rect 8345 11396 8349 11452
rect 8285 11392 8349 11396
rect 8365 11452 8429 11456
rect 8365 11396 8369 11452
rect 8369 11396 8425 11452
rect 8425 11396 8429 11452
rect 8365 11392 8429 11396
rect 8445 11452 8509 11456
rect 8445 11396 8449 11452
rect 8449 11396 8505 11452
rect 8505 11396 8509 11452
rect 8445 11392 8509 11396
rect 8525 11452 8589 11456
rect 8525 11396 8529 11452
rect 8529 11396 8585 11452
rect 8585 11396 8589 11452
rect 8525 11392 8589 11396
rect 15618 11452 15682 11456
rect 15618 11396 15622 11452
rect 15622 11396 15678 11452
rect 15678 11396 15682 11452
rect 15618 11392 15682 11396
rect 15698 11452 15762 11456
rect 15698 11396 15702 11452
rect 15702 11396 15758 11452
rect 15758 11396 15762 11452
rect 15698 11392 15762 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 4698 10908 4762 10912
rect 4698 10852 4702 10908
rect 4702 10852 4758 10908
rect 4758 10852 4762 10908
rect 4698 10848 4762 10852
rect 4778 10908 4842 10912
rect 4778 10852 4782 10908
rect 4782 10852 4838 10908
rect 4838 10852 4842 10908
rect 4778 10848 4842 10852
rect 4858 10908 4922 10912
rect 4858 10852 4862 10908
rect 4862 10852 4918 10908
rect 4918 10852 4922 10908
rect 4858 10848 4922 10852
rect 11952 10908 12016 10912
rect 11952 10852 11956 10908
rect 11956 10852 12012 10908
rect 12012 10852 12016 10908
rect 11952 10848 12016 10852
rect 12032 10908 12096 10912
rect 12032 10852 12036 10908
rect 12036 10852 12092 10908
rect 12092 10852 12096 10908
rect 12032 10848 12096 10852
rect 12112 10908 12176 10912
rect 12112 10852 12116 10908
rect 12116 10852 12172 10908
rect 12172 10852 12176 10908
rect 12112 10848 12176 10852
rect 12192 10908 12256 10912
rect 12192 10852 12196 10908
rect 12196 10852 12252 10908
rect 12252 10852 12256 10908
rect 12192 10848 12256 10852
rect 19285 10908 19349 10912
rect 19285 10852 19289 10908
rect 19289 10852 19345 10908
rect 19345 10852 19349 10908
rect 19285 10848 19349 10852
rect 19365 10908 19429 10912
rect 19365 10852 19369 10908
rect 19369 10852 19425 10908
rect 19425 10852 19429 10908
rect 19365 10848 19429 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 13492 10780 13556 10844
rect 8285 10364 8349 10368
rect 8285 10308 8289 10364
rect 8289 10308 8345 10364
rect 8345 10308 8349 10364
rect 8285 10304 8349 10308
rect 8365 10364 8429 10368
rect 8365 10308 8369 10364
rect 8369 10308 8425 10364
rect 8425 10308 8429 10364
rect 8365 10304 8429 10308
rect 8445 10364 8509 10368
rect 8445 10308 8449 10364
rect 8449 10308 8505 10364
rect 8505 10308 8509 10364
rect 8445 10304 8509 10308
rect 8525 10364 8589 10368
rect 8525 10308 8529 10364
rect 8529 10308 8585 10364
rect 8585 10308 8589 10364
rect 8525 10304 8589 10308
rect 15618 10364 15682 10368
rect 15618 10308 15622 10364
rect 15622 10308 15678 10364
rect 15678 10308 15682 10364
rect 15618 10304 15682 10308
rect 15698 10364 15762 10368
rect 15698 10308 15702 10364
rect 15702 10308 15758 10364
rect 15758 10308 15762 10364
rect 15698 10304 15762 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 11284 10100 11348 10164
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 4698 9820 4762 9824
rect 4698 9764 4702 9820
rect 4702 9764 4758 9820
rect 4758 9764 4762 9820
rect 4698 9760 4762 9764
rect 4778 9820 4842 9824
rect 4778 9764 4782 9820
rect 4782 9764 4838 9820
rect 4838 9764 4842 9820
rect 4778 9760 4842 9764
rect 4858 9820 4922 9824
rect 4858 9764 4862 9820
rect 4862 9764 4918 9820
rect 4918 9764 4922 9820
rect 4858 9760 4922 9764
rect 11952 9820 12016 9824
rect 11952 9764 11956 9820
rect 11956 9764 12012 9820
rect 12012 9764 12016 9820
rect 11952 9760 12016 9764
rect 12032 9820 12096 9824
rect 12032 9764 12036 9820
rect 12036 9764 12092 9820
rect 12092 9764 12096 9820
rect 12032 9760 12096 9764
rect 12112 9820 12176 9824
rect 12112 9764 12116 9820
rect 12116 9764 12172 9820
rect 12172 9764 12176 9820
rect 12112 9760 12176 9764
rect 12192 9820 12256 9824
rect 12192 9764 12196 9820
rect 12196 9764 12252 9820
rect 12252 9764 12256 9820
rect 12192 9760 12256 9764
rect 19285 9820 19349 9824
rect 19285 9764 19289 9820
rect 19289 9764 19345 9820
rect 19345 9764 19349 9820
rect 19285 9760 19349 9764
rect 19365 9820 19429 9824
rect 19365 9764 19369 9820
rect 19369 9764 19425 9820
rect 19425 9764 19429 9820
rect 19365 9760 19429 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 7604 9692 7668 9756
rect 9628 9556 9692 9620
rect 18828 9556 18892 9620
rect 8285 9276 8349 9280
rect 8285 9220 8289 9276
rect 8289 9220 8345 9276
rect 8345 9220 8349 9276
rect 8285 9216 8349 9220
rect 8365 9276 8429 9280
rect 8365 9220 8369 9276
rect 8369 9220 8425 9276
rect 8425 9220 8429 9276
rect 8365 9216 8429 9220
rect 8445 9276 8509 9280
rect 8445 9220 8449 9276
rect 8449 9220 8505 9276
rect 8505 9220 8509 9276
rect 8445 9216 8509 9220
rect 8525 9276 8589 9280
rect 8525 9220 8529 9276
rect 8529 9220 8585 9276
rect 8585 9220 8589 9276
rect 8525 9216 8589 9220
rect 15618 9276 15682 9280
rect 15618 9220 15622 9276
rect 15622 9220 15678 9276
rect 15678 9220 15682 9276
rect 15618 9216 15682 9220
rect 15698 9276 15762 9280
rect 15698 9220 15702 9276
rect 15702 9220 15758 9276
rect 15758 9220 15762 9276
rect 15698 9216 15762 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 9996 8876 10060 8940
rect 16804 8876 16868 8940
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 4698 8732 4762 8736
rect 4698 8676 4702 8732
rect 4702 8676 4758 8732
rect 4758 8676 4762 8732
rect 4698 8672 4762 8676
rect 4778 8732 4842 8736
rect 4778 8676 4782 8732
rect 4782 8676 4838 8732
rect 4838 8676 4842 8732
rect 4778 8672 4842 8676
rect 4858 8732 4922 8736
rect 4858 8676 4862 8732
rect 4862 8676 4918 8732
rect 4918 8676 4922 8732
rect 4858 8672 4922 8676
rect 11952 8732 12016 8736
rect 11952 8676 11956 8732
rect 11956 8676 12012 8732
rect 12012 8676 12016 8732
rect 11952 8672 12016 8676
rect 12032 8732 12096 8736
rect 12032 8676 12036 8732
rect 12036 8676 12092 8732
rect 12092 8676 12096 8732
rect 12032 8672 12096 8676
rect 12112 8732 12176 8736
rect 12112 8676 12116 8732
rect 12116 8676 12172 8732
rect 12172 8676 12176 8732
rect 12112 8672 12176 8676
rect 12192 8732 12256 8736
rect 12192 8676 12196 8732
rect 12196 8676 12252 8732
rect 12252 8676 12256 8732
rect 12192 8672 12256 8676
rect 19285 8732 19349 8736
rect 19285 8676 19289 8732
rect 19289 8676 19345 8732
rect 19345 8676 19349 8732
rect 19285 8672 19349 8676
rect 19365 8732 19429 8736
rect 19365 8676 19369 8732
rect 19369 8676 19425 8732
rect 19425 8676 19429 8732
rect 19365 8672 19429 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 8285 8188 8349 8192
rect 8285 8132 8289 8188
rect 8289 8132 8345 8188
rect 8345 8132 8349 8188
rect 8285 8128 8349 8132
rect 8365 8188 8429 8192
rect 8365 8132 8369 8188
rect 8369 8132 8425 8188
rect 8425 8132 8429 8188
rect 8365 8128 8429 8132
rect 8445 8188 8509 8192
rect 8445 8132 8449 8188
rect 8449 8132 8505 8188
rect 8505 8132 8509 8188
rect 8445 8128 8509 8132
rect 8525 8188 8589 8192
rect 8525 8132 8529 8188
rect 8529 8132 8585 8188
rect 8585 8132 8589 8188
rect 8525 8128 8589 8132
rect 15618 8188 15682 8192
rect 15618 8132 15622 8188
rect 15622 8132 15678 8188
rect 15678 8132 15682 8188
rect 15618 8128 15682 8132
rect 15698 8188 15762 8192
rect 15698 8132 15702 8188
rect 15702 8132 15758 8188
rect 15758 8132 15762 8188
rect 15698 8128 15762 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 9076 7924 9140 7988
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 4698 7644 4762 7648
rect 4698 7588 4702 7644
rect 4702 7588 4758 7644
rect 4758 7588 4762 7644
rect 4698 7584 4762 7588
rect 4778 7644 4842 7648
rect 4778 7588 4782 7644
rect 4782 7588 4838 7644
rect 4838 7588 4842 7644
rect 4778 7584 4842 7588
rect 4858 7644 4922 7648
rect 4858 7588 4862 7644
rect 4862 7588 4918 7644
rect 4918 7588 4922 7644
rect 4858 7584 4922 7588
rect 11952 7644 12016 7648
rect 11952 7588 11956 7644
rect 11956 7588 12012 7644
rect 12012 7588 12016 7644
rect 11952 7584 12016 7588
rect 12032 7644 12096 7648
rect 12032 7588 12036 7644
rect 12036 7588 12092 7644
rect 12092 7588 12096 7644
rect 12032 7584 12096 7588
rect 12112 7644 12176 7648
rect 12112 7588 12116 7644
rect 12116 7588 12172 7644
rect 12172 7588 12176 7644
rect 12112 7584 12176 7588
rect 12192 7644 12256 7648
rect 12192 7588 12196 7644
rect 12196 7588 12252 7644
rect 12252 7588 12256 7644
rect 12192 7584 12256 7588
rect 19285 7644 19349 7648
rect 19285 7588 19289 7644
rect 19289 7588 19345 7644
rect 19345 7588 19349 7644
rect 19285 7584 19349 7588
rect 19365 7644 19429 7648
rect 19365 7588 19369 7644
rect 19369 7588 19425 7644
rect 19425 7588 19429 7644
rect 19365 7584 19429 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 8285 7100 8349 7104
rect 8285 7044 8289 7100
rect 8289 7044 8345 7100
rect 8345 7044 8349 7100
rect 8285 7040 8349 7044
rect 8365 7100 8429 7104
rect 8365 7044 8369 7100
rect 8369 7044 8425 7100
rect 8425 7044 8429 7100
rect 8365 7040 8429 7044
rect 8445 7100 8509 7104
rect 8445 7044 8449 7100
rect 8449 7044 8505 7100
rect 8505 7044 8509 7100
rect 8445 7040 8509 7044
rect 8525 7100 8589 7104
rect 8525 7044 8529 7100
rect 8529 7044 8585 7100
rect 8585 7044 8589 7100
rect 8525 7040 8589 7044
rect 15618 7100 15682 7104
rect 15618 7044 15622 7100
rect 15622 7044 15678 7100
rect 15678 7044 15682 7100
rect 15618 7040 15682 7044
rect 15698 7100 15762 7104
rect 15698 7044 15702 7100
rect 15702 7044 15758 7100
rect 15758 7044 15762 7100
rect 15698 7040 15762 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 60 6700 124 6764
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 4698 6556 4762 6560
rect 4698 6500 4702 6556
rect 4702 6500 4758 6556
rect 4758 6500 4762 6556
rect 4698 6496 4762 6500
rect 4778 6556 4842 6560
rect 4778 6500 4782 6556
rect 4782 6500 4838 6556
rect 4838 6500 4842 6556
rect 4778 6496 4842 6500
rect 4858 6556 4922 6560
rect 4858 6500 4862 6556
rect 4862 6500 4918 6556
rect 4918 6500 4922 6556
rect 4858 6496 4922 6500
rect 11952 6556 12016 6560
rect 11952 6500 11956 6556
rect 11956 6500 12012 6556
rect 12012 6500 12016 6556
rect 11952 6496 12016 6500
rect 12032 6556 12096 6560
rect 12032 6500 12036 6556
rect 12036 6500 12092 6556
rect 12092 6500 12096 6556
rect 12032 6496 12096 6500
rect 12112 6556 12176 6560
rect 12112 6500 12116 6556
rect 12116 6500 12172 6556
rect 12172 6500 12176 6556
rect 12112 6496 12176 6500
rect 12192 6556 12256 6560
rect 12192 6500 12196 6556
rect 12196 6500 12252 6556
rect 12252 6500 12256 6556
rect 12192 6496 12256 6500
rect 19285 6556 19349 6560
rect 19285 6500 19289 6556
rect 19289 6500 19345 6556
rect 19345 6500 19349 6556
rect 19285 6496 19349 6500
rect 19365 6556 19429 6560
rect 19365 6500 19369 6556
rect 19369 6500 19425 6556
rect 19425 6500 19429 6556
rect 19365 6496 19429 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 60 6292 124 6356
rect 7972 6292 8036 6356
rect 8285 6012 8349 6016
rect 8285 5956 8289 6012
rect 8289 5956 8345 6012
rect 8345 5956 8349 6012
rect 8285 5952 8349 5956
rect 8365 6012 8429 6016
rect 8365 5956 8369 6012
rect 8369 5956 8425 6012
rect 8425 5956 8429 6012
rect 8365 5952 8429 5956
rect 8445 6012 8509 6016
rect 8445 5956 8449 6012
rect 8449 5956 8505 6012
rect 8505 5956 8509 6012
rect 8445 5952 8509 5956
rect 8525 6012 8589 6016
rect 8525 5956 8529 6012
rect 8529 5956 8585 6012
rect 8585 5956 8589 6012
rect 8525 5952 8589 5956
rect 15618 6012 15682 6016
rect 15618 5956 15622 6012
rect 15622 5956 15678 6012
rect 15678 5956 15682 6012
rect 15618 5952 15682 5956
rect 15698 6012 15762 6016
rect 15698 5956 15702 6012
rect 15702 5956 15758 6012
rect 15758 5956 15762 6012
rect 15698 5952 15762 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 5212 5748 5276 5812
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 4698 5468 4762 5472
rect 4698 5412 4702 5468
rect 4702 5412 4758 5468
rect 4758 5412 4762 5468
rect 4698 5408 4762 5412
rect 4778 5468 4842 5472
rect 4778 5412 4782 5468
rect 4782 5412 4838 5468
rect 4838 5412 4842 5468
rect 4778 5408 4842 5412
rect 4858 5468 4922 5472
rect 4858 5412 4862 5468
rect 4862 5412 4918 5468
rect 4918 5412 4922 5468
rect 4858 5408 4922 5412
rect 11952 5468 12016 5472
rect 11952 5412 11956 5468
rect 11956 5412 12012 5468
rect 12012 5412 12016 5468
rect 11952 5408 12016 5412
rect 12032 5468 12096 5472
rect 12032 5412 12036 5468
rect 12036 5412 12092 5468
rect 12092 5412 12096 5468
rect 12032 5408 12096 5412
rect 12112 5468 12176 5472
rect 12112 5412 12116 5468
rect 12116 5412 12172 5468
rect 12172 5412 12176 5468
rect 12112 5408 12176 5412
rect 12192 5468 12256 5472
rect 12192 5412 12196 5468
rect 12196 5412 12252 5468
rect 12252 5412 12256 5468
rect 12192 5408 12256 5412
rect 19285 5468 19349 5472
rect 19285 5412 19289 5468
rect 19289 5412 19345 5468
rect 19345 5412 19349 5468
rect 19285 5408 19349 5412
rect 19365 5468 19429 5472
rect 19365 5412 19369 5468
rect 19369 5412 19425 5468
rect 19425 5412 19429 5468
rect 19365 5408 19429 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 9260 5204 9324 5268
rect 8285 4924 8349 4928
rect 8285 4868 8289 4924
rect 8289 4868 8345 4924
rect 8345 4868 8349 4924
rect 8285 4864 8349 4868
rect 8365 4924 8429 4928
rect 8365 4868 8369 4924
rect 8369 4868 8425 4924
rect 8425 4868 8429 4924
rect 8365 4864 8429 4868
rect 8445 4924 8509 4928
rect 8445 4868 8449 4924
rect 8449 4868 8505 4924
rect 8505 4868 8509 4924
rect 8445 4864 8509 4868
rect 8525 4924 8589 4928
rect 8525 4868 8529 4924
rect 8529 4868 8585 4924
rect 8585 4868 8589 4924
rect 8525 4864 8589 4868
rect 15618 4924 15682 4928
rect 15618 4868 15622 4924
rect 15622 4868 15678 4924
rect 15678 4868 15682 4924
rect 15618 4864 15682 4868
rect 15698 4924 15762 4928
rect 15698 4868 15702 4924
rect 15702 4868 15758 4924
rect 15758 4868 15762 4924
rect 15698 4864 15762 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 5212 4388 5276 4452
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 4698 4380 4762 4384
rect 4698 4324 4702 4380
rect 4702 4324 4758 4380
rect 4758 4324 4762 4380
rect 4698 4320 4762 4324
rect 4778 4380 4842 4384
rect 4778 4324 4782 4380
rect 4782 4324 4838 4380
rect 4838 4324 4842 4380
rect 4778 4320 4842 4324
rect 4858 4380 4922 4384
rect 4858 4324 4862 4380
rect 4862 4324 4918 4380
rect 4918 4324 4922 4380
rect 4858 4320 4922 4324
rect 11952 4380 12016 4384
rect 11952 4324 11956 4380
rect 11956 4324 12012 4380
rect 12012 4324 12016 4380
rect 11952 4320 12016 4324
rect 12032 4380 12096 4384
rect 12032 4324 12036 4380
rect 12036 4324 12092 4380
rect 12092 4324 12096 4380
rect 12032 4320 12096 4324
rect 12112 4380 12176 4384
rect 12112 4324 12116 4380
rect 12116 4324 12172 4380
rect 12172 4324 12176 4380
rect 12112 4320 12176 4324
rect 12192 4380 12256 4384
rect 12192 4324 12196 4380
rect 12196 4324 12252 4380
rect 12252 4324 12256 4380
rect 12192 4320 12256 4324
rect 19285 4380 19349 4384
rect 19285 4324 19289 4380
rect 19289 4324 19345 4380
rect 19345 4324 19349 4380
rect 19285 4320 19349 4324
rect 19365 4380 19429 4384
rect 19365 4324 19369 4380
rect 19369 4324 19425 4380
rect 19425 4324 19429 4380
rect 19365 4320 19429 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 8285 3836 8349 3840
rect 8285 3780 8289 3836
rect 8289 3780 8345 3836
rect 8345 3780 8349 3836
rect 8285 3776 8349 3780
rect 8365 3836 8429 3840
rect 8365 3780 8369 3836
rect 8369 3780 8425 3836
rect 8425 3780 8429 3836
rect 8365 3776 8429 3780
rect 8445 3836 8509 3840
rect 8445 3780 8449 3836
rect 8449 3780 8505 3836
rect 8505 3780 8509 3836
rect 8445 3776 8509 3780
rect 8525 3836 8589 3840
rect 8525 3780 8529 3836
rect 8529 3780 8585 3836
rect 8585 3780 8589 3836
rect 8525 3776 8589 3780
rect 15618 3836 15682 3840
rect 15618 3780 15622 3836
rect 15622 3780 15678 3836
rect 15678 3780 15682 3836
rect 15618 3776 15682 3780
rect 15698 3836 15762 3840
rect 15698 3780 15702 3836
rect 15702 3780 15758 3836
rect 15758 3780 15762 3836
rect 15698 3776 15762 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 6684 3436 6748 3500
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 4698 3292 4762 3296
rect 4698 3236 4702 3292
rect 4702 3236 4758 3292
rect 4758 3236 4762 3292
rect 4698 3232 4762 3236
rect 4778 3292 4842 3296
rect 4778 3236 4782 3292
rect 4782 3236 4838 3292
rect 4838 3236 4842 3292
rect 4778 3232 4842 3236
rect 4858 3292 4922 3296
rect 4858 3236 4862 3292
rect 4862 3236 4918 3292
rect 4918 3236 4922 3292
rect 4858 3232 4922 3236
rect 11952 3292 12016 3296
rect 11952 3236 11956 3292
rect 11956 3236 12012 3292
rect 12012 3236 12016 3292
rect 11952 3232 12016 3236
rect 12032 3292 12096 3296
rect 12032 3236 12036 3292
rect 12036 3236 12092 3292
rect 12092 3236 12096 3292
rect 12032 3232 12096 3236
rect 12112 3292 12176 3296
rect 12112 3236 12116 3292
rect 12116 3236 12172 3292
rect 12172 3236 12176 3292
rect 12112 3232 12176 3236
rect 12192 3292 12256 3296
rect 12192 3236 12196 3292
rect 12196 3236 12252 3292
rect 12252 3236 12256 3292
rect 12192 3232 12256 3236
rect 19285 3292 19349 3296
rect 19285 3236 19289 3292
rect 19289 3236 19345 3292
rect 19345 3236 19349 3292
rect 19285 3232 19349 3236
rect 19365 3292 19429 3296
rect 19365 3236 19369 3292
rect 19369 3236 19425 3292
rect 19425 3236 19429 3292
rect 19365 3232 19429 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 8285 2748 8349 2752
rect 8285 2692 8289 2748
rect 8289 2692 8345 2748
rect 8345 2692 8349 2748
rect 8285 2688 8349 2692
rect 8365 2748 8429 2752
rect 8365 2692 8369 2748
rect 8369 2692 8425 2748
rect 8425 2692 8429 2748
rect 8365 2688 8429 2692
rect 8445 2748 8509 2752
rect 8445 2692 8449 2748
rect 8449 2692 8505 2748
rect 8505 2692 8509 2748
rect 8445 2688 8509 2692
rect 8525 2748 8589 2752
rect 8525 2692 8529 2748
rect 8529 2692 8585 2748
rect 8585 2692 8589 2748
rect 8525 2688 8589 2692
rect 15618 2748 15682 2752
rect 15618 2692 15622 2748
rect 15622 2692 15678 2748
rect 15678 2692 15682 2748
rect 15618 2688 15682 2692
rect 15698 2748 15762 2752
rect 15698 2692 15702 2748
rect 15702 2692 15758 2748
rect 15758 2692 15762 2748
rect 15698 2688 15762 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 4108 2484 4172 2548
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 4698 2204 4762 2208
rect 4698 2148 4702 2204
rect 4702 2148 4758 2204
rect 4758 2148 4762 2204
rect 4698 2144 4762 2148
rect 4778 2204 4842 2208
rect 4778 2148 4782 2204
rect 4782 2148 4838 2204
rect 4838 2148 4842 2204
rect 4778 2144 4842 2148
rect 4858 2204 4922 2208
rect 4858 2148 4862 2204
rect 4862 2148 4918 2204
rect 4918 2148 4922 2204
rect 4858 2144 4922 2148
rect 11952 2204 12016 2208
rect 11952 2148 11956 2204
rect 11956 2148 12012 2204
rect 12012 2148 12016 2204
rect 11952 2144 12016 2148
rect 12032 2204 12096 2208
rect 12032 2148 12036 2204
rect 12036 2148 12092 2204
rect 12092 2148 12096 2204
rect 12032 2144 12096 2148
rect 12112 2204 12176 2208
rect 12112 2148 12116 2204
rect 12116 2148 12172 2204
rect 12172 2148 12176 2204
rect 12112 2144 12176 2148
rect 12192 2204 12256 2208
rect 12192 2148 12196 2204
rect 12196 2148 12252 2204
rect 12252 2148 12256 2204
rect 12192 2144 12256 2148
rect 19285 2204 19349 2208
rect 19285 2148 19289 2204
rect 19289 2148 19345 2204
rect 19345 2148 19349 2204
rect 19285 2144 19349 2148
rect 19365 2204 19429 2208
rect 19365 2148 19369 2204
rect 19369 2148 19425 2204
rect 19425 2148 19429 2204
rect 19365 2144 19429 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 8708 1396 8772 1460
<< metal4 >>
rect 4610 19616 4931 19632
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4931 19616
rect 4610 18528 4931 19552
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4931 18528
rect 4610 17440 4931 18464
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4931 17440
rect 4610 16352 4931 17376
rect 8277 19072 8597 19632
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 17984 8597 19008
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 7603 16964 7669 16965
rect 7603 16900 7604 16964
rect 7668 16900 7669 16964
rect 7603 16899 7669 16900
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4931 16352
rect 4107 15332 4173 15333
rect 4107 15268 4108 15332
rect 4172 15268 4173 15332
rect 4107 15267 4173 15268
rect 59 13700 125 13701
rect 59 13636 60 13700
rect 124 13636 125 13700
rect 59 13635 125 13636
rect 62 13429 122 13635
rect 59 13428 125 13429
rect 59 13364 60 13428
rect 124 13364 125 13428
rect 59 13363 125 13364
rect 59 6764 125 6765
rect 59 6700 60 6764
rect 124 6700 125 6764
rect 59 6699 125 6700
rect 62 6357 122 6699
rect 59 6356 125 6357
rect 59 6292 60 6356
rect 124 6292 125 6356
rect 59 6291 125 6292
rect 4110 2549 4170 15267
rect 4610 15264 4931 16288
rect 6683 16012 6749 16013
rect 6683 15948 6684 16012
rect 6748 15948 6749 16012
rect 6683 15947 6749 15948
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4931 15264
rect 4610 14176 4931 15200
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4931 14176
rect 4610 13088 4931 14112
rect 5211 13428 5277 13429
rect 5211 13364 5212 13428
rect 5276 13364 5277 13428
rect 5211 13363 5277 13364
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4931 13088
rect 4610 12000 4931 13024
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4931 12000
rect 4610 10912 4931 11936
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4931 10912
rect 4610 9824 4931 10848
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4931 9824
rect 4610 8736 4931 9760
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4931 8736
rect 4610 7648 4931 8672
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4931 7648
rect 4610 6560 4931 7584
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4931 6560
rect 4610 5472 4931 6496
rect 5214 5813 5274 13363
rect 5211 5812 5277 5813
rect 5211 5748 5212 5812
rect 5276 5748 5277 5812
rect 5211 5747 5277 5748
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4931 5472
rect 4610 4384 4931 5408
rect 5214 4453 5274 5747
rect 5211 4452 5277 4453
rect 5211 4388 5212 4452
rect 5276 4388 5277 4452
rect 5211 4387 5277 4388
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4931 4384
rect 4610 3296 4931 4320
rect 6686 3501 6746 15947
rect 7606 9757 7666 16899
rect 8277 16896 8597 17920
rect 11944 19616 12264 19632
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 18528 12264 19552
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 17440 12264 18464
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 9995 16964 10061 16965
rect 9995 16900 9996 16964
rect 10060 16900 10061 16964
rect 9995 16899 10061 16900
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 15808 8597 16832
rect 9443 16828 9509 16829
rect 9443 16764 9444 16828
rect 9508 16764 9509 16828
rect 9443 16763 9509 16764
rect 9075 16556 9141 16557
rect 9075 16492 9076 16556
rect 9140 16492 9141 16556
rect 9075 16491 9141 16492
rect 8707 16284 8773 16285
rect 8707 16220 8708 16284
rect 8772 16220 8773 16284
rect 8707 16219 8773 16220
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 14720 8597 15744
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 7787 14516 7853 14517
rect 7787 14452 7788 14516
rect 7852 14452 7853 14516
rect 7787 14451 7853 14452
rect 7790 13293 7850 14451
rect 8277 13632 8597 14656
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 7971 13564 8037 13565
rect 7971 13500 7972 13564
rect 8036 13500 8037 13564
rect 7971 13499 8037 13500
rect 7787 13292 7853 13293
rect 7787 13228 7788 13292
rect 7852 13228 7853 13292
rect 7787 13227 7853 13228
rect 7603 9756 7669 9757
rect 7603 9692 7604 9756
rect 7668 9692 7669 9756
rect 7603 9691 7669 9692
rect 7974 6357 8034 13499
rect 8277 12544 8597 13568
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 11456 8597 12480
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 10368 8597 11392
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 9280 8597 10304
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 8192 8597 9216
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 7104 8597 8128
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 7971 6356 8037 6357
rect 7971 6292 7972 6356
rect 8036 6292 8037 6356
rect 7971 6291 8037 6292
rect 8277 6016 8597 7040
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 4928 8597 5952
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 3840 8597 4864
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 6683 3500 6749 3501
rect 6683 3436 6684 3500
rect 6748 3436 6749 3500
rect 6683 3435 6749 3436
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4931 3296
rect 4107 2548 4173 2549
rect 4107 2484 4108 2548
rect 4172 2484 4173 2548
rect 4107 2483 4173 2484
rect 4610 2208 4931 3232
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4931 2208
rect 4610 2128 4931 2144
rect 8277 2752 8597 3776
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2128 8597 2688
rect 8710 1461 8770 16219
rect 9078 7989 9138 16491
rect 9259 15332 9325 15333
rect 9259 15268 9260 15332
rect 9324 15268 9325 15332
rect 9259 15267 9325 15268
rect 9075 7988 9141 7989
rect 9075 7924 9076 7988
rect 9140 7924 9141 7988
rect 9075 7923 9141 7924
rect 9262 5269 9322 15267
rect 9446 12205 9506 16763
rect 9627 14516 9693 14517
rect 9627 14452 9628 14516
rect 9692 14452 9693 14516
rect 9627 14451 9693 14452
rect 9443 12204 9509 12205
rect 9443 12140 9444 12204
rect 9508 12140 9509 12204
rect 9443 12139 9509 12140
rect 9630 9621 9690 14451
rect 9627 9620 9693 9621
rect 9627 9556 9628 9620
rect 9692 9556 9693 9620
rect 9627 9555 9693 9556
rect 9998 8941 10058 16899
rect 11944 16352 12264 17376
rect 15610 19072 15930 19632
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 17984 15930 19008
rect 19277 19616 19597 19632
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 18528 19597 19552
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 16803 18052 16869 18053
rect 16803 17988 16804 18052
rect 16868 17988 16869 18052
rect 16803 17987 16869 17988
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 13491 17236 13557 17237
rect 13491 17172 13492 17236
rect 13556 17172 13557 17236
rect 13491 17171 13557 17172
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11283 15876 11349 15877
rect 11283 15812 11284 15876
rect 11348 15812 11349 15876
rect 11283 15811 11349 15812
rect 11286 10165 11346 15811
rect 11944 15264 12264 16288
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11651 14788 11717 14789
rect 11651 14724 11652 14788
rect 11716 14724 11717 14788
rect 11651 14723 11717 14724
rect 11654 13973 11714 14723
rect 11944 14176 12264 15200
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11651 13972 11717 13973
rect 11651 13908 11652 13972
rect 11716 13908 11717 13972
rect 11651 13907 11717 13908
rect 11944 13088 12264 14112
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 12000 12264 13024
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 10912 12264 11936
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11283 10164 11349 10165
rect 11283 10100 11284 10164
rect 11348 10100 11349 10164
rect 11283 10099 11349 10100
rect 11944 9824 12264 10848
rect 13494 10845 13554 17171
rect 15610 16896 15930 17920
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 15808 15930 16832
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 14720 15930 15744
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 13632 15930 14656
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 12544 15930 13568
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 11456 15930 12480
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 13491 10844 13557 10845
rect 13491 10780 13492 10844
rect 13556 10780 13557 10844
rect 13491 10779 13557 10780
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 9995 8940 10061 8941
rect 9995 8876 9996 8940
rect 10060 8876 10061 8940
rect 9995 8875 10061 8876
rect 11944 8736 12264 9760
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 7648 12264 8672
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 6560 12264 7584
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 5472 12264 6496
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 9259 5268 9325 5269
rect 9259 5204 9260 5268
rect 9324 5204 9325 5268
rect 9259 5203 9325 5204
rect 11944 4384 12264 5408
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 3296 12264 4320
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 2208 12264 3232
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2128 12264 2144
rect 15610 10368 15930 11392
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 9280 15930 10304
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 8192 15930 9216
rect 16806 8941 16866 17987
rect 19277 17440 19597 18464
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 16352 19597 17376
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 15264 19597 16288
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 18827 15060 18893 15061
rect 18827 14996 18828 15060
rect 18892 14996 18893 15060
rect 18827 14995 18893 14996
rect 18830 9621 18890 14995
rect 19277 14176 19597 15200
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 13088 19597 14112
rect 21587 13700 21653 13701
rect 21587 13636 21588 13700
rect 21652 13636 21653 13700
rect 21587 13635 21653 13636
rect 21590 13429 21650 13635
rect 21587 13428 21653 13429
rect 21587 13364 21588 13428
rect 21652 13364 21653 13428
rect 21587 13363 21653 13364
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 12000 19597 13024
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 10912 19597 11936
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 9824 19597 10848
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 18827 9620 18893 9621
rect 18827 9556 18828 9620
rect 18892 9556 18893 9620
rect 18827 9555 18893 9556
rect 16803 8940 16869 8941
rect 16803 8876 16804 8940
rect 16868 8876 16869 8940
rect 16803 8875 16869 8876
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 7104 15930 8128
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 6016 15930 7040
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 4928 15930 5952
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 3840 15930 4864
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 2752 15930 3776
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2128 15930 2688
rect 19277 8736 19597 9760
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 7648 19597 8672
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 6560 19597 7584
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 5472 19597 6496
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 4384 19597 5408
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 3296 19597 4320
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 2208 19597 3232
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2128 19597 2144
rect 8707 1460 8773 1461
rect 8707 1396 8708 1460
rect 8772 1396 8773 1460
rect 8707 1395 8773 1396
use scs8hd_nor2_4  _081_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__C tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_12
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _065_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 866 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__C
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _146_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_33
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_40
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 4968 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_44 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_80 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_101
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_97
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_161
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_174
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_200 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_conb_1  _133_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_or3_4  _057_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_69
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_2_82
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_188
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_201 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _042_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_or3_4  _059_
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_83
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_155
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_163
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _063_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_77
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_4  _076_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_170
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_188
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 774 592
use scs8hd_or2_4  _054_
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 682 592
use scs8hd_decap_8  FILLER_4_203
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_or3_4  _061_
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__C
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_21
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use scs8hd_nand2_4  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _098_
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 866 592
use scs8hd_or2_4  _124_
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _106_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_109
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_97
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_nor3_4  _109_
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_124
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _108_
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_140 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 130 592
use scs8hd_or4_4  _068_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_nor3_4  _107_
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_99
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_103
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_120
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 15364 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_14
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_18
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 130 592
use scs8hd_or2_4  _084_
timestamp 1586364061
transform 1 0 12512 0 1 7072
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_198
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_202
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_206
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_11
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_6  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 590 592
use scs8hd_or2_4  _117_
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_101
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_183
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_131
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_202
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_111
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_17
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_67
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 1050 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_103
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_162
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_13
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_153
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 2300 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_101
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_185
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _134_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_90
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_103
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_13
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_133
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 590 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_172
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_184
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_188
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_209
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 314 592
use scs8hd_or3_4  _053_
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_166
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use scs8hd_inv_8  _048_
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__053__C
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_20
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_24
timestamp 1586364061
transform 1 0 3312 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_38
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_209
timestamp 1586364061
transform 1 0 20332 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_34
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _062_
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_157
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 406 592
use scs8hd_conb_1  _138_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_8  _049_
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_57
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_8  _044_
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_157
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_6
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_42
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_68
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _055_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__D
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__D
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_151
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 18124 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_188
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_211
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_77
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_or4_4  _091_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_118
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 774 592
use scs8hd_inv_8  _050_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_conb_1  _137_
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_164
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _136_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_174
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_167
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_176
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 314 592
use scs8hd_conb_1  _139_
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_193
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_181
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_192
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 314 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_198
timestamp 1586364061
transform 1 0 19320 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_203
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_211
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_96
timestamp 1586364061
transform 1 0 9936 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_115
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _141_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_182
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_193
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _140_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_120
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 774 592
use scs8hd_decap_6  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_160
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_164
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_187
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_191
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_211
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_101
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_133
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_137
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_181
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_63
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 590 592
use scs8hd_decap_4  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_116
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_125
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_129
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_133
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_137
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_144
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_148
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_154
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 130 592
<< labels >>
rlabel metal2 s 2594 0 2650 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 3698 0 3754 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 824 480 944 6 address[2]
port 2 nsew default input
rlabel metal3 s 21520 824 22000 944 6 address[3]
port 3 nsew default input
rlabel metal3 s 21520 2592 22000 2712 6 address[4]
port 4 nsew default input
rlabel metal3 s 21520 4496 22000 4616 6 address[5]
port 5 nsew default input
rlabel metal3 s 21520 6264 22000 6384 6 address[6]
port 6 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 846 21520 902 22000 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 2594 21520 2650 22000 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal3 s 21520 8168 22000 8288 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 4434 21520 4490 22000 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 6274 21520 6330 22000 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal3 s 0 2592 480 2712 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 8114 21520 8170 22000 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal3 s 21520 9936 22000 10056 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal3 s 21520 11840 22000 11960 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal2 s 9954 21520 10010 22000 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal2 s 11794 21520 11850 22000 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 13634 21520 13690 22000 6 chany_top_in[1]
port 26 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 15474 21520 15530 22000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 14738 0 14794 480 6 chany_top_in[6]
port 31 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chany_top_in[7]
port 32 nsew default input
rlabel metal3 s 21520 13608 22000 13728 6 chany_top_in[8]
port 33 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal3 s 21520 15512 22000 15632 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal3 s 21520 17280 22000 17400 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal3 s 21520 19184 22000 19304 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 data_in
port 43 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 44 nsew default input
rlabel metal2 s 19154 0 19210 480 6 left_grid_pin_1_
port 45 nsew default tristate
rlabel metal2 s 17314 21520 17370 22000 6 left_grid_pin_5_
port 46 nsew default tristate
rlabel metal2 s 19154 21520 19210 22000 6 left_grid_pin_9_
port 47 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 right_grid_pin_0_
port 48 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 right_grid_pin_10_
port 49 nsew default tristate
rlabel metal2 s 20994 21520 21050 22000 6 right_grid_pin_12_
port 50 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 right_grid_pin_14_
port 51 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 right_grid_pin_2_
port 52 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 right_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 right_grid_pin_6_
port 54 nsew default tristate
rlabel metal3 s 21520 20952 22000 21072 6 right_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 4611 2128 4931 19632 6 vpwr
port 56 nsew default input
rlabel metal4 s 8277 2128 8597 19632 6 vgnd
port 57 nsew default input
<< end >>
