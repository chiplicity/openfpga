version https://git-lfs.github.com/spec/v1
oid sha256:4b6f54141fe07933884e58f0a34b152bc962b4db2b98147b177837c609700b2d
size 36423643
