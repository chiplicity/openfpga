magic
tech sky130A
magscale 1 2
timestamp 1604667829
<< locali >>
rect 12633 13175 12667 13481
rect 21649 12631 21683 12937
rect 8309 11679 8343 11781
rect 23857 10999 23891 11101
rect 6101 10523 6135 10693
<< viali >>
rect 24317 21097 24351 21131
rect 25329 21097 25363 21131
rect 24133 20961 24167 20995
rect 25145 20961 25179 20995
rect 19441 20757 19475 20791
rect 25697 20757 25731 20791
rect 26065 20757 26099 20791
rect 1593 20553 1627 20587
rect 7205 20553 7239 20587
rect 9597 20553 9631 20587
rect 12633 20553 12667 20587
rect 14749 20553 14783 20587
rect 17141 20553 17175 20587
rect 18245 20553 18279 20587
rect 21097 20553 21131 20587
rect 24317 20553 24351 20587
rect 19993 20417 20027 20451
rect 25513 20417 25547 20451
rect 26157 20417 26191 20451
rect 1409 20349 1443 20383
rect 7021 20349 7055 20383
rect 7481 20349 7515 20383
rect 9413 20349 9447 20383
rect 12449 20349 12483 20383
rect 12909 20349 12943 20383
rect 14565 20349 14599 20383
rect 15025 20349 15059 20383
rect 16957 20349 16991 20383
rect 18061 20349 18095 20383
rect 18521 20349 18555 20383
rect 19717 20349 19751 20383
rect 20913 20349 20947 20383
rect 21373 20349 21407 20383
rect 24133 20349 24167 20383
rect 19809 20281 19843 20315
rect 1961 20213 1995 20247
rect 9965 20213 9999 20247
rect 17509 20213 17543 20247
rect 19165 20213 19199 20247
rect 19349 20213 19383 20247
rect 23489 20213 23523 20247
rect 24041 20213 24075 20247
rect 24961 20213 24995 20247
rect 25605 20213 25639 20247
rect 25973 20213 26007 20247
rect 26065 20213 26099 20247
rect 11897 20009 11931 20043
rect 12449 20009 12483 20043
rect 17877 20009 17911 20043
rect 24041 19941 24075 19975
rect 12357 19873 12391 19907
rect 15669 19873 15703 19907
rect 15761 19873 15795 19907
rect 18245 19873 18279 19907
rect 18337 19873 18371 19907
rect 25237 19873 25271 19907
rect 12633 19805 12667 19839
rect 15853 19805 15887 19839
rect 18429 19805 18463 19839
rect 19441 19805 19475 19839
rect 25329 19805 25363 19839
rect 25513 19805 25547 19839
rect 26525 19805 26559 19839
rect 24409 19737 24443 19771
rect 24869 19737 24903 19771
rect 1685 19669 1719 19703
rect 4905 19669 4939 19703
rect 10885 19669 10919 19703
rect 11989 19669 12023 19703
rect 13001 19669 13035 19703
rect 14933 19669 14967 19703
rect 15301 19669 15335 19703
rect 16405 19669 16439 19703
rect 24777 19669 24811 19703
rect 25881 19669 25915 19703
rect 14841 19465 14875 19499
rect 22201 19465 22235 19499
rect 24685 19465 24719 19499
rect 26341 19465 26375 19499
rect 16405 19397 16439 19431
rect 4721 19329 4755 19363
rect 5365 19329 5399 19363
rect 11345 19329 11379 19363
rect 13093 19329 13127 19363
rect 13829 19329 13863 19363
rect 14749 19329 14783 19363
rect 15393 19329 15427 19363
rect 16957 19329 16991 19363
rect 25145 19329 25179 19363
rect 25329 19329 25363 19363
rect 26985 19329 27019 19363
rect 2237 19261 2271 19295
rect 2789 19261 2823 19295
rect 9045 19261 9079 19295
rect 9505 19261 9539 19295
rect 10701 19261 10735 19295
rect 11253 19261 11287 19295
rect 12817 19261 12851 19295
rect 14381 19261 14415 19295
rect 15209 19261 15243 19295
rect 15945 19261 15979 19295
rect 19349 19261 19383 19295
rect 19533 19261 19567 19295
rect 22017 19261 22051 19295
rect 22477 19261 22511 19295
rect 24225 19261 24259 19295
rect 25053 19261 25087 19295
rect 25881 19261 25915 19295
rect 26709 19261 26743 19295
rect 5273 19193 5307 19227
rect 10333 19193 10367 19227
rect 11161 19193 11195 19227
rect 16865 19193 16899 19227
rect 19073 19193 19107 19227
rect 19778 19193 19812 19227
rect 1685 19125 1719 19159
rect 2053 19125 2087 19159
rect 2421 19125 2455 19159
rect 3157 19125 3191 19159
rect 4813 19125 4847 19159
rect 5181 19125 5215 19159
rect 8125 19125 8159 19159
rect 9229 19125 9263 19159
rect 10793 19125 10827 19159
rect 11989 19125 12023 19159
rect 12449 19125 12483 19159
rect 12909 19125 12943 19159
rect 13461 19125 13495 19159
rect 15301 19125 15335 19159
rect 16313 19125 16347 19159
rect 16773 19125 16807 19159
rect 17877 19125 17911 19159
rect 18337 19125 18371 19159
rect 18705 19125 18739 19159
rect 20913 19125 20947 19159
rect 24501 19125 24535 19159
rect 26249 19125 26283 19159
rect 26801 19125 26835 19159
rect 27353 19125 27387 19159
rect 1593 18921 1627 18955
rect 6837 18921 6871 18955
rect 8033 18921 8067 18955
rect 10241 18921 10275 18955
rect 13185 18921 13219 18955
rect 15853 18921 15887 18955
rect 19257 18921 19291 18955
rect 22569 18921 22603 18955
rect 25329 18921 25363 18955
rect 26525 18921 26559 18955
rect 26985 18921 27019 18955
rect 1961 18853 1995 18887
rect 23857 18853 23891 18887
rect 24216 18853 24250 18887
rect 26893 18853 26927 18887
rect 5365 18785 5399 18819
rect 8401 18785 8435 18819
rect 10609 18785 10643 18819
rect 12061 18785 12095 18819
rect 16681 18785 16715 18819
rect 17785 18785 17819 18819
rect 18144 18785 18178 18819
rect 22477 18785 22511 18819
rect 2053 18717 2087 18751
rect 2145 18717 2179 18751
rect 5457 18717 5491 18751
rect 5641 18717 5675 18751
rect 8493 18717 8527 18751
rect 8585 18717 8619 18751
rect 10149 18717 10183 18751
rect 10701 18717 10735 18751
rect 10885 18717 10919 18751
rect 11805 18717 11839 18751
rect 16773 18717 16807 18751
rect 16957 18717 16991 18751
rect 17877 18717 17911 18751
rect 20913 18717 20947 18751
rect 22017 18717 22051 18751
rect 22661 18717 22695 18751
rect 23949 18717 23983 18751
rect 27077 18717 27111 18751
rect 2605 18581 2639 18615
rect 2973 18581 3007 18615
rect 3433 18581 3467 18615
rect 3709 18581 3743 18615
rect 4905 18581 4939 18615
rect 4997 18581 5031 18615
rect 7849 18581 7883 18615
rect 11713 18581 11747 18615
rect 15025 18581 15059 18615
rect 15577 18581 15611 18615
rect 16313 18581 16347 18615
rect 19901 18581 19935 18615
rect 20361 18581 20395 18615
rect 22109 18581 22143 18615
rect 23489 18581 23523 18615
rect 3065 18377 3099 18411
rect 4997 18377 5031 18411
rect 6377 18377 6411 18411
rect 7021 18377 7055 18411
rect 10517 18377 10551 18411
rect 11253 18377 11287 18411
rect 12173 18377 12207 18411
rect 12449 18377 12483 18411
rect 16589 18377 16623 18411
rect 17509 18377 17543 18411
rect 18797 18377 18831 18411
rect 20361 18377 20395 18411
rect 21557 18377 21591 18411
rect 27077 18377 27111 18411
rect 1501 18309 1535 18343
rect 11805 18309 11839 18343
rect 20177 18309 20211 18343
rect 22017 18309 22051 18343
rect 27997 18309 28031 18343
rect 2053 18241 2087 18275
rect 3525 18241 3559 18275
rect 3617 18241 3651 18275
rect 5641 18241 5675 18275
rect 6009 18241 6043 18275
rect 11345 18241 11379 18275
rect 13001 18241 13035 18275
rect 18705 18241 18739 18275
rect 19441 18241 19475 18275
rect 20913 18241 20947 18275
rect 22477 18241 22511 18275
rect 22661 18241 22695 18275
rect 24685 18241 24719 18275
rect 3433 18173 3467 18207
rect 4537 18173 4571 18207
rect 6837 18173 6871 18207
rect 8493 18173 8527 18207
rect 8749 18173 8783 18207
rect 15025 18173 15059 18207
rect 15209 18173 15243 18207
rect 19165 18173 19199 18207
rect 20729 18173 20763 18207
rect 21833 18173 21867 18207
rect 25513 18173 25547 18207
rect 25697 18173 25731 18207
rect 27629 18173 27663 18207
rect 1961 18105 1995 18139
rect 5365 18105 5399 18139
rect 8033 18105 8067 18139
rect 12817 18105 12851 18139
rect 13829 18105 13863 18139
rect 14749 18105 14783 18139
rect 15476 18105 15510 18139
rect 19257 18105 19291 18139
rect 19809 18105 19843 18139
rect 20821 18105 20855 18139
rect 22385 18105 22419 18139
rect 23029 18105 23063 18139
rect 24041 18105 24075 18139
rect 24593 18105 24627 18139
rect 25942 18105 25976 18139
rect 1869 18037 1903 18071
rect 2605 18037 2639 18071
rect 2881 18037 2915 18071
rect 4169 18037 4203 18071
rect 4813 18037 4847 18071
rect 5457 18037 5491 18071
rect 7573 18037 7607 18071
rect 8309 18037 8343 18071
rect 9873 18037 9907 18071
rect 10885 18037 10919 18071
rect 12909 18037 12943 18071
rect 13553 18037 13587 18071
rect 17141 18037 17175 18071
rect 18245 18037 18279 18071
rect 23397 18037 23431 18071
rect 24133 18037 24167 18071
rect 24501 18037 24535 18071
rect 25237 18037 25271 18071
rect 2881 17833 2915 17867
rect 4537 17833 4571 17867
rect 4997 17833 5031 17867
rect 6469 17833 6503 17867
rect 9505 17833 9539 17867
rect 11437 17833 11471 17867
rect 12909 17833 12943 17867
rect 14933 17833 14967 17867
rect 18061 17833 18095 17867
rect 18613 17833 18647 17867
rect 19165 17833 19199 17867
rect 20453 17833 20487 17867
rect 21189 17833 21223 17867
rect 22109 17833 22143 17867
rect 26249 17833 26283 17867
rect 3433 17765 3467 17799
rect 5356 17765 5390 17799
rect 16926 17765 16960 17799
rect 21741 17765 21775 17799
rect 26893 17765 26927 17799
rect 1768 17697 1802 17731
rect 3801 17697 3835 17731
rect 5089 17697 5123 17731
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 10149 17697 10183 17731
rect 11529 17697 11563 17731
rect 11796 17697 11830 17731
rect 16681 17697 16715 17731
rect 19533 17697 19567 17731
rect 22457 17697 22491 17731
rect 24777 17697 24811 17731
rect 25237 17697 25271 17731
rect 26985 17697 27019 17731
rect 1501 17629 1535 17663
rect 4077 17629 4111 17663
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 10241 17629 10275 17663
rect 15301 17629 15335 17663
rect 19625 17629 19659 17663
rect 19717 17629 19751 17663
rect 22201 17629 22235 17663
rect 25329 17629 25363 17663
rect 25513 17629 25547 17663
rect 27169 17629 27203 17663
rect 7941 17561 7975 17595
rect 9689 17561 9723 17595
rect 25973 17561 26007 17595
rect 8033 17493 8067 17527
rect 10701 17493 10735 17527
rect 16313 17493 16347 17527
rect 18981 17493 19015 17527
rect 23581 17493 23615 17527
rect 24133 17493 24167 17527
rect 24869 17493 24903 17527
rect 26525 17493 26559 17527
rect 2973 17289 3007 17323
rect 5457 17289 5491 17323
rect 7573 17289 7607 17323
rect 9413 17289 9447 17323
rect 10517 17289 10551 17323
rect 11529 17289 11563 17323
rect 12173 17289 12207 17323
rect 12449 17289 12483 17323
rect 17141 17289 17175 17323
rect 21373 17289 21407 17323
rect 21833 17289 21867 17323
rect 22845 17289 22879 17323
rect 25881 17289 25915 17323
rect 26433 17289 26467 17323
rect 10057 17221 10091 17255
rect 16773 17221 16807 17255
rect 7021 17153 7055 17187
rect 11069 17153 11103 17187
rect 13093 17153 13127 17187
rect 21741 17153 21775 17187
rect 22385 17153 22419 17187
rect 23397 17153 23431 17187
rect 26893 17153 26927 17187
rect 26985 17153 27019 17187
rect 27813 17153 27847 17187
rect 1593 17085 1627 17119
rect 4077 17085 4111 17119
rect 4344 17085 4378 17119
rect 7941 17085 7975 17119
rect 8033 17085 8067 17119
rect 10333 17085 10367 17119
rect 10885 17085 10919 17119
rect 14657 17085 14691 17119
rect 14841 17085 14875 17119
rect 18429 17085 18463 17119
rect 18613 17085 18647 17119
rect 20637 17085 20671 17119
rect 22201 17085 22235 17119
rect 23949 17085 23983 17119
rect 24205 17085 24239 17119
rect 26801 17085 26835 17119
rect 1860 17017 1894 17051
rect 3617 17017 3651 17051
rect 3985 17017 4019 17051
rect 6101 17017 6135 17051
rect 8300 17017 8334 17051
rect 10977 17017 11011 17051
rect 12909 17017 12943 17051
rect 15086 17017 15120 17051
rect 18858 17017 18892 17051
rect 21005 17017 21039 17051
rect 22293 17017 22327 17051
rect 6561 16949 6595 16983
rect 12817 16949 12851 16983
rect 13461 16949 13495 16983
rect 16221 16949 16255 16983
rect 19993 16949 20027 16983
rect 25329 16949 25363 16983
rect 26341 16949 26375 16983
rect 27445 16949 27479 16983
rect 28181 16949 28215 16983
rect 1685 16745 1719 16779
rect 2053 16745 2087 16779
rect 3157 16745 3191 16779
rect 3525 16745 3559 16779
rect 3801 16745 3835 16779
rect 4445 16745 4479 16779
rect 5641 16745 5675 16779
rect 6469 16745 6503 16779
rect 6929 16745 6963 16779
rect 8033 16745 8067 16779
rect 9965 16745 9999 16779
rect 10425 16745 10459 16779
rect 12909 16745 12943 16779
rect 13093 16745 13127 16779
rect 17325 16745 17359 16779
rect 18613 16745 18647 16779
rect 19625 16745 19659 16779
rect 19993 16745 20027 16779
rect 21557 16745 21591 16779
rect 23029 16745 23063 16779
rect 24041 16745 24075 16779
rect 24409 16745 24443 16779
rect 26525 16745 26559 16779
rect 5917 16677 5951 16711
rect 10876 16677 10910 16711
rect 13461 16677 13495 16711
rect 15761 16677 15795 16711
rect 17233 16677 17267 16711
rect 21189 16677 21223 16711
rect 23673 16677 23707 16711
rect 25329 16677 25363 16711
rect 26985 16677 27019 16711
rect 2145 16609 2179 16643
rect 2697 16609 2731 16643
rect 6837 16609 6871 16643
rect 8401 16609 8435 16643
rect 12633 16609 12667 16643
rect 13553 16609 13587 16643
rect 15669 16609 15703 16643
rect 18981 16609 19015 16643
rect 19073 16609 19107 16643
rect 21916 16609 21950 16643
rect 24777 16609 24811 16643
rect 25237 16609 25271 16643
rect 26893 16609 26927 16643
rect 2237 16541 2271 16575
rect 4537 16541 4571 16575
rect 4721 16541 4755 16575
rect 7113 16541 7147 16575
rect 8493 16541 8527 16575
rect 8677 16541 8711 16575
rect 10609 16541 10643 16575
rect 13737 16541 13771 16575
rect 15853 16541 15887 16575
rect 17417 16541 17451 16575
rect 18429 16541 18463 16575
rect 19165 16541 19199 16575
rect 21649 16541 21683 16575
rect 25421 16541 25455 16575
rect 26249 16541 26283 16575
rect 27169 16541 27203 16575
rect 4077 16473 4111 16507
rect 6377 16473 6411 16507
rect 7573 16473 7607 16507
rect 15301 16473 15335 16507
rect 16865 16473 16899 16507
rect 24869 16473 24903 16507
rect 5273 16405 5307 16439
rect 7941 16405 7975 16439
rect 9045 16405 9079 16439
rect 11989 16405 12023 16439
rect 15025 16405 15059 16439
rect 1593 16201 1627 16235
rect 2697 16201 2731 16235
rect 3065 16201 3099 16235
rect 3157 16201 3191 16235
rect 4537 16201 4571 16235
rect 6285 16201 6319 16235
rect 6561 16201 6595 16235
rect 9873 16201 9907 16235
rect 11069 16201 11103 16235
rect 14197 16201 14231 16235
rect 16405 16201 16439 16235
rect 17233 16201 17267 16235
rect 18245 16201 18279 16235
rect 21281 16201 21315 16235
rect 21833 16201 21867 16235
rect 23489 16201 23523 16235
rect 25053 16201 25087 16235
rect 28089 16201 28123 16235
rect 4261 16133 4295 16167
rect 14749 16133 14783 16167
rect 16957 16133 16991 16167
rect 27537 16133 27571 16167
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 3709 16065 3743 16099
rect 5825 16065 5859 16099
rect 7573 16065 7607 16099
rect 12817 16065 12851 16099
rect 15761 16065 15795 16099
rect 15853 16065 15887 16099
rect 18429 16065 18463 16099
rect 21005 16065 21039 16099
rect 22477 16065 22511 16099
rect 23673 16065 23707 16099
rect 26157 16065 26191 16099
rect 7297 15997 7331 16031
rect 8493 15997 8527 16031
rect 11897 15997 11931 16031
rect 13084 15997 13118 16031
rect 15669 15997 15703 16031
rect 22201 15997 22235 16031
rect 26424 15997 26458 16031
rect 1961 15929 1995 15963
rect 3525 15929 3559 15963
rect 5089 15929 5123 15963
rect 8738 15929 8772 15963
rect 12633 15929 12667 15963
rect 15209 15929 15243 15963
rect 17877 15929 17911 15963
rect 18674 15929 18708 15963
rect 20361 15929 20395 15963
rect 23121 15929 23155 15963
rect 23918 15929 23952 15963
rect 25973 15929 26007 15963
rect 3617 15861 3651 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 5641 15861 5675 15895
rect 6929 15861 6963 15895
rect 7389 15861 7423 15895
rect 8125 15861 8159 15895
rect 10609 15861 10643 15895
rect 11345 15861 11379 15895
rect 12173 15861 12207 15895
rect 15301 15861 15335 15895
rect 19809 15861 19843 15895
rect 21741 15861 21775 15895
rect 22293 15861 22327 15895
rect 25605 15861 25639 15895
rect 1685 15657 1719 15691
rect 4629 15657 4663 15691
rect 6285 15657 6319 15691
rect 7389 15657 7423 15691
rect 7849 15657 7883 15691
rect 8033 15657 8067 15691
rect 9413 15657 9447 15691
rect 10609 15657 10643 15691
rect 13737 15657 13771 15691
rect 14657 15657 14691 15691
rect 15117 15657 15151 15691
rect 16681 15657 16715 15691
rect 17233 15657 17267 15691
rect 18429 15657 18463 15691
rect 21833 15657 21867 15691
rect 23305 15657 23339 15691
rect 24869 15657 24903 15691
rect 26157 15657 26191 15691
rect 26893 15657 26927 15691
rect 2237 15589 2271 15623
rect 6929 15589 6963 15623
rect 10149 15589 10183 15623
rect 15568 15589 15602 15623
rect 18889 15589 18923 15623
rect 24777 15589 24811 15623
rect 2145 15521 2179 15555
rect 2789 15521 2823 15555
rect 4353 15521 4387 15555
rect 4905 15521 4939 15555
rect 5172 15521 5206 15555
rect 8401 15521 8435 15555
rect 12072 15521 12106 15555
rect 18797 15521 18831 15555
rect 22192 15521 22226 15555
rect 25237 15521 25271 15555
rect 2329 15453 2363 15487
rect 3525 15453 3559 15487
rect 8493 15453 8527 15487
rect 8585 15453 8619 15487
rect 10701 15453 10735 15487
rect 10793 15453 10827 15487
rect 11621 15453 11655 15487
rect 11805 15453 11839 15487
rect 15301 15453 15335 15487
rect 18981 15453 19015 15487
rect 19441 15453 19475 15487
rect 21925 15453 21959 15487
rect 25329 15453 25363 15487
rect 25513 15453 25547 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 1777 15385 1811 15419
rect 10241 15385 10275 15419
rect 13185 15385 13219 15419
rect 24225 15385 24259 15419
rect 3249 15317 3283 15351
rect 9045 15317 9079 15351
rect 11345 15317 11379 15351
rect 21465 15317 21499 15351
rect 23949 15317 23983 15351
rect 26525 15317 26559 15351
rect 3157 15113 3191 15147
rect 6653 15113 6687 15147
rect 7389 15113 7423 15147
rect 9689 15113 9723 15147
rect 10793 15113 10827 15147
rect 16221 15113 16255 15147
rect 17785 15113 17819 15147
rect 18613 15113 18647 15147
rect 21741 15113 21775 15147
rect 23397 15113 23431 15147
rect 25697 15113 25731 15147
rect 28089 15113 28123 15147
rect 10333 15045 10367 15079
rect 14381 15045 14415 15079
rect 16405 15045 16439 15079
rect 18889 15045 18923 15079
rect 23673 15045 23707 15079
rect 25973 15045 26007 15079
rect 4261 14977 4295 15011
rect 11345 14977 11379 15011
rect 13001 14977 13035 15011
rect 13461 14977 13495 15011
rect 15485 14977 15519 15011
rect 16957 14977 16991 15011
rect 17417 14977 17451 15011
rect 19073 14977 19107 15011
rect 21281 14977 21315 15011
rect 22201 14977 22235 15011
rect 22385 14977 22419 15011
rect 24225 14977 24259 15011
rect 26157 14977 26191 15011
rect 1777 14909 1811 14943
rect 2044 14909 2078 14943
rect 7665 14909 7699 14943
rect 8309 14909 8343 14943
rect 11161 14909 11195 14943
rect 11897 14909 11931 14943
rect 16865 14909 16899 14943
rect 22109 14909 22143 14943
rect 26424 14909 26458 14943
rect 4528 14841 4562 14875
rect 8554 14841 8588 14875
rect 11253 14841 11287 14875
rect 12817 14841 12851 14875
rect 14013 14841 14047 14875
rect 15301 14841 15335 14875
rect 19340 14841 19374 14875
rect 21649 14841 21683 14875
rect 22753 14841 22787 14875
rect 24041 14841 24075 14875
rect 1685 14773 1719 14807
rect 3801 14773 3835 14807
rect 4169 14773 4203 14807
rect 5641 14773 5675 14807
rect 6193 14773 6227 14807
rect 6837 14773 6871 14807
rect 8033 14773 8067 14807
rect 10701 14773 10735 14807
rect 12173 14773 12207 14807
rect 12449 14773 12483 14807
rect 12909 14773 12943 14807
rect 14657 14773 14691 14807
rect 14841 14773 14875 14807
rect 15209 14773 15243 14807
rect 15853 14773 15887 14807
rect 16773 14773 16807 14807
rect 18061 14773 18095 14807
rect 20453 14773 20487 14807
rect 24133 14773 24167 14807
rect 24961 14773 24995 14807
rect 25237 14773 25271 14807
rect 27537 14773 27571 14807
rect 2881 14569 2915 14603
rect 3801 14569 3835 14603
rect 4721 14569 4755 14603
rect 7941 14569 7975 14603
rect 8033 14569 8067 14603
rect 8401 14569 8435 14603
rect 11529 14569 11563 14603
rect 12173 14569 12207 14603
rect 14749 14569 14783 14603
rect 15577 14569 15611 14603
rect 18429 14569 18463 14603
rect 19717 14569 19751 14603
rect 20361 14569 20395 14603
rect 21373 14569 21407 14603
rect 24409 14569 24443 14603
rect 25421 14569 25455 14603
rect 26249 14569 26283 14603
rect 26985 14569 27019 14603
rect 5702 14501 5736 14535
rect 12541 14501 12575 14535
rect 15117 14501 15151 14535
rect 16672 14501 16706 14535
rect 24501 14501 24535 14535
rect 25145 14501 25179 14535
rect 27629 14501 27663 14535
rect 1501 14433 1535 14467
rect 1768 14433 1802 14467
rect 4077 14433 4111 14467
rect 8493 14433 8527 14467
rect 9505 14433 9539 14467
rect 10416 14433 10450 14467
rect 12889 14433 12923 14467
rect 18797 14433 18831 14467
rect 19625 14433 19659 14467
rect 21824 14433 21858 14467
rect 26893 14433 26927 14467
rect 5457 14365 5491 14399
rect 8677 14365 8711 14399
rect 10149 14365 10183 14399
rect 12633 14365 12667 14399
rect 16405 14365 16439 14399
rect 19901 14365 19935 14399
rect 21557 14365 21591 14399
rect 24593 14365 24627 14399
rect 27169 14365 27203 14399
rect 9045 14297 9079 14331
rect 14013 14297 14047 14331
rect 19165 14297 19199 14331
rect 24041 14297 24075 14331
rect 26525 14297 26559 14331
rect 3433 14229 3467 14263
rect 4261 14229 4295 14263
rect 5181 14229 5215 14263
rect 6837 14229 6871 14263
rect 7389 14229 7423 14263
rect 10057 14229 10091 14263
rect 17785 14229 17819 14263
rect 19257 14229 19291 14263
rect 22937 14229 22971 14263
rect 23857 14229 23891 14263
rect 25789 14229 25823 14263
rect 4169 14025 4203 14059
rect 4721 14025 4755 14059
rect 6653 14025 6687 14059
rect 9229 14025 9263 14059
rect 10701 14025 10735 14059
rect 12173 14025 12207 14059
rect 13553 14025 13587 14059
rect 15025 14025 15059 14059
rect 16773 14025 16807 14059
rect 17877 14025 17911 14059
rect 18705 14025 18739 14059
rect 20085 14025 20119 14059
rect 20269 14025 20303 14059
rect 21833 14025 21867 14059
rect 23489 14025 23523 14059
rect 26709 14025 26743 14059
rect 27905 14025 27939 14059
rect 28273 14025 28307 14059
rect 4997 13957 5031 13991
rect 10793 13957 10827 13991
rect 25789 13957 25823 13991
rect 5825 13889 5859 13923
rect 7389 13889 7423 13923
rect 9689 13889 9723 13923
rect 9873 13889 9907 13923
rect 11345 13889 11379 13923
rect 11805 13889 11839 13923
rect 13001 13889 13035 13923
rect 13829 13889 13863 13923
rect 15577 13889 15611 13923
rect 19257 13889 19291 13923
rect 20821 13889 20855 13923
rect 22477 13889 22511 13923
rect 27537 13889 27571 13923
rect 1685 13821 1719 13855
rect 1869 13821 1903 13855
rect 5641 13821 5675 13855
rect 7205 13821 7239 13855
rect 7849 13821 7883 13855
rect 8309 13821 8343 13855
rect 9137 13821 9171 13855
rect 14841 13821 14875 13855
rect 15485 13821 15519 13855
rect 18521 13821 18555 13855
rect 19717 13821 19751 13855
rect 20729 13821 20763 13855
rect 22845 13821 22879 13855
rect 24041 13821 24075 13855
rect 24409 13821 24443 13855
rect 2136 13753 2170 13787
rect 5549 13753 5583 13787
rect 7297 13753 7331 13787
rect 8769 13753 8803 13787
rect 11161 13753 11195 13787
rect 12817 13753 12851 13787
rect 19073 13753 19107 13787
rect 19165 13753 19199 13787
rect 20637 13753 20671 13787
rect 21741 13753 21775 13787
rect 22293 13753 22327 13787
rect 24654 13753 24688 13787
rect 26433 13753 26467 13787
rect 27261 13753 27295 13787
rect 27353 13753 27387 13787
rect 3249 13685 3283 13719
rect 5181 13685 5215 13719
rect 6285 13685 6319 13719
rect 6837 13685 6871 13719
rect 9597 13685 9631 13719
rect 10333 13685 10367 13719
rect 11253 13685 11287 13719
rect 12449 13685 12483 13719
rect 12909 13685 12943 13719
rect 14013 13685 14047 13719
rect 15393 13685 15427 13719
rect 16497 13685 16531 13719
rect 21281 13685 21315 13719
rect 22201 13685 22235 13719
rect 26893 13685 26927 13719
rect 4813 13481 4847 13515
rect 5273 13481 5307 13515
rect 5917 13481 5951 13515
rect 9321 13481 9355 13515
rect 10333 13481 10367 13515
rect 10701 13481 10735 13515
rect 11161 13481 11195 13515
rect 12633 13481 12667 13515
rect 13093 13481 13127 13515
rect 15761 13481 15795 13515
rect 19349 13481 19383 13515
rect 20269 13481 20303 13515
rect 23213 13481 23247 13515
rect 23765 13481 23799 13515
rect 25329 13481 25363 13515
rect 26341 13481 26375 13515
rect 26893 13481 26927 13515
rect 27629 13481 27663 13515
rect 6285 13413 6319 13447
rect 2513 13345 2547 13379
rect 3525 13345 3559 13379
rect 6736 13345 6770 13379
rect 11529 13345 11563 13379
rect 2605 13277 2639 13311
rect 2789 13277 2823 13311
rect 5365 13277 5399 13311
rect 5457 13277 5491 13311
rect 6469 13277 6503 13311
rect 11621 13277 11655 13311
rect 11713 13277 11747 13311
rect 4905 13209 4939 13243
rect 8769 13209 8803 13243
rect 14749 13413 14783 13447
rect 17408 13413 17442 13447
rect 19625 13413 19659 13447
rect 15669 13345 15703 13379
rect 16313 13345 16347 13379
rect 21445 13345 21479 13379
rect 23949 13345 23983 13379
rect 24216 13345 24250 13379
rect 13185 13277 13219 13311
rect 13369 13277 13403 13311
rect 15853 13277 15887 13311
rect 17141 13277 17175 13311
rect 19809 13277 19843 13311
rect 21189 13277 21223 13311
rect 26985 13277 27019 13311
rect 27169 13277 27203 13311
rect 12725 13209 12759 13243
rect 13737 13209 13771 13243
rect 15301 13209 15335 13243
rect 25973 13209 26007 13243
rect 26525 13209 26559 13243
rect 1869 13141 1903 13175
rect 2145 13141 2179 13175
rect 3157 13141 3191 13175
rect 4261 13141 4295 13175
rect 7849 13141 7883 13175
rect 8401 13141 8435 13175
rect 9965 13141 9999 13175
rect 11069 13141 11103 13175
rect 12541 13141 12575 13175
rect 12633 13141 12667 13175
rect 15025 13141 15059 13175
rect 18521 13141 18555 13175
rect 20729 13141 20763 13175
rect 22569 13141 22603 13175
rect 3985 12937 4019 12971
rect 4997 12937 5031 12971
rect 6009 12937 6043 12971
rect 9413 12937 9447 12971
rect 11253 12937 11287 12971
rect 12449 12937 12483 12971
rect 13461 12937 13495 12971
rect 14841 12937 14875 12971
rect 15025 12937 15059 12971
rect 16037 12937 16071 12971
rect 16865 12937 16899 12971
rect 18613 12937 18647 12971
rect 20361 12937 20395 12971
rect 21649 12937 21683 12971
rect 21741 12937 21775 12971
rect 21925 12937 21959 12971
rect 23029 12937 23063 12971
rect 23397 12937 23431 12971
rect 24869 12937 24903 12971
rect 27353 12937 27387 12971
rect 3065 12869 3099 12903
rect 4537 12869 4571 12903
rect 4905 12869 4939 12903
rect 20269 12869 20303 12903
rect 21373 12869 21407 12903
rect 5549 12801 5583 12835
rect 7941 12801 7975 12835
rect 8309 12801 8343 12835
rect 13093 12801 13127 12835
rect 13921 12801 13955 12835
rect 14197 12801 14231 12835
rect 15485 12801 15519 12835
rect 15669 12801 15703 12835
rect 19165 12801 19199 12835
rect 19625 12801 19659 12835
rect 20821 12801 20855 12835
rect 21005 12801 21039 12835
rect 1685 12733 1719 12767
rect 5365 12733 5399 12767
rect 7665 12733 7699 12767
rect 9781 12733 9815 12767
rect 9873 12733 9907 12767
rect 10129 12733 10163 12767
rect 12817 12733 12851 12767
rect 12909 12733 12943 12767
rect 15393 12733 15427 12767
rect 1952 12665 1986 12699
rect 3617 12665 3651 12699
rect 7113 12665 7147 12699
rect 12265 12665 12299 12699
rect 17877 12665 17911 12699
rect 18981 12665 19015 12699
rect 24133 12869 24167 12903
rect 27077 12869 27111 12903
rect 22477 12801 22511 12835
rect 25053 12801 25087 12835
rect 22293 12733 22327 12767
rect 23949 12733 23983 12767
rect 24501 12733 24535 12767
rect 25320 12733 25354 12767
rect 27537 12733 27571 12767
rect 28089 12733 28123 12767
rect 5457 12597 5491 12631
rect 6469 12597 6503 12631
rect 7297 12597 7331 12631
rect 7757 12597 7791 12631
rect 8677 12597 8711 12631
rect 8861 12597 8895 12631
rect 11897 12597 11931 12631
rect 16497 12597 16531 12631
rect 17233 12597 17267 12631
rect 18521 12597 18555 12631
rect 19073 12597 19107 12631
rect 20729 12597 20763 12631
rect 21649 12597 21683 12631
rect 22385 12597 22419 12631
rect 26433 12597 26467 12631
rect 27721 12597 27755 12631
rect 2789 12393 2823 12427
rect 6561 12393 6595 12427
rect 7205 12393 7239 12427
rect 7573 12393 7607 12427
rect 10149 12393 10183 12427
rect 12725 12393 12759 12427
rect 13277 12393 13311 12427
rect 14565 12393 14599 12427
rect 15577 12393 15611 12427
rect 20729 12393 20763 12427
rect 22293 12393 22327 12427
rect 24317 12393 24351 12427
rect 24685 12393 24719 12427
rect 25881 12393 25915 12427
rect 26525 12393 26559 12427
rect 1961 12325 1995 12359
rect 11590 12325 11624 12359
rect 16773 12325 16807 12359
rect 18144 12325 18178 12359
rect 22845 12325 22879 12359
rect 1409 12257 1443 12291
rect 4804 12257 4838 12291
rect 7665 12257 7699 12291
rect 10057 12257 10091 12291
rect 11253 12257 11287 12291
rect 16681 12257 16715 12291
rect 20913 12257 20947 12291
rect 21180 12257 21214 12291
rect 23765 12257 23799 12291
rect 25237 12257 25271 12291
rect 26893 12257 26927 12291
rect 2329 12189 2363 12223
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 4537 12189 4571 12223
rect 7849 12189 7883 12223
rect 8585 12189 8619 12223
rect 10241 12189 10275 12223
rect 11345 12189 11379 12223
rect 16957 12189 16991 12223
rect 17877 12189 17911 12223
rect 20361 12189 20395 12223
rect 25329 12189 25363 12223
rect 25421 12189 25455 12223
rect 26985 12189 27019 12223
rect 27169 12189 27203 12223
rect 1593 12121 1627 12155
rect 3525 12121 3559 12155
rect 9321 12121 9355 12155
rect 16221 12121 16255 12155
rect 23673 12121 23707 12155
rect 26249 12121 26283 12155
rect 2421 12053 2455 12087
rect 3893 12053 3927 12087
rect 4261 12053 4295 12087
rect 5917 12053 5951 12087
rect 7113 12053 7147 12087
rect 8309 12053 8343 12087
rect 8953 12053 8987 12087
rect 9689 12053 9723 12087
rect 14933 12053 14967 12087
rect 16313 12053 16347 12087
rect 19257 12053 19291 12087
rect 23949 12053 23983 12087
rect 24869 12053 24903 12087
rect 2053 11849 2087 11883
rect 2513 11849 2547 11883
rect 3985 11849 4019 11883
rect 5181 11849 5215 11883
rect 7021 11849 7055 11883
rect 8125 11849 8159 11883
rect 9965 11849 9999 11883
rect 10517 11849 10551 11883
rect 10885 11849 10919 11883
rect 11713 11849 11747 11883
rect 14657 11849 14691 11883
rect 15945 11849 15979 11883
rect 17877 11849 17911 11883
rect 21465 11849 21499 11883
rect 23489 11849 23523 11883
rect 25053 11849 25087 11883
rect 25697 11849 25731 11883
rect 28089 11849 28123 11883
rect 4261 11781 4295 11815
rect 4721 11781 4755 11815
rect 8309 11781 8343 11815
rect 8401 11781 8435 11815
rect 11437 11781 11471 11815
rect 16313 11781 16347 11815
rect 21005 11781 21039 11815
rect 25973 11781 26007 11815
rect 2421 11713 2455 11747
rect 2973 11713 3007 11747
rect 3065 11713 3099 11747
rect 5825 11713 5859 11747
rect 7573 11713 7607 11747
rect 15393 11713 15427 11747
rect 17049 11713 17083 11747
rect 22017 11713 22051 11747
rect 23857 11713 23891 11747
rect 24501 11713 24535 11747
rect 24593 11713 24627 11747
rect 1409 11645 1443 11679
rect 4077 11645 4111 11679
rect 5549 11645 5583 11679
rect 7389 11645 7423 11679
rect 8309 11645 8343 11679
rect 8585 11645 8619 11679
rect 8841 11645 8875 11679
rect 15209 11645 15243 11679
rect 18337 11645 18371 11679
rect 18889 11645 18923 11679
rect 18981 11645 19015 11679
rect 21925 11645 21959 11679
rect 22477 11645 22511 11679
rect 24409 11645 24443 11679
rect 26157 11645 26191 11679
rect 2881 11577 2915 11611
rect 3617 11577 3651 11611
rect 5641 11577 5675 11611
rect 15301 11577 15335 11611
rect 16865 11577 16899 11611
rect 19226 11577 19260 11611
rect 21833 11577 21867 11611
rect 26402 11577 26436 11611
rect 1593 11509 1627 11543
rect 4997 11509 5031 11543
rect 6193 11509 6227 11543
rect 6653 11509 6687 11543
rect 7481 11509 7515 11543
rect 14841 11509 14875 11543
rect 16405 11509 16439 11543
rect 16773 11509 16807 11543
rect 17417 11509 17451 11543
rect 20361 11509 20395 11543
rect 21281 11509 21315 11543
rect 24041 11509 24075 11543
rect 27537 11509 27571 11543
rect 1593 11305 1627 11339
rect 2421 11305 2455 11339
rect 2881 11305 2915 11339
rect 5641 11305 5675 11339
rect 6285 11305 6319 11339
rect 8493 11305 8527 11339
rect 10057 11305 10091 11339
rect 14841 11305 14875 11339
rect 16313 11305 16347 11339
rect 17325 11305 17359 11339
rect 17509 11305 17543 11339
rect 19257 11305 19291 11339
rect 19625 11305 19659 11339
rect 20269 11305 20303 11339
rect 21465 11305 21499 11339
rect 21925 11305 21959 11339
rect 22201 11305 22235 11339
rect 22753 11305 22787 11339
rect 23949 11305 23983 11339
rect 24409 11305 24443 11339
rect 25053 11305 25087 11339
rect 25421 11305 25455 11339
rect 26893 11305 26927 11339
rect 26985 11305 27019 11339
rect 3709 11237 3743 11271
rect 4506 11237 4540 11271
rect 6653 11237 6687 11271
rect 7021 11237 7055 11271
rect 7380 11237 7414 11271
rect 9045 11237 9079 11271
rect 9413 11237 9447 11271
rect 16957 11237 16991 11271
rect 17877 11237 17911 11271
rect 17969 11237 18003 11271
rect 19717 11237 19751 11271
rect 22845 11237 22879 11271
rect 26157 11237 26191 11271
rect 2789 11169 2823 11203
rect 18521 11169 18555 11203
rect 21281 11169 21315 11203
rect 23673 11169 23707 11203
rect 24317 11169 24351 11203
rect 2329 11101 2363 11135
rect 3065 11101 3099 11135
rect 4261 11101 4295 11135
rect 7113 11101 7147 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 16405 11101 16439 11135
rect 16497 11101 16531 11135
rect 18061 11101 18095 11135
rect 19901 11101 19935 11135
rect 22937 11101 22971 11135
rect 23857 11101 23891 11135
rect 24593 11101 24627 11135
rect 27077 11101 27111 11135
rect 9689 11033 9723 11067
rect 15945 11033 15979 11067
rect 18981 11033 19015 11067
rect 22385 11033 22419 11067
rect 26525 11033 26559 11067
rect 21189 10965 21223 10999
rect 23857 10965 23891 10999
rect 3065 10761 3099 10795
rect 3617 10761 3651 10795
rect 5181 10761 5215 10795
rect 6285 10761 6319 10795
rect 7481 10761 7515 10795
rect 8861 10761 8895 10795
rect 15945 10761 15979 10795
rect 16405 10761 16439 10795
rect 17601 10761 17635 10795
rect 18061 10761 18095 10795
rect 19165 10761 19199 10795
rect 19441 10761 19475 10795
rect 21189 10761 21223 10795
rect 22477 10761 22511 10795
rect 23121 10761 23155 10795
rect 23489 10761 23523 10795
rect 27169 10761 27203 10795
rect 27905 10761 27939 10795
rect 6101 10693 6135 10727
rect 9045 10693 9079 10727
rect 17233 10693 17267 10727
rect 21097 10693 21131 10727
rect 26157 10693 26191 10727
rect 2697 10625 2731 10659
rect 4077 10625 4111 10659
rect 4261 10625 4295 10659
rect 5825 10625 5859 10659
rect 3525 10557 3559 10591
rect 4721 10557 4755 10591
rect 5641 10557 5675 10591
rect 8033 10625 8067 10659
rect 9597 10625 9631 10659
rect 18521 10625 18555 10659
rect 18613 10625 18647 10659
rect 20177 10625 20211 10659
rect 21649 10625 21683 10659
rect 21833 10625 21867 10659
rect 23673 10625 23707 10659
rect 26709 10625 26743 10659
rect 27537 10625 27571 10659
rect 7941 10557 7975 10591
rect 9505 10557 9539 10591
rect 18429 10557 18463 10591
rect 19993 10557 20027 10591
rect 20085 10557 20119 10591
rect 26617 10557 26651 10591
rect 1961 10489 1995 10523
rect 2421 10489 2455 10523
rect 3985 10489 4019 10523
rect 6101 10489 6135 10523
rect 7297 10489 7331 10523
rect 7849 10489 7883 10523
rect 9413 10489 9447 10523
rect 23940 10489 23974 10523
rect 25605 10489 25639 10523
rect 25973 10489 26007 10523
rect 26525 10489 26559 10523
rect 2053 10421 2087 10455
rect 2513 10421 2547 10455
rect 5089 10421 5123 10455
rect 5549 10421 5583 10455
rect 6653 10421 6687 10455
rect 8585 10421 8619 10455
rect 10057 10421 10091 10455
rect 10425 10421 10459 10455
rect 16773 10421 16807 10455
rect 19625 10421 19659 10455
rect 20729 10421 20763 10455
rect 21557 10421 21591 10455
rect 25053 10421 25087 10455
rect 2329 10217 2363 10251
rect 2789 10217 2823 10251
rect 3525 10217 3559 10251
rect 5457 10217 5491 10251
rect 7941 10217 7975 10251
rect 8493 10217 8527 10251
rect 9689 10217 9723 10251
rect 10241 10217 10275 10251
rect 17601 10217 17635 10251
rect 18245 10217 18279 10251
rect 18889 10217 18923 10251
rect 19717 10217 19751 10251
rect 20729 10217 20763 10251
rect 21557 10217 21591 10251
rect 22017 10217 22051 10251
rect 22661 10217 22695 10251
rect 23029 10217 23063 10251
rect 23489 10217 23523 10251
rect 26249 10217 26283 10251
rect 27077 10217 27111 10251
rect 27629 10217 27663 10251
rect 4344 10149 4378 10183
rect 9137 10149 9171 10183
rect 18337 10149 18371 10183
rect 19349 10149 19383 10183
rect 21925 10149 21959 10183
rect 23826 10149 23860 10183
rect 2881 10081 2915 10115
rect 6817 10081 6851 10115
rect 20085 10081 20119 10115
rect 21281 10081 21315 10115
rect 23581 10081 23615 10115
rect 26525 10081 26559 10115
rect 1961 10013 1995 10047
rect 2973 10013 3007 10047
rect 3893 10013 3927 10047
rect 4077 10013 4111 10047
rect 6561 10013 6595 10047
rect 18429 10013 18463 10047
rect 22201 10013 22235 10047
rect 17877 9945 17911 9979
rect 2421 9877 2455 9911
rect 6101 9877 6135 9911
rect 6377 9877 6411 9911
rect 24961 9877 24995 9911
rect 26709 9877 26743 9911
rect 1777 9673 1811 9707
rect 3341 9673 3375 9707
rect 3617 9673 3651 9707
rect 21557 9673 21591 9707
rect 23029 9673 23063 9707
rect 26341 9673 26375 9707
rect 1869 9605 1903 9639
rect 2881 9605 2915 9639
rect 7481 9605 7515 9639
rect 8585 9605 8619 9639
rect 17141 9605 17175 9639
rect 18061 9605 18095 9639
rect 19625 9605 19659 9639
rect 21097 9605 21131 9639
rect 23857 9605 23891 9639
rect 26617 9605 26651 9639
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 4261 9537 4295 9571
rect 5825 9537 5859 9571
rect 6193 9537 6227 9571
rect 7941 9537 7975 9571
rect 8033 9537 8067 9571
rect 17417 9537 17451 9571
rect 17785 9537 17819 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 19073 9537 19107 9571
rect 20177 9537 20211 9571
rect 20729 9537 20763 9571
rect 22201 9537 22235 9571
rect 22569 9537 22603 9571
rect 23489 9537 23523 9571
rect 24501 9537 24535 9571
rect 25421 9537 25455 9571
rect 4721 9469 4755 9503
rect 5549 9469 5583 9503
rect 9045 9469 9079 9503
rect 18429 9469 18463 9503
rect 20085 9469 20119 9503
rect 21373 9469 21407 9503
rect 22017 9469 22051 9503
rect 26433 9469 26467 9503
rect 26985 9469 27019 9503
rect 27537 9469 27571 9503
rect 28089 9469 28123 9503
rect 3985 9401 4019 9435
rect 4997 9401 5031 9435
rect 19533 9401 19567 9435
rect 21925 9401 21959 9435
rect 24225 9401 24259 9435
rect 24869 9401 24903 9435
rect 2237 9333 2271 9367
rect 4077 9333 4111 9367
rect 5181 9333 5215 9367
rect 5641 9333 5675 9367
rect 6561 9333 6595 9367
rect 7389 9333 7423 9367
rect 7849 9333 7883 9367
rect 19993 9333 20027 9367
rect 24317 9333 24351 9367
rect 27721 9333 27755 9367
rect 1961 9129 1995 9163
rect 4353 9129 4387 9163
rect 5457 9129 5491 9163
rect 7941 9129 7975 9163
rect 18153 9129 18187 9163
rect 18521 9129 18555 9163
rect 19717 9129 19751 9163
rect 21649 9129 21683 9163
rect 21925 9129 21959 9163
rect 23581 9129 23615 9163
rect 24041 9129 24075 9163
rect 24409 9129 24443 9163
rect 24777 9129 24811 9163
rect 2329 9061 2363 9095
rect 6184 9061 6218 9095
rect 24869 9061 24903 9095
rect 2789 8993 2823 9027
rect 3709 8993 3743 9027
rect 4721 8993 4755 9027
rect 26525 8993 26559 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 4813 8925 4847 8959
rect 4905 8925 4939 8959
rect 5917 8925 5951 8959
rect 24961 8925 24995 8959
rect 2421 8789 2455 8823
rect 5825 8789 5859 8823
rect 7297 8789 7331 8823
rect 8401 8789 8435 8823
rect 26709 8789 26743 8823
rect 1961 8585 1995 8619
rect 3065 8585 3099 8619
rect 6837 8585 6871 8619
rect 24501 8585 24535 8619
rect 24869 8585 24903 8619
rect 25237 8585 25271 8619
rect 25513 8585 25547 8619
rect 27353 8585 27387 8619
rect 27721 8585 27755 8619
rect 3617 8517 3651 8551
rect 5181 8517 5215 8551
rect 6193 8517 6227 8551
rect 8401 8517 8435 8551
rect 26617 8517 26651 8551
rect 26985 8517 27019 8551
rect 1869 8449 1903 8483
rect 2513 8449 2547 8483
rect 3525 8449 3559 8483
rect 4077 8449 4111 8483
rect 4169 8449 4203 8483
rect 5825 8449 5859 8483
rect 7389 8449 7423 8483
rect 7849 8449 7883 8483
rect 8309 8449 8343 8483
rect 8861 8449 8895 8483
rect 8953 8449 8987 8483
rect 2329 8381 2363 8415
rect 3985 8381 4019 8415
rect 4721 8381 4755 8415
rect 5641 8381 5675 8415
rect 7205 8381 7239 8415
rect 25329 8381 25363 8415
rect 25881 8381 25915 8415
rect 26433 8381 26467 8415
rect 27537 8381 27571 8415
rect 28089 8381 28123 8415
rect 2421 8313 2455 8347
rect 5089 8313 5123 8347
rect 5549 8313 5583 8347
rect 7297 8313 7331 8347
rect 6561 8245 6595 8279
rect 8769 8245 8803 8279
rect 1593 8041 1627 8075
rect 2145 8041 2179 8075
rect 2697 8041 2731 8075
rect 3065 8041 3099 8075
rect 3617 8041 3651 8075
rect 4997 8041 5031 8075
rect 5181 8041 5215 8075
rect 5549 8041 5583 8075
rect 5641 8041 5675 8075
rect 6745 8041 6779 8075
rect 25513 8041 25547 8075
rect 4721 7973 4755 8007
rect 1409 7905 1443 7939
rect 2513 7905 2547 7939
rect 4077 7905 4111 7939
rect 6285 7905 6319 7939
rect 7113 7905 7147 7939
rect 25329 7905 25363 7939
rect 26525 7905 26559 7939
rect 5733 7837 5767 7871
rect 7205 7837 7239 7871
rect 7297 7837 7331 7871
rect 4261 7769 4295 7803
rect 6561 7701 6595 7735
rect 8401 7701 8435 7735
rect 26709 7701 26743 7735
rect 2329 7497 2363 7531
rect 2697 7497 2731 7531
rect 3801 7497 3835 7531
rect 4169 7497 4203 7531
rect 4537 7497 4571 7531
rect 5273 7497 5307 7531
rect 5733 7497 5767 7531
rect 6101 7497 6135 7531
rect 25421 7497 25455 7531
rect 27353 7497 27387 7531
rect 1593 7429 1627 7463
rect 4905 7429 4939 7463
rect 27721 7429 27755 7463
rect 2053 7361 2087 7395
rect 3525 7361 3559 7395
rect 1409 7293 1443 7327
rect 2513 7293 2547 7327
rect 3617 7293 3651 7327
rect 4721 7293 4755 7327
rect 26433 7293 26467 7327
rect 26985 7293 27019 7327
rect 27537 7293 27571 7327
rect 28089 7293 28123 7327
rect 3157 7225 3191 7259
rect 7113 7225 7147 7259
rect 6561 7157 6595 7191
rect 7389 7157 7423 7191
rect 26617 7157 26651 7191
rect 3065 6953 3099 6987
rect 3617 6953 3651 6987
rect 5733 6953 5767 6987
rect 6101 6885 6135 6919
rect 1409 6817 1443 6851
rect 2053 6817 2087 6851
rect 2329 6817 2363 6851
rect 2513 6817 2547 6851
rect 4077 6817 4111 6851
rect 4721 6817 4755 6851
rect 4997 6817 5031 6851
rect 6193 6817 6227 6851
rect 26525 6817 26559 6851
rect 6377 6749 6411 6783
rect 1593 6681 1627 6715
rect 2697 6681 2731 6715
rect 4261 6613 4295 6647
rect 26709 6613 26743 6647
rect 4169 6409 4203 6443
rect 5733 6409 5767 6443
rect 6193 6409 6227 6443
rect 26341 6409 26375 6443
rect 26617 6409 26651 6443
rect 27077 6409 27111 6443
rect 1593 6341 1627 6375
rect 2053 6341 2087 6375
rect 3525 6341 3559 6375
rect 3157 6273 3191 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 3617 6205 3651 6239
rect 26433 6205 26467 6239
rect 2329 6069 2363 6103
rect 2697 6069 2731 6103
rect 3801 6069 3835 6103
rect 6561 6069 6595 6103
rect 2329 5865 2363 5899
rect 3157 5865 3191 5899
rect 3617 5865 3651 5899
rect 2053 5797 2087 5831
rect 1409 5729 1443 5763
rect 2513 5729 2547 5763
rect 26525 5729 26559 5763
rect 1593 5593 1627 5627
rect 26709 5593 26743 5627
rect 2697 5525 2731 5559
rect 2053 5321 2087 5355
rect 2513 5321 2547 5355
rect 27353 5321 27387 5355
rect 1409 5117 1443 5151
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 1593 4981 1627 5015
rect 26617 4981 26651 5015
rect 1685 4777 1719 4811
rect 2053 3145 2087 3179
rect 1409 2941 1443 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 1593 2805 1627 2839
rect 26617 2805 26651 2839
rect 6285 2601 6319 2635
rect 8309 2601 8343 2635
rect 6745 2465 6779 2499
rect 7196 2465 7230 2499
rect 6929 2397 6963 2431
<< metal1 >>
rect 3510 23400 3516 23452
rect 3568 23440 3574 23452
rect 11974 23440 11980 23452
rect 3568 23412 11980 23440
rect 3568 23400 3574 23412
rect 11974 23400 11980 23412
rect 12032 23400 12038 23452
rect 3510 22516 3516 22568
rect 3568 22556 3574 22568
rect 7926 22556 7932 22568
rect 3568 22528 7932 22556
rect 3568 22516 3574 22528
rect 7926 22516 7932 22528
rect 7984 22516 7990 22568
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 24305 21131 24363 21137
rect 24305 21097 24317 21131
rect 24351 21097 24363 21131
rect 24305 21091 24363 21097
rect 25317 21131 25375 21137
rect 25317 21097 25329 21131
rect 25363 21128 25375 21131
rect 27154 21128 27160 21140
rect 25363 21100 27160 21128
rect 25363 21097 25375 21100
rect 25317 21091 25375 21097
rect 24320 21060 24348 21091
rect 27154 21088 27160 21100
rect 27212 21088 27218 21140
rect 28994 21060 29000 21072
rect 24320 21032 29000 21060
rect 28994 21020 29000 21032
rect 29052 21020 29058 21072
rect 23842 20952 23848 21004
rect 23900 20992 23906 21004
rect 24121 20995 24179 21001
rect 24121 20992 24133 20995
rect 23900 20964 24133 20992
rect 23900 20952 23906 20964
rect 24121 20961 24133 20964
rect 24167 20961 24179 20995
rect 24121 20955 24179 20961
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20992 25191 20995
rect 25179 20964 26096 20992
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 5718 20788 5724 20800
rect 4120 20760 5724 20788
rect 4120 20748 4126 20760
rect 5718 20748 5724 20760
rect 5776 20748 5782 20800
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 19978 20788 19984 20800
rect 19475 20760 19984 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 19978 20748 19984 20760
rect 20036 20748 20042 20800
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 25130 20788 25136 20800
rect 21508 20760 25136 20788
rect 21508 20748 21514 20760
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 25682 20788 25688 20800
rect 25643 20760 25688 20788
rect 25682 20748 25688 20760
rect 25740 20748 25746 20800
rect 26068 20797 26096 20964
rect 26053 20791 26111 20797
rect 26053 20757 26065 20791
rect 26099 20788 26111 20791
rect 26602 20788 26608 20800
rect 26099 20760 26608 20788
rect 26099 20757 26111 20760
rect 26053 20751 26111 20757
rect 26602 20748 26608 20760
rect 26660 20748 26666 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 992 20556 1593 20584
rect 992 20544 998 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 7193 20587 7251 20593
rect 7193 20553 7205 20587
rect 7239 20584 7251 20587
rect 8202 20584 8208 20596
rect 7239 20556 8208 20584
rect 7239 20553 7251 20556
rect 7193 20547 7251 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9585 20587 9643 20593
rect 9585 20553 9597 20587
rect 9631 20584 9643 20587
rect 10226 20584 10232 20596
rect 9631 20556 10232 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 12621 20587 12679 20593
rect 12621 20553 12633 20587
rect 12667 20584 12679 20587
rect 13998 20584 14004 20596
rect 12667 20556 14004 20584
rect 12667 20553 12679 20556
rect 12621 20547 12679 20553
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 14737 20587 14795 20593
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 15838 20584 15844 20596
rect 14783 20556 15844 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 17129 20587 17187 20593
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17770 20584 17776 20596
rect 17175 20556 17776 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 19610 20584 19616 20596
rect 18279 20556 19616 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 21542 20584 21548 20596
rect 21131 20556 21548 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 24305 20587 24363 20593
rect 24305 20553 24317 20587
rect 24351 20584 24363 20587
rect 25222 20584 25228 20596
rect 24351 20556 25228 20584
rect 24351 20553 24363 20556
rect 24305 20547 24363 20553
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 19978 20448 19984 20460
rect 19939 20420 19984 20448
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20448 25559 20451
rect 25774 20448 25780 20460
rect 25547 20420 25780 20448
rect 25547 20417 25559 20420
rect 25501 20411 25559 20417
rect 25774 20408 25780 20420
rect 25832 20448 25838 20460
rect 26145 20451 26203 20457
rect 26145 20448 26157 20451
rect 25832 20420 26157 20448
rect 25832 20408 25838 20420
rect 26145 20417 26157 20420
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 7009 20383 7067 20389
rect 1443 20352 1992 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1964 20256 1992 20352
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7098 20380 7104 20392
rect 7055 20352 7104 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7098 20340 7104 20352
rect 7156 20380 7162 20392
rect 7469 20383 7527 20389
rect 7469 20380 7481 20383
rect 7156 20352 7481 20380
rect 7156 20340 7162 20352
rect 7469 20349 7481 20352
rect 7515 20349 7527 20383
rect 7469 20343 7527 20349
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 9447 20352 9996 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 9968 20256 9996 20352
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12492 20352 12909 20380
rect 12492 20340 12498 20352
rect 12897 20349 12909 20352
rect 12943 20349 12955 20383
rect 12897 20343 12955 20349
rect 14553 20383 14611 20389
rect 14553 20349 14565 20383
rect 14599 20380 14611 20383
rect 14826 20380 14832 20392
rect 14599 20352 14832 20380
rect 14599 20349 14611 20352
rect 14553 20343 14611 20349
rect 14826 20340 14832 20352
rect 14884 20380 14890 20392
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 14884 20352 15025 20380
rect 14884 20340 14890 20352
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20380 17003 20383
rect 16991 20352 17540 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 17512 20256 17540 20352
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 17644 20352 18061 20380
rect 17644 20340 17650 20352
rect 18049 20349 18061 20352
rect 18095 20380 18107 20383
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18095 20352 18521 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 19705 20383 19763 20389
rect 19705 20380 19717 20383
rect 18509 20343 18567 20349
rect 19168 20352 19717 20380
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 9950 20244 9956 20256
rect 9911 20216 9956 20244
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 17494 20244 17500 20256
rect 17455 20216 17500 20244
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 19168 20253 19196 20352
rect 19705 20349 19717 20352
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 20772 20352 20913 20380
rect 20772 20340 20778 20352
rect 20901 20349 20913 20352
rect 20947 20380 20959 20383
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 20947 20352 21373 20380
rect 20947 20349 20959 20352
rect 20901 20343 20959 20349
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 24121 20383 24179 20389
rect 24121 20380 24133 20383
rect 21361 20343 21419 20349
rect 24044 20352 24133 20380
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 19797 20315 19855 20321
rect 19797 20312 19809 20315
rect 19484 20284 19809 20312
rect 19484 20272 19490 20284
rect 19797 20281 19809 20284
rect 19843 20281 19855 20315
rect 19797 20275 19855 20281
rect 24044 20256 24072 20352
rect 24121 20349 24133 20352
rect 24167 20349 24179 20383
rect 24121 20343 24179 20349
rect 25682 20272 25688 20324
rect 25740 20312 25746 20324
rect 25740 20284 26096 20312
rect 25740 20272 25746 20284
rect 19153 20247 19211 20253
rect 19153 20244 19165 20247
rect 18656 20216 19165 20244
rect 18656 20204 18662 20216
rect 19153 20213 19165 20216
rect 19199 20213 19211 20247
rect 19334 20244 19340 20256
rect 19295 20216 19340 20244
rect 19153 20207 19211 20213
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 23477 20247 23535 20253
rect 23477 20213 23489 20247
rect 23523 20244 23535 20247
rect 23842 20244 23848 20256
rect 23523 20216 23848 20244
rect 23523 20213 23535 20216
rect 23477 20207 23535 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 24026 20244 24032 20256
rect 23987 20216 24032 20244
rect 24026 20204 24032 20216
rect 24084 20204 24090 20256
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 25222 20244 25228 20256
rect 24995 20216 25228 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 25590 20244 25596 20256
rect 25551 20216 25596 20244
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 25866 20204 25872 20256
rect 25924 20244 25930 20256
rect 26068 20253 26096 20284
rect 25961 20247 26019 20253
rect 25961 20244 25973 20247
rect 25924 20216 25973 20244
rect 25924 20204 25930 20216
rect 25961 20213 25973 20216
rect 26007 20213 26019 20247
rect 25961 20207 26019 20213
rect 26053 20247 26111 20253
rect 26053 20213 26065 20247
rect 26099 20244 26111 20247
rect 26142 20244 26148 20256
rect 26099 20216 26148 20244
rect 26099 20213 26111 20216
rect 26053 20207 26111 20213
rect 26142 20204 26148 20216
rect 26200 20204 26206 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 12250 20040 12256 20052
rect 11931 20012 12256 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 12250 20000 12256 20012
rect 12308 20040 12314 20052
rect 12437 20043 12495 20049
rect 12437 20040 12449 20043
rect 12308 20012 12449 20040
rect 12308 20000 12314 20012
rect 12437 20009 12449 20012
rect 12483 20009 12495 20043
rect 12437 20003 12495 20009
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 17552 20012 17877 20040
rect 17552 20000 17558 20012
rect 17865 20009 17877 20012
rect 17911 20009 17923 20043
rect 17865 20003 17923 20009
rect 24029 19975 24087 19981
rect 24029 19941 24041 19975
rect 24075 19972 24087 19975
rect 25590 19972 25596 19984
rect 24075 19944 25596 19972
rect 24075 19941 24087 19944
rect 24029 19935 24087 19941
rect 25590 19932 25596 19944
rect 25648 19932 25654 19984
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 11940 19876 12357 19904
rect 11940 19864 11946 19876
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 15654 19904 15660 19916
rect 15615 19876 15660 19904
rect 12345 19867 12403 19873
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 15804 19876 15849 19904
rect 15804 19864 15810 19876
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 18012 19876 18245 19904
rect 18012 19864 18018 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18690 19904 18696 19916
rect 18371 19876 18696 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 25222 19904 25228 19916
rect 25183 19876 25228 19904
rect 25222 19864 25228 19876
rect 25280 19864 25286 19916
rect 12618 19836 12624 19848
rect 12579 19808 12624 19836
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 15838 19836 15844 19848
rect 15799 19808 15844 19836
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 18417 19799 18475 19805
rect 18322 19728 18328 19780
rect 18380 19768 18386 19780
rect 18432 19768 18460 19799
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 25317 19839 25375 19845
rect 25317 19805 25329 19839
rect 25363 19805 25375 19839
rect 25317 19799 25375 19805
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 25774 19836 25780 19848
rect 25547 19808 25780 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 18380 19740 18460 19768
rect 24397 19771 24455 19777
rect 18380 19728 18386 19740
rect 24397 19737 24409 19771
rect 24443 19768 24455 19771
rect 24857 19771 24915 19777
rect 24857 19768 24869 19771
rect 24443 19740 24869 19768
rect 24443 19737 24455 19740
rect 24397 19731 24455 19737
rect 24857 19737 24869 19740
rect 24903 19768 24915 19771
rect 25130 19768 25136 19780
rect 24903 19740 25136 19768
rect 24903 19737 24915 19740
rect 24857 19731 24915 19737
rect 25130 19728 25136 19740
rect 25188 19728 25194 19780
rect 1673 19703 1731 19709
rect 1673 19669 1685 19703
rect 1719 19700 1731 19703
rect 1946 19700 1952 19712
rect 1719 19672 1952 19700
rect 1719 19669 1731 19672
rect 1673 19663 1731 19669
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 4893 19703 4951 19709
rect 4893 19669 4905 19703
rect 4939 19700 4951 19703
rect 5074 19700 5080 19712
rect 4939 19672 5080 19700
rect 4939 19669 4951 19672
rect 4893 19663 4951 19669
rect 5074 19660 5080 19672
rect 5132 19660 5138 19712
rect 10873 19703 10931 19709
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 10962 19700 10968 19712
rect 10919 19672 10968 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 11977 19703 12035 19709
rect 11977 19669 11989 19703
rect 12023 19700 12035 19703
rect 12342 19700 12348 19712
rect 12023 19672 12348 19700
rect 12023 19669 12035 19672
rect 11977 19663 12035 19669
rect 12342 19660 12348 19672
rect 12400 19660 12406 19712
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 12989 19703 13047 19709
rect 12989 19700 13001 19703
rect 12860 19672 13001 19700
rect 12860 19660 12866 19672
rect 12989 19669 13001 19672
rect 13035 19669 13047 19703
rect 12989 19663 13047 19669
rect 14921 19703 14979 19709
rect 14921 19669 14933 19703
rect 14967 19700 14979 19703
rect 15102 19700 15108 19712
rect 14967 19672 15108 19700
rect 14967 19669 14979 19672
rect 14921 19663 14979 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 16390 19700 16396 19712
rect 16351 19672 16396 19700
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 24765 19703 24823 19709
rect 24765 19669 24777 19703
rect 24811 19700 24823 19703
rect 24946 19700 24952 19712
rect 24811 19672 24952 19700
rect 24811 19669 24823 19672
rect 24765 19663 24823 19669
rect 24946 19660 24952 19672
rect 25004 19700 25010 19712
rect 25332 19700 25360 19799
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 26510 19836 26516 19848
rect 26471 19808 26516 19836
rect 26510 19796 26516 19808
rect 26568 19796 26574 19848
rect 25866 19700 25872 19712
rect 25004 19672 25360 19700
rect 25827 19672 25872 19700
rect 25004 19660 25010 19672
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 14826 19496 14832 19508
rect 14787 19468 14832 19496
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 22189 19499 22247 19505
rect 22189 19465 22201 19499
rect 22235 19496 22247 19499
rect 23382 19496 23388 19508
rect 22235 19468 23388 19496
rect 22235 19465 22247 19468
rect 22189 19459 22247 19465
rect 23382 19456 23388 19468
rect 23440 19456 23446 19508
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24673 19499 24731 19505
rect 24673 19496 24685 19499
rect 24084 19468 24685 19496
rect 24084 19456 24090 19468
rect 24673 19465 24685 19468
rect 24719 19465 24731 19499
rect 24673 19459 24731 19465
rect 25866 19456 25872 19508
rect 25924 19496 25930 19508
rect 26329 19499 26387 19505
rect 26329 19496 26341 19499
rect 25924 19468 26341 19496
rect 25924 19456 25930 19468
rect 26329 19465 26341 19468
rect 26375 19465 26387 19499
rect 26329 19459 26387 19465
rect 15746 19388 15752 19440
rect 15804 19428 15810 19440
rect 16393 19431 16451 19437
rect 16393 19428 16405 19431
rect 15804 19400 16405 19428
rect 15804 19388 15810 19400
rect 16393 19397 16405 19400
rect 16439 19397 16451 19431
rect 25774 19428 25780 19440
rect 16393 19391 16451 19397
rect 24964 19400 25780 19428
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19360 4767 19363
rect 5350 19360 5356 19372
rect 4755 19332 5356 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 5350 19320 5356 19332
rect 5408 19320 5414 19372
rect 11330 19360 11336 19372
rect 10980 19332 11336 19360
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 2240 19224 2268 19255
rect 2774 19252 2780 19304
rect 2832 19292 2838 19304
rect 9030 19292 9036 19304
rect 2832 19264 2877 19292
rect 8991 19264 9036 19292
rect 2832 19252 2838 19264
rect 9030 19252 9036 19264
rect 9088 19292 9094 19304
rect 9493 19295 9551 19301
rect 9493 19292 9505 19295
rect 9088 19264 9505 19292
rect 9088 19252 9094 19264
rect 9493 19261 9505 19264
rect 9539 19261 9551 19295
rect 9493 19255 9551 19261
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 10980 19292 11008 19332
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 12618 19360 12624 19372
rect 11756 19332 12624 19360
rect 11756 19320 11762 19332
rect 12618 19320 12624 19332
rect 12676 19360 12682 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12676 19332 13093 19360
rect 12676 19320 12682 19332
rect 13081 19329 13093 19332
rect 13127 19360 13139 19363
rect 13817 19363 13875 19369
rect 13817 19360 13829 19363
rect 13127 19332 13829 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13817 19329 13829 19332
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19360 14795 19363
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 14783 19332 15393 19360
rect 14783 19329 14795 19332
rect 14737 19323 14795 19329
rect 15381 19329 15393 19332
rect 15427 19360 15439 19363
rect 16482 19360 16488 19372
rect 15427 19332 16488 19360
rect 15427 19329 15439 19332
rect 15381 19323 15439 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16945 19363 17003 19369
rect 16945 19360 16957 19363
rect 16592 19332 16957 19360
rect 10735 19264 11008 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 11112 19264 11253 19292
rect 11112 19252 11118 19264
rect 11241 19261 11253 19264
rect 11287 19292 11299 19295
rect 12526 19292 12532 19304
rect 11287 19264 12532 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12802 19292 12808 19304
rect 12763 19264 12808 19292
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 14415 19264 15209 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 15197 19261 15209 19264
rect 15243 19292 15255 19295
rect 15286 19292 15292 19304
rect 15243 19264 15292 19292
rect 15243 19261 15255 19264
rect 15197 19255 15255 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15470 19252 15476 19304
rect 15528 19292 15534 19304
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15528 19264 15945 19292
rect 15528 19252 15534 19264
rect 15933 19261 15945 19264
rect 15979 19292 15991 19295
rect 16592 19292 16620 19332
rect 16945 19329 16957 19332
rect 16991 19360 17003 19363
rect 17402 19360 17408 19372
rect 16991 19332 17408 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 24964 19360 24992 19400
rect 25774 19388 25780 19400
rect 25832 19388 25838 19440
rect 25130 19360 25136 19372
rect 24872 19332 24992 19360
rect 25091 19332 25136 19360
rect 15979 19264 16620 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 17736 19264 19349 19292
rect 17736 19252 17742 19264
rect 19337 19261 19349 19264
rect 19383 19292 19395 19295
rect 19521 19295 19579 19301
rect 19521 19292 19533 19295
rect 19383 19264 19533 19292
rect 19383 19261 19395 19264
rect 19337 19255 19395 19261
rect 19521 19261 19533 19264
rect 19567 19261 19579 19295
rect 19521 19255 19579 19261
rect 21818 19252 21824 19304
rect 21876 19292 21882 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21876 19264 22017 19292
rect 21876 19252 21882 19264
rect 22005 19261 22017 19264
rect 22051 19292 22063 19295
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 22051 19264 22477 19292
rect 22051 19261 22063 19264
rect 22005 19255 22063 19261
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 24210 19292 24216 19304
rect 24123 19264 24216 19292
rect 22465 19255 22523 19261
rect 24210 19252 24216 19264
rect 24268 19292 24274 19304
rect 24872 19292 24900 19332
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25314 19360 25320 19372
rect 25275 19332 25320 19360
rect 25314 19320 25320 19332
rect 25372 19320 25378 19372
rect 26973 19363 27031 19369
rect 26973 19329 26985 19363
rect 27019 19360 27031 19363
rect 27338 19360 27344 19372
rect 27019 19332 27344 19360
rect 27019 19329 27031 19332
rect 26973 19323 27031 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 24268 19264 24900 19292
rect 25041 19295 25099 19301
rect 24268 19252 24274 19264
rect 25041 19261 25053 19295
rect 25087 19292 25099 19295
rect 25590 19292 25596 19304
rect 25087 19264 25596 19292
rect 25087 19261 25099 19264
rect 25041 19255 25099 19261
rect 25590 19252 25596 19264
rect 25648 19252 25654 19304
rect 25869 19295 25927 19301
rect 25869 19261 25881 19295
rect 25915 19292 25927 19295
rect 26510 19292 26516 19304
rect 25915 19264 26516 19292
rect 25915 19261 25927 19264
rect 25869 19255 25927 19261
rect 26510 19252 26516 19264
rect 26568 19292 26574 19304
rect 26697 19295 26755 19301
rect 26697 19292 26709 19295
rect 26568 19264 26709 19292
rect 26568 19252 26574 19264
rect 26697 19261 26709 19264
rect 26743 19261 26755 19295
rect 26697 19255 26755 19261
rect 2792 19224 2820 19252
rect 2240 19196 2820 19224
rect 4890 19184 4896 19236
rect 4948 19224 4954 19236
rect 5261 19227 5319 19233
rect 5261 19224 5273 19227
rect 4948 19196 5273 19224
rect 4948 19184 4954 19196
rect 5261 19193 5273 19196
rect 5307 19193 5319 19227
rect 5261 19187 5319 19193
rect 10321 19227 10379 19233
rect 10321 19193 10333 19227
rect 10367 19224 10379 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10367 19196 11161 19224
rect 10367 19193 10379 19196
rect 10321 19187 10379 19193
rect 11149 19193 11161 19196
rect 11195 19224 11207 19227
rect 16850 19224 16856 19236
rect 11195 19196 12480 19224
rect 16811 19196 16856 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 1673 19159 1731 19165
rect 1673 19125 1685 19159
rect 1719 19156 1731 19159
rect 2041 19159 2099 19165
rect 2041 19156 2053 19159
rect 1719 19128 2053 19156
rect 1719 19125 1731 19128
rect 1673 19119 1731 19125
rect 2041 19125 2053 19128
rect 2087 19156 2099 19159
rect 2130 19156 2136 19168
rect 2087 19128 2136 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 2406 19156 2412 19168
rect 2367 19128 2412 19156
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 3142 19156 3148 19168
rect 3103 19128 3148 19156
rect 3142 19116 3148 19128
rect 3200 19116 3206 19168
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5074 19116 5080 19168
rect 5132 19156 5138 19168
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 5132 19128 5181 19156
rect 5132 19116 5138 19128
rect 5169 19125 5181 19128
rect 5215 19125 5227 19159
rect 8110 19156 8116 19168
rect 8071 19128 8116 19156
rect 5169 19119 5227 19125
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 9214 19156 9220 19168
rect 9175 19128 9220 19156
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 10778 19156 10784 19168
rect 10739 19128 10784 19156
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12452 19165 12480 19196
rect 16850 19184 16856 19196
rect 16908 19184 16914 19236
rect 19061 19227 19119 19233
rect 19061 19193 19073 19227
rect 19107 19224 19119 19227
rect 19766 19227 19824 19233
rect 19766 19224 19778 19227
rect 19107 19196 19778 19224
rect 19107 19193 19119 19196
rect 19061 19187 19119 19193
rect 19766 19193 19778 19196
rect 19812 19224 19824 19227
rect 19978 19224 19984 19236
rect 19812 19196 19984 19224
rect 19812 19193 19824 19196
rect 19766 19187 19824 19193
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 11977 19159 12035 19165
rect 11977 19156 11989 19159
rect 11940 19128 11989 19156
rect 11940 19116 11946 19128
rect 11977 19125 11989 19128
rect 12023 19125 12035 19159
rect 11977 19119 12035 19125
rect 12437 19159 12495 19165
rect 12437 19125 12449 19159
rect 12483 19125 12495 19159
rect 12437 19119 12495 19125
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 13354 19156 13360 19168
rect 12943 19128 13360 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13354 19116 13360 19128
rect 13412 19156 13418 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 13412 19128 13461 19156
rect 13412 19116 13418 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 15289 19159 15347 19165
rect 15289 19156 15301 19159
rect 15160 19128 15301 19156
rect 15160 19116 15166 19128
rect 15289 19125 15301 19128
rect 15335 19125 15347 19159
rect 15289 19119 15347 19125
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19156 16359 19159
rect 16758 19156 16764 19168
rect 16347 19128 16764 19156
rect 16347 19125 16359 19128
rect 16301 19119 16359 19125
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 17862 19156 17868 19168
rect 17823 19128 17868 19156
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18322 19156 18328 19168
rect 18283 19128 18328 19156
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 18690 19156 18696 19168
rect 18651 19128 18696 19156
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20496 19128 20913 19156
rect 20496 19116 20502 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 24486 19156 24492 19168
rect 24447 19128 24492 19156
rect 20901 19119 20959 19125
rect 24486 19116 24492 19128
rect 24544 19116 24550 19168
rect 25590 19116 25596 19168
rect 25648 19156 25654 19168
rect 26237 19159 26295 19165
rect 26237 19156 26249 19159
rect 25648 19128 26249 19156
rect 25648 19116 25654 19128
rect 26237 19125 26249 19128
rect 26283 19156 26295 19159
rect 26789 19159 26847 19165
rect 26789 19156 26801 19159
rect 26283 19128 26801 19156
rect 26283 19125 26295 19128
rect 26237 19119 26295 19125
rect 26789 19125 26801 19128
rect 26835 19125 26847 19159
rect 27338 19156 27344 19168
rect 27299 19128 27344 19156
rect 26789 19119 26847 19125
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 3142 18952 3148 18964
rect 1627 18924 3148 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 3142 18912 3148 18924
rect 3200 18912 3206 18964
rect 4798 18912 4804 18964
rect 4856 18952 4862 18964
rect 6822 18952 6828 18964
rect 4856 18924 6828 18952
rect 4856 18912 4862 18924
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 8021 18955 8079 18961
rect 8021 18921 8033 18955
rect 8067 18952 8079 18955
rect 9030 18952 9036 18964
rect 8067 18924 9036 18952
rect 8067 18921 8079 18924
rect 8021 18915 8079 18921
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 10226 18952 10232 18964
rect 10187 18924 10232 18952
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 13173 18955 13231 18961
rect 13173 18952 13185 18955
rect 10928 18924 13185 18952
rect 10928 18912 10934 18924
rect 13096 18896 13124 18924
rect 13173 18921 13185 18924
rect 13219 18921 13231 18955
rect 13173 18915 13231 18921
rect 15746 18912 15752 18964
rect 15804 18952 15810 18964
rect 15841 18955 15899 18961
rect 15841 18952 15853 18955
rect 15804 18924 15853 18952
rect 15804 18912 15810 18924
rect 15841 18921 15853 18924
rect 15887 18921 15899 18955
rect 15841 18915 15899 18921
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 18380 18924 19257 18952
rect 18380 18912 18386 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 22554 18952 22560 18964
rect 22515 18924 22560 18952
rect 19245 18915 19303 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 24486 18912 24492 18964
rect 24544 18952 24550 18964
rect 25314 18952 25320 18964
rect 24544 18924 25320 18952
rect 24544 18912 24550 18924
rect 25314 18912 25320 18924
rect 25372 18912 25378 18964
rect 26326 18912 26332 18964
rect 26384 18952 26390 18964
rect 26513 18955 26571 18961
rect 26513 18952 26525 18955
rect 26384 18924 26525 18952
rect 26384 18912 26390 18924
rect 26513 18921 26525 18924
rect 26559 18921 26571 18955
rect 26970 18952 26976 18964
rect 26931 18924 26976 18952
rect 26513 18915 26571 18921
rect 26970 18912 26976 18924
rect 27028 18912 27034 18964
rect 1946 18884 1952 18896
rect 1907 18856 1952 18884
rect 1946 18844 1952 18856
rect 2004 18884 2010 18896
rect 2682 18884 2688 18896
rect 2004 18856 2688 18884
rect 2004 18844 2010 18856
rect 2682 18844 2688 18856
rect 2740 18844 2746 18896
rect 13078 18844 13084 18896
rect 13136 18844 13142 18896
rect 24210 18893 24216 18896
rect 23845 18887 23903 18893
rect 23845 18853 23857 18887
rect 23891 18884 23903 18887
rect 24204 18884 24216 18893
rect 23891 18856 24216 18884
rect 23891 18853 23903 18856
rect 23845 18847 23903 18853
rect 24204 18847 24216 18856
rect 24210 18844 24216 18847
rect 24268 18844 24274 18896
rect 26881 18887 26939 18893
rect 26881 18853 26893 18887
rect 26927 18884 26939 18887
rect 27062 18884 27068 18896
rect 26927 18856 27068 18884
rect 26927 18853 26939 18856
rect 26881 18847 26939 18853
rect 27062 18844 27068 18856
rect 27120 18844 27126 18896
rect 4706 18776 4712 18828
rect 4764 18816 4770 18828
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 4764 18788 5365 18816
rect 4764 18776 4770 18788
rect 5353 18785 5365 18788
rect 5399 18785 5411 18819
rect 5353 18779 5411 18785
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 8168 18788 8401 18816
rect 8168 18776 8174 18788
rect 8389 18785 8401 18788
rect 8435 18816 8447 18819
rect 9582 18816 9588 18828
rect 8435 18788 9588 18816
rect 8435 18785 8447 18788
rect 8389 18779 8447 18785
rect 9582 18776 9588 18788
rect 9640 18776 9646 18828
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10597 18819 10655 18825
rect 10597 18816 10609 18819
rect 9732 18788 10609 18816
rect 9732 18776 9738 18788
rect 10597 18785 10609 18788
rect 10643 18816 10655 18819
rect 10778 18816 10784 18828
rect 10643 18788 10784 18816
rect 10643 18785 10655 18788
rect 10597 18779 10655 18785
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 12049 18819 12107 18825
rect 12049 18816 12061 18819
rect 11388 18788 12061 18816
rect 11388 18776 11394 18788
rect 12049 18785 12061 18788
rect 12095 18785 12107 18819
rect 12049 18779 12107 18785
rect 16298 18776 16304 18828
rect 16356 18816 16362 18828
rect 18138 18825 18144 18828
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 16356 18788 16681 18816
rect 16356 18776 16362 18788
rect 16669 18785 16681 18788
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 17773 18819 17831 18825
rect 17773 18785 17785 18819
rect 17819 18816 17831 18819
rect 18132 18816 18144 18825
rect 17819 18788 18144 18816
rect 17819 18785 17831 18788
rect 17773 18779 17831 18785
rect 18132 18779 18144 18788
rect 18138 18776 18144 18779
rect 18196 18776 18202 18828
rect 21634 18776 21640 18828
rect 21692 18816 21698 18828
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 21692 18788 22477 18816
rect 21692 18776 21698 18788
rect 22465 18785 22477 18788
rect 22511 18816 22523 18819
rect 23382 18816 23388 18828
rect 22511 18788 23388 18816
rect 22511 18785 22523 18788
rect 22465 18779 22523 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18717 2099 18751
rect 2041 18711 2099 18717
rect 2056 18680 2084 18711
rect 2130 18708 2136 18760
rect 2188 18748 2194 18760
rect 5442 18748 5448 18760
rect 2188 18720 2233 18748
rect 5403 18720 5448 18748
rect 2188 18708 2194 18720
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 5626 18748 5632 18760
rect 5587 18720 5632 18748
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 8481 18751 8539 18757
rect 8481 18748 8493 18751
rect 7852 18720 8493 18748
rect 2056 18652 3464 18680
rect 3436 18624 3464 18652
rect 1578 18572 1584 18624
rect 1636 18612 1642 18624
rect 2593 18615 2651 18621
rect 2593 18612 2605 18615
rect 1636 18584 2605 18612
rect 1636 18572 1642 18584
rect 2593 18581 2605 18584
rect 2639 18581 2651 18615
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2593 18575 2651 18581
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3418 18612 3424 18624
rect 3379 18584 3424 18612
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 3694 18612 3700 18624
rect 3655 18584 3700 18612
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 4890 18612 4896 18624
rect 4851 18584 4896 18612
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 4985 18615 5043 18621
rect 4985 18581 4997 18615
rect 5031 18612 5043 18615
rect 5258 18612 5264 18624
rect 5031 18584 5264 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 7852 18621 7880 18720
rect 8481 18717 8493 18720
rect 8527 18717 8539 18751
rect 8481 18711 8539 18717
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 10137 18751 10195 18757
rect 8628 18720 8673 18748
rect 8628 18708 8634 18720
rect 10137 18717 10149 18751
rect 10183 18748 10195 18751
rect 10686 18748 10692 18760
rect 10183 18720 10692 18748
rect 10183 18717 10195 18720
rect 10137 18711 10195 18717
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 10870 18748 10876 18760
rect 10831 18720 10876 18748
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11790 18748 11796 18760
rect 11751 18720 11796 18748
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18748 17003 18751
rect 17494 18748 17500 18760
rect 16991 18720 17500 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 16776 18680 16804 18711
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17678 18708 17684 18760
rect 17736 18748 17742 18760
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17736 18720 17877 18748
rect 17736 18708 17742 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20772 18720 20913 18748
rect 20772 18708 20778 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18748 22063 18751
rect 22646 18748 22652 18760
rect 22051 18720 22652 18748
rect 22051 18717 22063 18720
rect 22005 18711 22063 18717
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 23934 18748 23940 18760
rect 23895 18720 23940 18748
rect 23934 18708 23940 18720
rect 23992 18708 23998 18760
rect 26326 18708 26332 18760
rect 26384 18748 26390 18760
rect 27065 18751 27123 18757
rect 27065 18748 27077 18751
rect 26384 18720 27077 18748
rect 26384 18708 26390 18720
rect 27065 18717 27077 18720
rect 27111 18748 27123 18751
rect 27338 18748 27344 18760
rect 27111 18720 27344 18748
rect 27111 18717 27123 18720
rect 27065 18711 27123 18717
rect 27338 18708 27344 18720
rect 27396 18708 27402 18760
rect 16724 18652 16804 18680
rect 16724 18640 16730 18652
rect 7837 18615 7895 18621
rect 7837 18612 7849 18615
rect 6972 18584 7849 18612
rect 6972 18572 6978 18584
rect 7837 18581 7849 18584
rect 7883 18581 7895 18615
rect 11698 18612 11704 18624
rect 11659 18584 11704 18612
rect 7837 18575 7895 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 15010 18612 15016 18624
rect 14971 18584 15016 18612
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15565 18615 15623 18621
rect 15565 18581 15577 18615
rect 15611 18612 15623 18615
rect 15746 18612 15752 18624
rect 15611 18584 15752 18612
rect 15611 18581 15623 18584
rect 15565 18575 15623 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 16301 18615 16359 18621
rect 16301 18581 16313 18615
rect 16347 18612 16359 18615
rect 16390 18612 16396 18624
rect 16347 18584 16396 18612
rect 16347 18581 16359 18584
rect 16301 18575 16359 18581
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 19886 18612 19892 18624
rect 19847 18584 19892 18612
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 20349 18615 20407 18621
rect 20349 18612 20361 18615
rect 20036 18584 20361 18612
rect 20036 18572 20042 18584
rect 20349 18581 20361 18584
rect 20395 18581 20407 18615
rect 20349 18575 20407 18581
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 23477 18615 23535 18621
rect 22152 18584 22197 18612
rect 22152 18572 22158 18584
rect 23477 18581 23489 18615
rect 23523 18612 23535 18615
rect 24670 18612 24676 18624
rect 23523 18584 24676 18612
rect 23523 18581 23535 18584
rect 23477 18575 23535 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3053 18411 3111 18417
rect 3053 18408 3065 18411
rect 2832 18380 3065 18408
rect 2832 18368 2838 18380
rect 3053 18377 3065 18380
rect 3099 18377 3111 18411
rect 4982 18408 4988 18420
rect 4895 18380 4988 18408
rect 3053 18371 3111 18377
rect 4982 18368 4988 18380
rect 5040 18408 5046 18420
rect 5442 18408 5448 18420
rect 5040 18380 5448 18408
rect 5040 18368 5046 18380
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 5684 18380 6377 18408
rect 5684 18368 5690 18380
rect 6365 18377 6377 18380
rect 6411 18408 6423 18411
rect 6454 18408 6460 18420
rect 6411 18380 6460 18408
rect 6411 18377 6423 18380
rect 6365 18371 6423 18377
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 6546 18368 6552 18420
rect 6604 18408 6610 18420
rect 7009 18411 7067 18417
rect 7009 18408 7021 18411
rect 6604 18380 7021 18408
rect 6604 18368 6610 18380
rect 7009 18377 7021 18380
rect 7055 18377 7067 18411
rect 7009 18371 7067 18377
rect 10505 18411 10563 18417
rect 10505 18377 10517 18411
rect 10551 18408 10563 18411
rect 10870 18408 10876 18420
rect 10551 18380 10876 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 11241 18411 11299 18417
rect 11241 18377 11253 18411
rect 11287 18408 11299 18411
rect 11330 18408 11336 18420
rect 11287 18380 11336 18408
rect 11287 18377 11299 18380
rect 11241 18371 11299 18377
rect 11330 18368 11336 18380
rect 11388 18408 11394 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 11388 18380 12173 18408
rect 11388 18368 11394 18380
rect 12161 18377 12173 18380
rect 12207 18408 12219 18411
rect 12207 18380 12296 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 1489 18343 1547 18349
rect 1489 18309 1501 18343
rect 1535 18340 1547 18343
rect 3694 18340 3700 18352
rect 1535 18312 3700 18340
rect 1535 18309 1547 18312
rect 1489 18303 1547 18309
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 3528 18281 3556 18312
rect 3694 18300 3700 18312
rect 3752 18300 3758 18352
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 11790 18340 11796 18352
rect 11572 18312 11796 18340
rect 11572 18300 11578 18312
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 12268 18340 12296 18380
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 16574 18408 16580 18420
rect 12492 18380 12537 18408
rect 16535 18380 16580 18408
rect 12492 18368 12498 18380
rect 16574 18368 16580 18380
rect 16632 18368 16638 18420
rect 17494 18408 17500 18420
rect 17455 18380 17500 18408
rect 17494 18368 17500 18380
rect 17552 18408 17558 18420
rect 17770 18408 17776 18420
rect 17552 18380 17776 18408
rect 17552 18368 17558 18380
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 17862 18368 17868 18420
rect 17920 18408 17926 18420
rect 18785 18411 18843 18417
rect 18785 18408 18797 18411
rect 17920 18380 18797 18408
rect 17920 18368 17926 18380
rect 18785 18377 18797 18380
rect 18831 18377 18843 18411
rect 18785 18371 18843 18377
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 20349 18411 20407 18417
rect 20349 18408 20361 18411
rect 19944 18380 20361 18408
rect 19944 18368 19950 18380
rect 20349 18377 20361 18380
rect 20395 18377 20407 18411
rect 20349 18371 20407 18377
rect 21545 18411 21603 18417
rect 21545 18377 21557 18411
rect 21591 18408 21603 18411
rect 22554 18408 22560 18420
rect 21591 18380 22560 18408
rect 21591 18377 21603 18380
rect 21545 18371 21603 18377
rect 22554 18368 22560 18380
rect 22612 18368 22618 18420
rect 25866 18368 25872 18420
rect 25924 18408 25930 18420
rect 27065 18411 27123 18417
rect 27065 18408 27077 18411
rect 25924 18380 27077 18408
rect 25924 18368 25930 18380
rect 27065 18377 27077 18380
rect 27111 18377 27123 18411
rect 27065 18371 27123 18377
rect 12894 18340 12900 18352
rect 12268 18312 12900 18340
rect 12894 18300 12900 18312
rect 12952 18340 12958 18352
rect 20162 18340 20168 18352
rect 12952 18312 13032 18340
rect 20123 18312 20168 18340
rect 12952 18300 12958 18312
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 5626 18272 5632 18284
rect 5539 18244 5632 18272
rect 3605 18235 3663 18241
rect 2958 18204 2964 18216
rect 2056 18176 2964 18204
rect 1578 18096 1584 18148
rect 1636 18136 1642 18148
rect 1949 18139 2007 18145
rect 1949 18136 1961 18139
rect 1636 18108 1961 18136
rect 1636 18096 1642 18108
rect 1949 18105 1961 18108
rect 1995 18105 2007 18139
rect 1949 18099 2007 18105
rect 1670 18028 1676 18080
rect 1728 18068 1734 18080
rect 1857 18071 1915 18077
rect 1857 18068 1869 18071
rect 1728 18040 1869 18068
rect 1728 18028 1734 18040
rect 1857 18037 1869 18040
rect 1903 18068 1915 18071
rect 2056 18068 2084 18176
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3200 18176 3433 18204
rect 3200 18164 3206 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3620 18204 3648 18235
rect 5626 18232 5632 18244
rect 5684 18272 5690 18284
rect 5997 18275 6055 18281
rect 5997 18272 6009 18275
rect 5684 18244 6009 18272
rect 5684 18232 5690 18244
rect 5997 18241 6009 18244
rect 6043 18241 6055 18275
rect 11333 18275 11391 18281
rect 5997 18235 6055 18241
rect 7576 18244 8616 18272
rect 3421 18167 3479 18173
rect 3528 18176 3648 18204
rect 4525 18207 4583 18213
rect 3528 18136 3556 18176
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4706 18204 4712 18216
rect 4571 18176 4712 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 6822 18204 6828 18216
rect 6783 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 5353 18139 5411 18145
rect 5353 18136 5365 18139
rect 2884 18108 3556 18136
rect 4172 18108 5365 18136
rect 2884 18080 2912 18108
rect 4172 18080 4200 18108
rect 5353 18105 5365 18108
rect 5399 18105 5411 18139
rect 5353 18099 5411 18105
rect 2590 18068 2596 18080
rect 1903 18040 2084 18068
rect 2551 18040 2596 18068
rect 1903 18037 1915 18040
rect 1857 18031 1915 18037
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 2866 18068 2872 18080
rect 2827 18040 2872 18068
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 4154 18068 4160 18080
rect 4115 18040 4160 18068
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4798 18068 4804 18080
rect 4759 18040 4804 18068
rect 4798 18028 4804 18040
rect 4856 18068 4862 18080
rect 5445 18071 5503 18077
rect 5445 18068 5457 18071
rect 4856 18040 5457 18068
rect 4856 18028 4862 18040
rect 5445 18037 5457 18040
rect 5491 18037 5503 18071
rect 5445 18031 5503 18037
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7576 18077 7604 18244
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8168 18176 8493 18204
rect 8168 18164 8174 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8588 18204 8616 18244
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 12802 18272 12808 18284
rect 11379 18244 12808 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 13004 18281 13032 18312
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 21726 18300 21732 18352
rect 21784 18340 21790 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21784 18312 22017 18340
rect 21784 18300 21790 18312
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 26970 18300 26976 18352
rect 27028 18340 27034 18352
rect 27985 18343 28043 18349
rect 27985 18340 27997 18343
rect 27028 18312 27997 18340
rect 27028 18300 27034 18312
rect 27985 18309 27997 18312
rect 28031 18309 28043 18343
rect 27985 18303 28043 18309
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18693 18275 18751 18281
rect 18693 18272 18705 18275
rect 18196 18244 18705 18272
rect 18196 18232 18202 18244
rect 18693 18241 18705 18244
rect 18739 18272 18751 18275
rect 19426 18272 19432 18284
rect 18739 18244 19432 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 19978 18232 19984 18284
rect 20036 18272 20042 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20036 18244 20913 18272
rect 20036 18232 20042 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 22462 18272 22468 18284
rect 22423 18244 22468 18272
rect 20901 18235 20959 18241
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 22646 18272 22652 18284
rect 22607 18244 22652 18272
rect 22646 18232 22652 18244
rect 22704 18232 22710 18284
rect 24670 18272 24676 18284
rect 24631 18244 24676 18272
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 8737 18207 8795 18213
rect 8737 18204 8749 18207
rect 8588 18176 8749 18204
rect 8481 18167 8539 18173
rect 8737 18173 8749 18176
rect 8783 18204 8795 18207
rect 9306 18204 9312 18216
rect 8783 18176 9312 18204
rect 8783 18173 8795 18176
rect 8737 18167 8795 18173
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 14918 18164 14924 18216
rect 14976 18204 14982 18216
rect 15013 18207 15071 18213
rect 15013 18204 15025 18207
rect 14976 18176 15025 18204
rect 14976 18164 14982 18176
rect 15013 18173 15025 18176
rect 15059 18204 15071 18207
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15059 18176 15209 18204
rect 15059 18173 15071 18176
rect 15013 18167 15071 18173
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18204 19211 18207
rect 19886 18204 19892 18216
rect 19199 18176 19892 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 20714 18204 20720 18216
rect 20675 18176 20720 18204
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 21634 18164 21640 18216
rect 21692 18204 21698 18216
rect 21821 18207 21879 18213
rect 21821 18204 21833 18207
rect 21692 18176 21833 18204
rect 21692 18164 21698 18176
rect 21821 18173 21833 18176
rect 21867 18173 21879 18207
rect 25501 18207 25559 18213
rect 25501 18204 25513 18207
rect 21821 18167 21879 18173
rect 23952 18176 25513 18204
rect 23952 18148 23980 18176
rect 25501 18173 25513 18176
rect 25547 18204 25559 18207
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 25547 18176 25697 18204
rect 25547 18173 25559 18176
rect 25501 18167 25559 18173
rect 25685 18173 25697 18176
rect 25731 18173 25743 18207
rect 25685 18167 25743 18173
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 27617 18207 27675 18213
rect 27617 18204 27629 18207
rect 27120 18176 27629 18204
rect 27120 18164 27126 18176
rect 27617 18173 27629 18176
rect 27663 18173 27675 18207
rect 27617 18167 27675 18173
rect 8021 18139 8079 18145
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 8570 18136 8576 18148
rect 8067 18108 8576 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 8570 18096 8576 18108
rect 8628 18136 8634 18148
rect 8628 18108 8708 18136
rect 8628 18096 8634 18108
rect 7561 18071 7619 18077
rect 7561 18068 7573 18071
rect 7340 18040 7573 18068
rect 7340 18028 7346 18040
rect 7561 18037 7573 18040
rect 7607 18037 7619 18071
rect 7561 18031 7619 18037
rect 8110 18028 8116 18080
rect 8168 18068 8174 18080
rect 8297 18071 8355 18077
rect 8297 18068 8309 18071
rect 8168 18040 8309 18068
rect 8168 18028 8174 18040
rect 8297 18037 8309 18040
rect 8343 18037 8355 18071
rect 8680 18068 8708 18108
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 12400 18108 12817 18136
rect 12400 18096 12406 18108
rect 12805 18105 12817 18108
rect 12851 18136 12863 18139
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 12851 18108 13829 18136
rect 12851 18105 12863 18108
rect 12805 18099 12863 18105
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 13817 18099 13875 18105
rect 14737 18139 14795 18145
rect 14737 18105 14749 18139
rect 14783 18136 14795 18139
rect 15464 18139 15522 18145
rect 15464 18136 15476 18139
rect 14783 18108 15476 18136
rect 14783 18105 14795 18108
rect 14737 18099 14795 18105
rect 15464 18105 15476 18108
rect 15510 18136 15522 18139
rect 15746 18136 15752 18148
rect 15510 18108 15752 18136
rect 15510 18105 15522 18108
rect 15464 18099 15522 18105
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 19245 18139 19303 18145
rect 19245 18105 19257 18139
rect 19291 18136 19303 18139
rect 19334 18136 19340 18148
rect 19291 18108 19340 18136
rect 19291 18105 19303 18108
rect 19245 18099 19303 18105
rect 19334 18096 19340 18108
rect 19392 18136 19398 18148
rect 19797 18139 19855 18145
rect 19797 18136 19809 18139
rect 19392 18108 19809 18136
rect 19392 18096 19398 18108
rect 19797 18105 19809 18108
rect 19843 18105 19855 18139
rect 19797 18099 19855 18105
rect 20162 18096 20168 18148
rect 20220 18136 20226 18148
rect 20809 18139 20867 18145
rect 20809 18136 20821 18139
rect 20220 18108 20821 18136
rect 20220 18096 20226 18108
rect 20809 18105 20821 18108
rect 20855 18136 20867 18139
rect 21358 18136 21364 18148
rect 20855 18108 21364 18136
rect 20855 18105 20867 18108
rect 20809 18099 20867 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 21910 18096 21916 18148
rect 21968 18136 21974 18148
rect 22373 18139 22431 18145
rect 22373 18136 22385 18139
rect 21968 18108 22385 18136
rect 21968 18096 21974 18108
rect 22373 18105 22385 18108
rect 22419 18136 22431 18139
rect 23017 18139 23075 18145
rect 23017 18136 23029 18139
rect 22419 18108 23029 18136
rect 22419 18105 22431 18108
rect 22373 18099 22431 18105
rect 23017 18105 23029 18108
rect 23063 18105 23075 18139
rect 23934 18136 23940 18148
rect 23017 18099 23075 18105
rect 23400 18108 23940 18136
rect 23400 18080 23428 18108
rect 23934 18096 23940 18108
rect 23992 18096 23998 18148
rect 24029 18139 24087 18145
rect 24029 18105 24041 18139
rect 24075 18136 24087 18139
rect 24210 18136 24216 18148
rect 24075 18108 24216 18136
rect 24075 18105 24087 18108
rect 24029 18099 24087 18105
rect 24210 18096 24216 18108
rect 24268 18136 24274 18148
rect 24581 18139 24639 18145
rect 24581 18136 24593 18139
rect 24268 18108 24593 18136
rect 24268 18096 24274 18108
rect 24581 18105 24593 18108
rect 24627 18105 24639 18139
rect 25930 18139 25988 18145
rect 25930 18136 25942 18139
rect 24581 18099 24639 18105
rect 25332 18108 25942 18136
rect 25332 18080 25360 18108
rect 25930 18105 25942 18108
rect 25976 18136 25988 18139
rect 26234 18136 26240 18148
rect 25976 18108 26240 18136
rect 25976 18105 25988 18108
rect 25930 18099 25988 18105
rect 26234 18096 26240 18108
rect 26292 18096 26298 18148
rect 9861 18071 9919 18077
rect 9861 18068 9873 18071
rect 8680 18040 9873 18068
rect 8297 18031 8355 18037
rect 9861 18037 9873 18040
rect 9907 18068 9919 18071
rect 10134 18068 10140 18080
rect 9907 18040 10140 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10870 18068 10876 18080
rect 10831 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 12897 18071 12955 18077
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 13538 18068 13544 18080
rect 12943 18040 13544 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13630 18028 13636 18080
rect 13688 18068 13694 18080
rect 16666 18068 16672 18080
rect 13688 18040 16672 18068
rect 13688 18028 13694 18040
rect 16666 18028 16672 18040
rect 16724 18068 16730 18080
rect 17129 18071 17187 18077
rect 17129 18068 17141 18071
rect 16724 18040 17141 18068
rect 16724 18028 16730 18040
rect 17129 18037 17141 18040
rect 17175 18037 17187 18071
rect 17129 18031 17187 18037
rect 17678 18028 17684 18080
rect 17736 18068 17742 18080
rect 18233 18071 18291 18077
rect 18233 18068 18245 18071
rect 17736 18040 18245 18068
rect 17736 18028 17742 18040
rect 18233 18037 18245 18040
rect 18279 18037 18291 18071
rect 23382 18068 23388 18080
rect 23343 18040 23388 18068
rect 18233 18031 18291 18037
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 23474 18028 23480 18080
rect 23532 18068 23538 18080
rect 24121 18071 24179 18077
rect 24121 18068 24133 18071
rect 23532 18040 24133 18068
rect 23532 18028 23538 18040
rect 24121 18037 24133 18040
rect 24167 18037 24179 18071
rect 24121 18031 24179 18037
rect 24394 18028 24400 18080
rect 24452 18068 24458 18080
rect 24489 18071 24547 18077
rect 24489 18068 24501 18071
rect 24452 18040 24501 18068
rect 24452 18028 24458 18040
rect 24489 18037 24501 18040
rect 24535 18037 24547 18071
rect 24489 18031 24547 18037
rect 25225 18071 25283 18077
rect 25225 18037 25237 18071
rect 25271 18068 25283 18071
rect 25314 18068 25320 18080
rect 25271 18040 25320 18068
rect 25271 18037 25283 18040
rect 25225 18031 25283 18037
rect 25314 18028 25320 18040
rect 25372 18028 25378 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17864 2930 17876
rect 4338 17864 4344 17876
rect 2924 17836 4344 17864
rect 2924 17824 2930 17836
rect 4338 17824 4344 17836
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 4982 17864 4988 17876
rect 4943 17836 4988 17864
rect 4525 17827 4583 17833
rect 4982 17824 4988 17836
rect 5040 17824 5046 17876
rect 6454 17864 6460 17876
rect 6415 17836 6460 17864
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 9493 17867 9551 17873
rect 9493 17833 9505 17867
rect 9539 17864 9551 17867
rect 9674 17864 9680 17876
rect 9539 17836 9680 17864
rect 9539 17833 9551 17836
rect 9493 17827 9551 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 11425 17867 11483 17873
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 11698 17864 11704 17876
rect 11471 17836 11704 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 11698 17824 11704 17836
rect 11756 17864 11762 17876
rect 12894 17864 12900 17876
rect 11756 17836 11836 17864
rect 12855 17836 12900 17864
rect 11756 17824 11762 17836
rect 2590 17756 2596 17808
rect 2648 17796 2654 17808
rect 3421 17799 3479 17805
rect 3421 17796 3433 17799
rect 2648 17768 3433 17796
rect 2648 17756 2654 17768
rect 3421 17765 3433 17768
rect 3467 17796 3479 17799
rect 3510 17796 3516 17808
rect 3467 17768 3516 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3510 17756 3516 17768
rect 3568 17756 3574 17808
rect 5344 17799 5402 17805
rect 5344 17765 5356 17799
rect 5390 17796 5402 17799
rect 5626 17796 5632 17808
rect 5390 17768 5632 17796
rect 5390 17765 5402 17768
rect 5344 17759 5402 17765
rect 5626 17756 5632 17768
rect 5684 17756 5690 17808
rect 1756 17731 1814 17737
rect 1756 17697 1768 17731
rect 1802 17728 1814 17731
rect 2038 17728 2044 17740
rect 1802 17700 2044 17728
rect 1802 17697 1814 17700
rect 1756 17691 1814 17697
rect 2038 17688 2044 17700
rect 2096 17728 2102 17740
rect 2958 17728 2964 17740
rect 2096 17700 2964 17728
rect 2096 17688 2102 17700
rect 2958 17688 2964 17700
rect 3016 17728 3022 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 3016 17700 3801 17728
rect 3016 17688 3022 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17728 5135 17731
rect 5166 17728 5172 17740
rect 5123 17700 5172 17728
rect 5123 17697 5135 17700
rect 5077 17691 5135 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 7926 17688 7932 17740
rect 7984 17728 7990 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7984 17700 8401 17728
rect 7984 17688 7990 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 10042 17728 10048 17740
rect 10003 17700 10048 17728
rect 8389 17691 8447 17697
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10318 17728 10324 17740
rect 10183 17700 10324 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 11514 17728 11520 17740
rect 11475 17700 11520 17728
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11808 17737 11836 17836
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 14921 17867 14979 17873
rect 14921 17833 14933 17867
rect 14967 17864 14979 17867
rect 15010 17864 15016 17876
rect 14967 17836 15016 17864
rect 14967 17833 14979 17836
rect 14921 17827 14979 17833
rect 15010 17824 15016 17836
rect 15068 17864 15074 17876
rect 15470 17864 15476 17876
rect 15068 17836 15476 17864
rect 15068 17824 15074 17836
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 18012 17836 18061 17864
rect 18012 17824 18018 17836
rect 18049 17833 18061 17836
rect 18095 17864 18107 17867
rect 18506 17864 18512 17876
rect 18095 17836 18512 17864
rect 18095 17833 18107 17836
rect 18049 17827 18107 17833
rect 18506 17824 18512 17836
rect 18564 17864 18570 17876
rect 18601 17867 18659 17873
rect 18601 17864 18613 17867
rect 18564 17836 18613 17864
rect 18564 17824 18570 17836
rect 18601 17833 18613 17836
rect 18647 17833 18659 17867
rect 18601 17827 18659 17833
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 19153 17867 19211 17873
rect 19153 17864 19165 17867
rect 18748 17836 19165 17864
rect 18748 17824 18754 17836
rect 19153 17833 19165 17836
rect 19199 17833 19211 17867
rect 19153 17827 19211 17833
rect 20441 17867 20499 17873
rect 20441 17833 20453 17867
rect 20487 17864 20499 17867
rect 20622 17864 20628 17876
rect 20487 17836 20628 17864
rect 20487 17833 20499 17836
rect 20441 17827 20499 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 21177 17867 21235 17873
rect 21177 17833 21189 17867
rect 21223 17864 21235 17867
rect 21910 17864 21916 17876
rect 21223 17836 21916 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 22097 17867 22155 17873
rect 22097 17833 22109 17867
rect 22143 17864 22155 17867
rect 22278 17864 22284 17876
rect 22143 17836 22284 17864
rect 22143 17833 22155 17836
rect 22097 17827 22155 17833
rect 22278 17824 22284 17836
rect 22336 17864 22342 17876
rect 22462 17864 22468 17876
rect 22336 17836 22468 17864
rect 22336 17824 22342 17836
rect 22462 17824 22468 17836
rect 22520 17824 22526 17876
rect 26234 17864 26240 17876
rect 26195 17836 26240 17864
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 16574 17756 16580 17808
rect 16632 17796 16638 17808
rect 16914 17799 16972 17805
rect 16914 17796 16926 17799
rect 16632 17768 16926 17796
rect 16632 17756 16638 17768
rect 16914 17765 16926 17768
rect 16960 17765 16972 17799
rect 16914 17759 16972 17765
rect 19426 17756 19432 17808
rect 19484 17796 19490 17808
rect 21729 17799 21787 17805
rect 19484 17768 19748 17796
rect 19484 17756 19490 17768
rect 11784 17731 11842 17737
rect 11784 17697 11796 17731
rect 11830 17728 11842 17731
rect 13446 17728 13452 17740
rect 11830 17700 13452 17728
rect 11830 17697 11842 17700
rect 11784 17691 11842 17697
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 16666 17728 16672 17740
rect 14976 17700 16672 17728
rect 14976 17688 14982 17700
rect 16666 17688 16672 17700
rect 16724 17728 16730 17740
rect 17678 17728 17684 17740
rect 16724 17700 17684 17728
rect 16724 17688 16730 17700
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 18966 17688 18972 17740
rect 19024 17728 19030 17740
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 19024 17700 19533 17728
rect 19024 17688 19030 17700
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 1486 17660 1492 17672
rect 1447 17632 1492 17660
rect 1486 17620 1492 17632
rect 1544 17620 1550 17672
rect 4062 17660 4068 17672
rect 4023 17632 4068 17660
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 15289 17663 15347 17669
rect 10284 17632 10329 17660
rect 10284 17620 10290 17632
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 16482 17660 16488 17672
rect 15335 17632 16488 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 19720 17669 19748 17768
rect 21729 17765 21741 17799
rect 21775 17796 21787 17799
rect 22646 17796 22652 17808
rect 21775 17768 22652 17796
rect 21775 17765 21787 17768
rect 21729 17759 21787 17765
rect 22646 17756 22652 17768
rect 22704 17756 22710 17808
rect 26881 17799 26939 17805
rect 26881 17765 26893 17799
rect 26927 17796 26939 17799
rect 27246 17796 27252 17808
rect 26927 17768 27252 17796
rect 26927 17765 26939 17768
rect 26881 17759 26939 17765
rect 27246 17756 27252 17768
rect 27304 17756 27310 17808
rect 21358 17688 21364 17740
rect 21416 17728 21422 17740
rect 22445 17731 22503 17737
rect 22445 17728 22457 17731
rect 21416 17700 22457 17728
rect 21416 17688 21422 17700
rect 22445 17697 22457 17700
rect 22491 17728 22503 17731
rect 23014 17728 23020 17740
rect 22491 17700 23020 17728
rect 22491 17697 22503 17700
rect 22445 17691 22503 17697
rect 23014 17688 23020 17700
rect 23072 17688 23078 17740
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17728 24823 17731
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 24811 17700 25237 17728
rect 24811 17697 24823 17700
rect 24765 17691 24823 17697
rect 25225 17697 25237 17700
rect 25271 17728 25283 17731
rect 26973 17731 27031 17737
rect 25271 17700 25636 17728
rect 25271 17697 25283 17700
rect 25225 17691 25283 17697
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 20438 17660 20444 17672
rect 19751 17632 20444 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 7929 17595 7987 17601
rect 7929 17561 7941 17595
rect 7975 17592 7987 17595
rect 8680 17592 8708 17620
rect 7975 17564 8708 17592
rect 9677 17595 9735 17601
rect 7975 17561 7987 17564
rect 7929 17555 7987 17561
rect 9677 17561 9689 17595
rect 9723 17592 9735 17595
rect 10870 17592 10876 17604
rect 9723 17564 10876 17592
rect 9723 17561 9735 17564
rect 9677 17555 9735 17561
rect 10870 17552 10876 17564
rect 10928 17552 10934 17604
rect 19628 17592 19656 17623
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 22186 17660 22192 17672
rect 22147 17632 22192 17660
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 25317 17663 25375 17669
rect 25317 17660 25329 17663
rect 24780 17632 25329 17660
rect 24780 17604 24808 17632
rect 25317 17629 25329 17632
rect 25363 17629 25375 17663
rect 25498 17660 25504 17672
rect 25459 17632 25504 17660
rect 25317 17623 25375 17629
rect 25498 17620 25504 17632
rect 25556 17620 25562 17672
rect 25608 17660 25636 17700
rect 26973 17697 26985 17731
rect 27019 17728 27031 17731
rect 27430 17728 27436 17740
rect 27019 17700 27436 17728
rect 27019 17697 27031 17700
rect 26973 17691 27031 17697
rect 27430 17688 27436 17700
rect 27488 17688 27494 17740
rect 27157 17663 27215 17669
rect 25608 17632 27016 17660
rect 19794 17592 19800 17604
rect 19628 17564 19800 17592
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 24762 17552 24768 17604
rect 24820 17552 24826 17604
rect 25961 17595 26019 17601
rect 25961 17561 25973 17595
rect 26007 17592 26019 17595
rect 26878 17592 26884 17604
rect 26007 17564 26884 17592
rect 26007 17561 26019 17564
rect 25961 17555 26019 17561
rect 26878 17552 26884 17564
rect 26936 17552 26942 17604
rect 26988 17592 27016 17632
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 27706 17660 27712 17672
rect 27203 17632 27712 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 27706 17620 27712 17632
rect 27764 17620 27770 17672
rect 27798 17592 27804 17604
rect 26988 17564 27804 17592
rect 27798 17552 27804 17564
rect 27856 17552 27862 17604
rect 8018 17524 8024 17536
rect 7979 17496 8024 17524
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 10686 17524 10692 17536
rect 9364 17496 10692 17524
rect 9364 17484 9370 17496
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 16298 17524 16304 17536
rect 13320 17496 16304 17524
rect 13320 17484 13326 17496
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 18966 17524 18972 17536
rect 18927 17496 18972 17524
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 23566 17524 23572 17536
rect 23527 17496 23572 17524
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 24121 17527 24179 17533
rect 24121 17524 24133 17527
rect 23808 17496 24133 17524
rect 23808 17484 23814 17496
rect 24121 17493 24133 17496
rect 24167 17524 24179 17527
rect 24394 17524 24400 17536
rect 24167 17496 24400 17524
rect 24167 17493 24179 17496
rect 24121 17487 24179 17493
rect 24394 17484 24400 17496
rect 24452 17484 24458 17536
rect 24857 17527 24915 17533
rect 24857 17493 24869 17527
rect 24903 17524 24915 17527
rect 25222 17524 25228 17536
rect 24903 17496 25228 17524
rect 24903 17493 24915 17496
rect 24857 17487 24915 17493
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 26510 17524 26516 17536
rect 26471 17496 26516 17524
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 2958 17320 2964 17332
rect 2919 17292 2964 17320
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 5445 17323 5503 17329
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5626 17320 5632 17332
rect 5491 17292 5632 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 7561 17323 7619 17329
rect 7561 17320 7573 17323
rect 7524 17292 7573 17320
rect 7524 17280 7530 17292
rect 7561 17289 7573 17292
rect 7607 17320 7619 17323
rect 8386 17320 8392 17332
rect 7607 17292 8392 17320
rect 7607 17289 7619 17292
rect 7561 17283 7619 17289
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 9364 17292 9413 17320
rect 9364 17280 9370 17292
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 9732 17292 10517 17320
rect 9732 17280 9738 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 10505 17283 10563 17289
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 12032 17292 12173 17320
rect 12032 17280 12038 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 12161 17283 12219 17289
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12526 17320 12532 17332
rect 12483 17292 12532 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16632 17292 17141 17320
rect 16632 17280 16638 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 21358 17320 21364 17332
rect 21319 17292 21364 17320
rect 17129 17283 17187 17289
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 21818 17320 21824 17332
rect 21779 17292 21824 17320
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 22833 17323 22891 17329
rect 22833 17320 22845 17323
rect 22244 17292 22845 17320
rect 22244 17280 22250 17292
rect 22833 17289 22845 17292
rect 22879 17320 22891 17323
rect 23382 17320 23388 17332
rect 22879 17292 23388 17320
rect 22879 17289 22891 17292
rect 22833 17283 22891 17289
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 25774 17280 25780 17332
rect 25832 17320 25838 17332
rect 25869 17323 25927 17329
rect 25869 17320 25881 17323
rect 25832 17292 25881 17320
rect 25832 17280 25838 17292
rect 25869 17289 25881 17292
rect 25915 17289 25927 17323
rect 26418 17320 26424 17332
rect 26379 17292 26424 17320
rect 25869 17283 25927 17289
rect 10045 17255 10103 17261
rect 10045 17221 10057 17255
rect 10091 17252 10103 17255
rect 10318 17252 10324 17264
rect 10091 17224 10324 17252
rect 10091 17221 10103 17224
rect 10045 17215 10103 17221
rect 10318 17212 10324 17224
rect 10376 17212 10382 17264
rect 16666 17212 16672 17264
rect 16724 17252 16730 17264
rect 16761 17255 16819 17261
rect 16761 17252 16773 17255
rect 16724 17224 16773 17252
rect 16724 17212 16730 17224
rect 16761 17221 16773 17224
rect 16807 17221 16819 17255
rect 16761 17215 16819 17221
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7055 17156 8156 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 1486 17076 1492 17128
rect 1544 17116 1550 17128
rect 4338 17125 4344 17128
rect 1581 17119 1639 17125
rect 1581 17116 1593 17119
rect 1544 17088 1593 17116
rect 1544 17076 1550 17088
rect 1581 17085 1593 17088
rect 1627 17116 1639 17119
rect 4065 17119 4123 17125
rect 1627 17088 3188 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 3160 17060 3188 17088
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4332 17116 4344 17125
rect 4111 17088 4145 17116
rect 4299 17088 4344 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4332 17079 4344 17088
rect 1848 17051 1906 17057
rect 1848 17017 1860 17051
rect 1894 17048 1906 17051
rect 2222 17048 2228 17060
rect 1894 17020 2228 17048
rect 1894 17017 1906 17020
rect 1848 17011 1906 17017
rect 2222 17008 2228 17020
rect 2280 17008 2286 17060
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 3605 17051 3663 17057
rect 3605 17048 3617 17051
rect 3200 17020 3617 17048
rect 3200 17008 3206 17020
rect 3605 17017 3617 17020
rect 3651 17048 3663 17051
rect 3973 17051 4031 17057
rect 3973 17048 3985 17051
rect 3651 17020 3985 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 3973 17017 3985 17020
rect 4019 17048 4031 17051
rect 4080 17048 4108 17079
rect 4338 17076 4344 17079
rect 4396 17076 4402 17128
rect 7926 17116 7932 17128
rect 7887 17088 7932 17116
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17085 8079 17119
rect 8128 17116 8156 17156
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 10744 17156 11069 17184
rect 10744 17144 10750 17156
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13446 17184 13452 17196
rect 13127 17156 13452 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 21729 17187 21787 17193
rect 21729 17153 21741 17187
rect 21775 17184 21787 17187
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 21775 17156 22385 17184
rect 21775 17153 21787 17156
rect 21729 17147 21787 17153
rect 22373 17153 22385 17156
rect 22419 17184 22431 17187
rect 23385 17187 23443 17193
rect 23385 17184 23397 17187
rect 22419 17156 23397 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 23385 17153 23397 17156
rect 23431 17184 23443 17187
rect 23566 17184 23572 17196
rect 23431 17156 23572 17184
rect 23431 17153 23443 17156
rect 23385 17147 23443 17153
rect 23566 17144 23572 17156
rect 23624 17184 23630 17196
rect 23624 17156 24072 17184
rect 23624 17144 23630 17156
rect 10042 17116 10048 17128
rect 8128 17088 10048 17116
rect 8021 17079 8079 17085
rect 5166 17048 5172 17060
rect 4019 17020 5172 17048
rect 4019 17017 4031 17020
rect 3973 17011 4031 17017
rect 5166 17008 5172 17020
rect 5224 17048 5230 17060
rect 6089 17051 6147 17057
rect 6089 17048 6101 17051
rect 5224 17020 6101 17048
rect 5224 17008 5230 17020
rect 6089 17017 6101 17020
rect 6135 17048 6147 17051
rect 8036 17048 8064 17079
rect 10042 17076 10048 17088
rect 10100 17116 10106 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 10100 17088 10333 17116
rect 10100 17076 10106 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10870 17116 10876 17128
rect 10831 17088 10876 17116
rect 10321 17079 10379 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 14645 17119 14703 17125
rect 14645 17116 14657 17119
rect 12860 17088 14657 17116
rect 12860 17076 12866 17088
rect 14645 17085 14657 17088
rect 14691 17116 14703 17119
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14691 17088 14841 17116
rect 14691 17085 14703 17088
rect 14645 17079 14703 17085
rect 14829 17085 14841 17088
rect 14875 17116 14887 17119
rect 14918 17116 14924 17128
rect 14875 17088 14924 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 18417 17119 18475 17125
rect 18417 17116 18429 17119
rect 17736 17088 18429 17116
rect 17736 17076 17742 17088
rect 18417 17085 18429 17088
rect 18463 17116 18475 17119
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 18463 17088 18613 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 21818 17116 21824 17128
rect 20671 17088 21824 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 21818 17076 21824 17088
rect 21876 17116 21882 17128
rect 22189 17119 22247 17125
rect 22189 17116 22201 17119
rect 21876 17088 22201 17116
rect 21876 17076 21882 17088
rect 22189 17085 22201 17088
rect 22235 17085 22247 17119
rect 22189 17079 22247 17085
rect 23937 17119 23995 17125
rect 23937 17085 23949 17119
rect 23983 17085 23995 17119
rect 24044 17116 24072 17156
rect 24193 17119 24251 17125
rect 24193 17116 24205 17119
rect 24044 17088 24205 17116
rect 23937 17079 23995 17085
rect 24193 17085 24205 17088
rect 24239 17085 24251 17119
rect 25884 17116 25912 17283
rect 26418 17280 26424 17292
rect 26476 17280 26482 17332
rect 26326 17212 26332 17264
rect 26384 17252 26390 17264
rect 26384 17224 27016 17252
rect 26384 17212 26390 17224
rect 26878 17184 26884 17196
rect 26839 17156 26884 17184
rect 26878 17144 26884 17156
rect 26936 17144 26942 17196
rect 26988 17193 27016 17224
rect 26973 17187 27031 17193
rect 26973 17153 26985 17187
rect 27019 17184 27031 17187
rect 27522 17184 27528 17196
rect 27019 17156 27528 17184
rect 27019 17153 27031 17156
rect 26973 17147 27031 17153
rect 27522 17144 27528 17156
rect 27580 17184 27586 17196
rect 27801 17187 27859 17193
rect 27801 17184 27813 17187
rect 27580 17156 27813 17184
rect 27580 17144 27586 17156
rect 27801 17153 27813 17156
rect 27847 17153 27859 17187
rect 27801 17147 27859 17153
rect 26786 17116 26792 17128
rect 25884 17088 26792 17116
rect 24193 17079 24251 17085
rect 8110 17048 8116 17060
rect 6135 17020 8116 17048
rect 6135 17017 6147 17020
rect 6089 17011 6147 17017
rect 8110 17008 8116 17020
rect 8168 17008 8174 17060
rect 8288 17051 8346 17057
rect 8288 17017 8300 17051
rect 8334 17048 8346 17051
rect 8662 17048 8668 17060
rect 8334 17020 8668 17048
rect 8334 17017 8346 17020
rect 8288 17011 8346 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 10410 17008 10416 17060
rect 10468 17048 10474 17060
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 10468 17020 10977 17048
rect 10468 17008 10474 17020
rect 10965 17017 10977 17020
rect 11011 17017 11023 17051
rect 10965 17011 11023 17017
rect 12618 17008 12624 17060
rect 12676 17048 12682 17060
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 12676 17020 12909 17048
rect 12676 17008 12682 17020
rect 12897 17017 12909 17020
rect 12943 17017 12955 17051
rect 12897 17011 12955 17017
rect 15010 17008 15016 17060
rect 15068 17057 15074 17060
rect 15068 17051 15132 17057
rect 15068 17017 15086 17051
rect 15120 17017 15132 17051
rect 15068 17011 15132 17017
rect 15068 17008 15074 17011
rect 18506 17008 18512 17060
rect 18564 17048 18570 17060
rect 18846 17051 18904 17057
rect 18846 17048 18858 17051
rect 18564 17020 18858 17048
rect 18564 17008 18570 17020
rect 18846 17017 18858 17020
rect 18892 17017 18904 17051
rect 18846 17011 18904 17017
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17048 21051 17051
rect 21634 17048 21640 17060
rect 21039 17020 21640 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 21634 17008 21640 17020
rect 21692 17048 21698 17060
rect 22281 17051 22339 17057
rect 22281 17048 22293 17051
rect 21692 17020 22293 17048
rect 21692 17008 21698 17020
rect 22281 17017 22293 17020
rect 22327 17017 22339 17051
rect 22281 17011 22339 17017
rect 23382 17008 23388 17060
rect 23440 17048 23446 17060
rect 23952 17048 23980 17079
rect 26786 17076 26792 17088
rect 26844 17076 26850 17128
rect 24026 17048 24032 17060
rect 23440 17020 24032 17048
rect 23440 17008 23446 17020
rect 24026 17008 24032 17020
rect 24084 17008 24090 17060
rect 25498 17048 25504 17060
rect 25332 17020 25504 17048
rect 6549 16983 6607 16989
rect 6549 16949 6561 16983
rect 6595 16980 6607 16983
rect 6914 16980 6920 16992
rect 6595 16952 6920 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 6914 16940 6920 16952
rect 6972 16940 6978 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12032 16952 12817 16980
rect 12032 16940 12038 16952
rect 12805 16949 12817 16952
rect 12851 16980 12863 16983
rect 13170 16980 13176 16992
rect 12851 16952 13176 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 13446 16980 13452 16992
rect 13407 16952 13452 16980
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 15746 16940 15752 16992
rect 15804 16980 15810 16992
rect 16209 16983 16267 16989
rect 16209 16980 16221 16983
rect 15804 16952 16221 16980
rect 15804 16940 15810 16952
rect 16209 16949 16221 16952
rect 16255 16949 16267 16983
rect 16209 16943 16267 16949
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 19944 16952 19993 16980
rect 19944 16940 19950 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 21542 16940 21548 16992
rect 21600 16980 21606 16992
rect 22186 16980 22192 16992
rect 21600 16952 22192 16980
rect 21600 16940 21606 16952
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 25332 16989 25360 17020
rect 25498 17008 25504 17020
rect 25556 17048 25562 17060
rect 26418 17048 26424 17060
rect 25556 17020 26424 17048
rect 25556 17008 25562 17020
rect 26418 17008 26424 17020
rect 26476 17008 26482 17060
rect 25317 16983 25375 16989
rect 25317 16949 25329 16983
rect 25363 16949 25375 16983
rect 26326 16980 26332 16992
rect 26239 16952 26332 16980
rect 25317 16943 25375 16949
rect 26326 16940 26332 16952
rect 26384 16980 26390 16992
rect 27246 16980 27252 16992
rect 26384 16952 27252 16980
rect 26384 16940 26390 16952
rect 27246 16940 27252 16952
rect 27304 16940 27310 16992
rect 27430 16980 27436 16992
rect 27391 16952 27436 16980
rect 27430 16940 27436 16952
rect 27488 16940 27494 16992
rect 27706 16940 27712 16992
rect 27764 16980 27770 16992
rect 28169 16983 28227 16989
rect 28169 16980 28181 16983
rect 27764 16952 28181 16980
rect 27764 16940 27770 16952
rect 28169 16949 28181 16952
rect 28215 16949 28227 16983
rect 28169 16943 28227 16949
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 2041 16779 2099 16785
rect 2041 16745 2053 16779
rect 2087 16776 2099 16779
rect 2682 16776 2688 16788
rect 2087 16748 2688 16776
rect 2087 16745 2099 16748
rect 2041 16739 2099 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 3142 16776 3148 16788
rect 3103 16748 3148 16776
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16776 3574 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3568 16748 3801 16776
rect 3568 16736 3574 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 3804 16708 3832 16739
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4120 16748 4445 16776
rect 4120 16736 4126 16748
rect 4433 16745 4445 16748
rect 4479 16776 4491 16779
rect 4522 16776 4528 16788
rect 4479 16748 4528 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 5626 16776 5632 16788
rect 5587 16748 5632 16776
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 6730 16776 6736 16788
rect 6503 16748 6736 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 6914 16736 6920 16748
rect 6972 16776 6978 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 6972 16748 8033 16776
rect 6972 16736 6978 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 9953 16779 10011 16785
rect 9953 16745 9965 16779
rect 9999 16776 10011 16779
rect 10226 16776 10232 16788
rect 9999 16748 10232 16776
rect 9999 16745 10011 16748
rect 9953 16739 10011 16745
rect 4614 16708 4620 16720
rect 3804 16680 4620 16708
rect 4614 16668 4620 16680
rect 4672 16708 4678 16720
rect 5902 16708 5908 16720
rect 4672 16680 4752 16708
rect 5863 16680 5908 16708
rect 4672 16668 4678 16680
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2590 16640 2596 16652
rect 2179 16612 2596 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2590 16600 2596 16612
rect 2648 16640 2654 16652
rect 2685 16643 2743 16649
rect 2685 16640 2697 16643
rect 2648 16612 2697 16640
rect 2648 16600 2654 16612
rect 2685 16609 2697 16612
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 3016 16612 4108 16640
rect 3016 16600 3022 16612
rect 2222 16572 2228 16584
rect 2135 16544 2228 16572
rect 2222 16532 2228 16544
rect 2280 16572 2286 16584
rect 3510 16572 3516 16584
rect 2280 16544 3516 16572
rect 2280 16532 2286 16544
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 4080 16513 4108 16612
rect 4430 16532 4436 16584
rect 4488 16572 4494 16584
rect 4724 16581 4752 16680
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 8570 16640 8576 16652
rect 8435 16612 8576 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 4525 16575 4583 16581
rect 4525 16572 4537 16575
rect 4488 16544 4537 16572
rect 4488 16532 4494 16544
rect 4525 16541 4537 16544
rect 4571 16541 4583 16575
rect 4525 16535 4583 16541
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16541 4767 16575
rect 4709 16535 4767 16541
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7282 16572 7288 16584
rect 7147 16544 7288 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 4065 16507 4123 16513
rect 4065 16473 4077 16507
rect 4111 16473 4123 16507
rect 4065 16467 4123 16473
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 7116 16504 7144 16535
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 8478 16572 8484 16584
rect 8439 16544 8484 16572
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 9968 16572 9996 16739
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 10410 16776 10416 16788
rect 10371 16748 10416 16776
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 12802 16776 12808 16788
rect 11572 16748 12808 16776
rect 11572 16736 11578 16748
rect 12802 16736 12808 16748
rect 12860 16776 12866 16788
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12860 16748 12909 16776
rect 12860 16736 12866 16748
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 12897 16739 12955 16745
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13814 16776 13820 16788
rect 13127 16748 13820 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 17310 16776 17316 16788
rect 17271 16748 17316 16776
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 18966 16776 18972 16788
rect 18647 16748 18972 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 19484 16748 19625 16776
rect 19484 16736 19490 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 19981 16779 20039 16785
rect 19981 16776 19993 16779
rect 19852 16748 19993 16776
rect 19852 16736 19858 16748
rect 19981 16745 19993 16748
rect 20027 16745 20039 16779
rect 19981 16739 20039 16745
rect 21545 16779 21603 16785
rect 21545 16745 21557 16779
rect 21591 16776 21603 16779
rect 22002 16776 22008 16788
rect 21591 16748 22008 16776
rect 21591 16745 21603 16748
rect 21545 16739 21603 16745
rect 22002 16736 22008 16748
rect 22060 16736 22066 16788
rect 23014 16776 23020 16788
rect 22975 16748 23020 16776
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 24026 16776 24032 16788
rect 23987 16748 24032 16776
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 24397 16779 24455 16785
rect 24397 16745 24409 16779
rect 24443 16776 24455 16779
rect 25498 16776 25504 16788
rect 24443 16748 25504 16776
rect 24443 16745 24455 16748
rect 24397 16739 24455 16745
rect 25498 16736 25504 16748
rect 25556 16736 25562 16788
rect 26513 16779 26571 16785
rect 26513 16745 26525 16779
rect 26559 16776 26571 16779
rect 26878 16776 26884 16788
rect 26559 16748 26884 16776
rect 26559 16745 26571 16748
rect 26513 16739 26571 16745
rect 26878 16736 26884 16748
rect 26936 16736 26942 16788
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 10864 16711 10922 16717
rect 10864 16708 10876 16711
rect 10192 16680 10876 16708
rect 10192 16668 10198 16680
rect 10864 16677 10876 16680
rect 10910 16708 10922 16711
rect 10962 16708 10968 16720
rect 10910 16680 10968 16708
rect 10910 16677 10922 16680
rect 10864 16671 10922 16677
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 13262 16708 13268 16720
rect 12216 16680 13268 16708
rect 12216 16668 12222 16680
rect 13262 16668 13268 16680
rect 13320 16708 13326 16720
rect 13449 16711 13507 16717
rect 13449 16708 13461 16711
rect 13320 16680 13461 16708
rect 13320 16668 13326 16680
rect 13449 16677 13461 16680
rect 13495 16677 13507 16711
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 13449 16671 13507 16677
rect 15212 16680 15761 16708
rect 12618 16640 12624 16652
rect 12579 16612 12624 16640
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13630 16640 13636 16652
rect 13587 16612 13636 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 15212 16640 15240 16680
rect 15749 16677 15761 16680
rect 15795 16677 15807 16711
rect 15749 16671 15807 16677
rect 16482 16668 16488 16720
rect 16540 16708 16546 16720
rect 17218 16708 17224 16720
rect 16540 16680 17224 16708
rect 16540 16668 16546 16680
rect 17218 16668 17224 16680
rect 17276 16668 17282 16720
rect 18414 16668 18420 16720
rect 18472 16708 18478 16720
rect 19812 16708 19840 16736
rect 18472 16680 19840 16708
rect 21177 16711 21235 16717
rect 18472 16668 18478 16680
rect 21177 16677 21189 16711
rect 21223 16708 21235 16711
rect 21726 16708 21732 16720
rect 21223 16680 21732 16708
rect 21223 16677 21235 16680
rect 21177 16671 21235 16677
rect 21726 16668 21732 16680
rect 21784 16708 21790 16720
rect 22094 16708 22100 16720
rect 21784 16680 22100 16708
rect 21784 16668 21790 16680
rect 22094 16668 22100 16680
rect 22152 16668 22158 16720
rect 23661 16711 23719 16717
rect 23661 16677 23673 16711
rect 23707 16708 23719 16711
rect 24854 16708 24860 16720
rect 23707 16680 24860 16708
rect 23707 16677 23719 16680
rect 23661 16671 23719 16677
rect 24854 16668 24860 16680
rect 24912 16708 24918 16720
rect 25317 16711 25375 16717
rect 25317 16708 25329 16711
rect 24912 16680 25329 16708
rect 24912 16668 24918 16680
rect 25317 16677 25329 16680
rect 25363 16677 25375 16711
rect 25317 16671 25375 16677
rect 25866 16668 25872 16720
rect 25924 16708 25930 16720
rect 26973 16711 27031 16717
rect 26973 16708 26985 16711
rect 25924 16680 26985 16708
rect 25924 16668 25930 16680
rect 26973 16677 26985 16680
rect 27019 16677 27031 16711
rect 26973 16671 27031 16677
rect 15378 16640 15384 16652
rect 15120 16612 15240 16640
rect 15304 16612 15384 16640
rect 10594 16572 10600 16584
rect 8720 16544 9996 16572
rect 10555 16544 10600 16572
rect 8720 16532 8726 16544
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 13722 16572 13728 16584
rect 13683 16544 13728 16572
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 15120 16572 15148 16612
rect 13872 16544 15148 16572
rect 13872 16532 13878 16544
rect 7558 16504 7564 16516
rect 6411 16476 7144 16504
rect 7471 16476 7564 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 7558 16464 7564 16476
rect 7616 16504 7622 16516
rect 8680 16504 8708 16532
rect 15304 16513 15332 16612
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 16850 16600 16856 16652
rect 16908 16600 16914 16652
rect 18230 16600 18236 16652
rect 18288 16640 18294 16652
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18288 16612 18981 16640
rect 18288 16600 18294 16612
rect 18969 16609 18981 16612
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19116 16612 19161 16640
rect 19116 16600 19122 16612
rect 21266 16600 21272 16652
rect 21324 16640 21330 16652
rect 21904 16643 21962 16649
rect 21904 16640 21916 16643
rect 21324 16612 21916 16640
rect 21324 16600 21330 16612
rect 21904 16609 21916 16612
rect 21950 16640 21962 16643
rect 22646 16640 22652 16652
rect 21950 16612 22652 16640
rect 21950 16609 21962 16612
rect 21904 16603 21962 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 24762 16640 24768 16652
rect 24723 16612 24768 16640
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 24946 16640 24952 16652
rect 24872 16612 24952 16640
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 16868 16513 16896 16600
rect 17402 16572 17408 16584
rect 17363 16544 17408 16572
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 18417 16575 18475 16581
rect 18417 16572 18429 16575
rect 17736 16544 18429 16572
rect 17736 16532 17742 16544
rect 18417 16541 18429 16544
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 19153 16575 19211 16581
rect 19153 16541 19165 16575
rect 19199 16572 19211 16575
rect 19886 16572 19892 16584
rect 19199 16544 19892 16572
rect 19199 16541 19211 16544
rect 19153 16535 19211 16541
rect 7616 16476 8708 16504
rect 15289 16507 15347 16513
rect 7616 16464 7622 16476
rect 15289 16473 15301 16507
rect 15335 16473 15347 16507
rect 15289 16467 15347 16473
rect 16853 16507 16911 16513
rect 16853 16473 16865 16507
rect 16899 16473 16911 16507
rect 16853 16467 16911 16473
rect 18966 16464 18972 16516
rect 19024 16504 19030 16516
rect 19168 16504 19196 16535
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 21542 16532 21548 16584
rect 21600 16572 21606 16584
rect 21637 16575 21695 16581
rect 21637 16572 21649 16575
rect 21600 16544 21649 16572
rect 21600 16532 21606 16544
rect 21637 16541 21649 16544
rect 21683 16541 21695 16575
rect 21637 16535 21695 16541
rect 19024 16476 19196 16504
rect 19024 16464 19030 16476
rect 5261 16439 5319 16445
rect 5261 16405 5273 16439
rect 5307 16436 5319 16439
rect 5626 16436 5632 16448
rect 5307 16408 5632 16436
rect 5307 16405 5319 16408
rect 5261 16399 5319 16405
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8110 16436 8116 16448
rect 7975 16408 8116 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8110 16396 8116 16408
rect 8168 16436 8174 16448
rect 8386 16436 8392 16448
rect 8168 16408 8392 16436
rect 8168 16396 8174 16408
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 9030 16436 9036 16448
rect 8991 16408 9036 16436
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 11977 16439 12035 16445
rect 11977 16405 11989 16439
rect 12023 16436 12035 16439
rect 12342 16436 12348 16448
rect 12023 16408 12348 16436
rect 12023 16405 12035 16408
rect 11977 16399 12035 16405
rect 12342 16396 12348 16408
rect 12400 16396 12406 16448
rect 15010 16436 15016 16448
rect 14971 16408 15016 16436
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 21652 16436 21680 16535
rect 24872 16513 24900 16612
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 25222 16640 25228 16652
rect 25183 16612 25228 16640
rect 25222 16600 25228 16612
rect 25280 16600 25286 16652
rect 26878 16640 26884 16652
rect 26160 16612 26884 16640
rect 25314 16532 25320 16584
rect 25372 16572 25378 16584
rect 25409 16575 25467 16581
rect 25409 16572 25421 16575
rect 25372 16544 25421 16572
rect 25372 16532 25378 16544
rect 25409 16541 25421 16544
rect 25455 16541 25467 16575
rect 25409 16535 25467 16541
rect 25590 16532 25596 16584
rect 25648 16572 25654 16584
rect 26160 16572 26188 16612
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 25648 16544 26188 16572
rect 26237 16575 26295 16581
rect 25648 16532 25654 16544
rect 26237 16541 26249 16575
rect 26283 16572 26295 16575
rect 26418 16572 26424 16584
rect 26283 16544 26424 16572
rect 26283 16541 26295 16544
rect 26237 16535 26295 16541
rect 26418 16532 26424 16544
rect 26476 16572 26482 16584
rect 27154 16572 27160 16584
rect 26476 16544 27160 16572
rect 26476 16532 26482 16544
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 24857 16507 24915 16513
rect 24857 16473 24869 16507
rect 24903 16473 24915 16507
rect 24857 16467 24915 16473
rect 21910 16436 21916 16448
rect 21652 16408 21916 16436
rect 21910 16396 21916 16408
rect 21968 16396 21974 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2682 16232 2688 16244
rect 2643 16204 2688 16232
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 3050 16232 3056 16244
rect 3011 16204 3056 16232
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 3145 16235 3203 16241
rect 3145 16201 3157 16235
rect 3191 16232 3203 16235
rect 3418 16232 3424 16244
rect 3191 16204 3424 16232
rect 3191 16201 3203 16204
rect 3145 16195 3203 16201
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 4522 16232 4528 16244
rect 4483 16204 4528 16232
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6454 16232 6460 16244
rect 6319 16204 6460 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 4430 16164 4436 16176
rect 4295 16136 4436 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 4430 16124 4436 16136
rect 4488 16124 4494 16176
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 3510 16056 3516 16108
rect 3568 16096 3574 16108
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 3568 16068 3709 16096
rect 3568 16056 3574 16068
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 5810 16096 5816 16108
rect 5723 16068 5816 16096
rect 3697 16059 3755 16065
rect 5810 16056 5816 16068
rect 5868 16096 5874 16108
rect 6288 16096 6316 16195
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 6546 16192 6552 16244
rect 6604 16232 6610 16244
rect 9861 16235 9919 16241
rect 6604 16204 6649 16232
rect 6604 16192 6610 16204
rect 9861 16201 9873 16235
rect 9907 16232 9919 16235
rect 10226 16232 10232 16244
rect 9907 16204 10232 16232
rect 9907 16201 9919 16204
rect 9861 16195 9919 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 11054 16232 11060 16244
rect 11015 16204 11060 16232
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 14185 16235 14243 16241
rect 14185 16201 14197 16235
rect 14231 16232 14243 16235
rect 15010 16232 15016 16244
rect 14231 16204 15016 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 15010 16192 15016 16204
rect 15068 16232 15074 16244
rect 15562 16232 15568 16244
rect 15068 16204 15568 16232
rect 15068 16192 15074 16204
rect 15562 16192 15568 16204
rect 15620 16232 15626 16244
rect 16393 16235 16451 16241
rect 15620 16204 15884 16232
rect 15620 16192 15626 16204
rect 14734 16164 14740 16176
rect 14695 16136 14740 16164
rect 14734 16124 14740 16136
rect 14792 16164 14798 16176
rect 14792 16136 15792 16164
rect 14792 16124 14798 16136
rect 7558 16096 7564 16108
rect 5868 16068 6316 16096
rect 7519 16068 7564 16096
rect 5868 16056 5874 16068
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 12802 16096 12808 16108
rect 12763 16068 12808 16096
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 15764 16105 15792 16136
rect 15856 16105 15884 16204
rect 16393 16201 16405 16235
rect 16439 16232 16451 16235
rect 16482 16232 16488 16244
rect 16439 16204 16488 16232
rect 16439 16201 16451 16204
rect 16393 16195 16451 16201
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15841 16099 15899 16105
rect 15841 16065 15853 16099
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 6604 16000 7297 16028
rect 6604 15988 6610 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 13078 16037 13084 16040
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 8444 16000 8493 16028
rect 8444 15988 8450 16000
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 11885 16031 11943 16037
rect 11885 15997 11897 16031
rect 11931 16028 11943 16031
rect 13072 16028 13084 16037
rect 11931 16000 13084 16028
rect 11931 15997 11943 16000
rect 11885 15991 11943 15997
rect 13072 15991 13084 16000
rect 13078 15988 13084 15991
rect 13136 15988 13142 16040
rect 15470 15988 15476 16040
rect 15528 16028 15534 16040
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15528 16000 15669 16028
rect 15528 15988 15534 16000
rect 15657 15997 15669 16000
rect 15703 16028 15715 16031
rect 16408 16028 16436 16195
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 18230 16232 18236 16244
rect 18191 16204 18236 16232
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 21266 16232 21272 16244
rect 21227 16204 21272 16232
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 21818 16232 21824 16244
rect 21779 16204 21824 16232
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 24026 16232 24032 16244
rect 23523 16204 24032 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 16945 16167 17003 16173
rect 16945 16133 16957 16167
rect 16991 16164 17003 16167
rect 17310 16164 17316 16176
rect 16991 16136 17316 16164
rect 16991 16133 17003 16136
rect 16945 16127 17003 16133
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18230 16096 18236 16108
rect 17736 16068 18236 16096
rect 17736 16056 17742 16068
rect 18230 16056 18236 16068
rect 18288 16096 18294 16108
rect 18417 16099 18475 16105
rect 18417 16096 18429 16099
rect 18288 16068 18429 16096
rect 18288 16056 18294 16068
rect 18417 16065 18429 16068
rect 18463 16065 18475 16099
rect 18417 16059 18475 16065
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21358 16096 21364 16108
rect 21039 16068 21364 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 23676 16105 23704 16204
rect 24026 16192 24032 16204
rect 24084 16232 24090 16244
rect 24084 16204 24624 16232
rect 24084 16192 24090 16204
rect 24596 16164 24624 16204
rect 24670 16192 24676 16244
rect 24728 16232 24734 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24728 16204 25053 16232
rect 24728 16192 24734 16204
rect 25041 16201 25053 16204
rect 25087 16232 25099 16235
rect 25774 16232 25780 16244
rect 25087 16204 25780 16232
rect 25087 16201 25099 16204
rect 25041 16195 25099 16201
rect 25774 16192 25780 16204
rect 25832 16192 25838 16244
rect 27154 16192 27160 16244
rect 27212 16232 27218 16244
rect 28077 16235 28135 16241
rect 28077 16232 28089 16235
rect 27212 16204 28089 16232
rect 27212 16192 27218 16204
rect 28077 16201 28089 16204
rect 28123 16201 28135 16235
rect 28077 16195 28135 16201
rect 27522 16164 27528 16176
rect 24596 16136 26188 16164
rect 27483 16136 27528 16164
rect 26160 16108 26188 16136
rect 27522 16124 27528 16136
rect 27580 16124 27586 16176
rect 22465 16099 22523 16105
rect 22465 16065 22477 16099
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16065 23719 16099
rect 26142 16096 26148 16108
rect 26055 16068 26148 16096
rect 23661 16059 23719 16065
rect 15703 16000 16436 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 22189 16031 22247 16037
rect 22189 16028 22201 16031
rect 22152 16000 22201 16028
rect 22152 15988 22158 16000
rect 22189 15997 22201 16000
rect 22235 15997 22247 16031
rect 22189 15991 22247 15997
rect 22370 15988 22376 16040
rect 22428 16028 22434 16040
rect 22480 16028 22508 16059
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 26418 16037 26424 16040
rect 26412 16028 26424 16037
rect 22428 16000 22508 16028
rect 26379 16000 26424 16028
rect 22428 15988 22434 16000
rect 26412 15991 26424 16000
rect 26418 15988 26424 15991
rect 26476 15988 26482 16040
rect 1946 15960 1952 15972
rect 1907 15932 1952 15960
rect 1946 15920 1952 15932
rect 2004 15920 2010 15972
rect 3050 15920 3056 15972
rect 3108 15960 3114 15972
rect 3418 15960 3424 15972
rect 3108 15932 3424 15960
rect 3108 15920 3114 15932
rect 3418 15920 3424 15932
rect 3476 15960 3482 15972
rect 3513 15963 3571 15969
rect 3513 15960 3525 15963
rect 3476 15932 3525 15960
rect 3476 15920 3482 15932
rect 3513 15929 3525 15932
rect 3559 15929 3571 15963
rect 3513 15923 3571 15929
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 5077 15963 5135 15969
rect 5077 15960 5089 15963
rect 5040 15932 5089 15960
rect 5040 15920 5046 15932
rect 5077 15929 5089 15932
rect 5123 15960 5135 15963
rect 5123 15932 5580 15960
rect 5123 15929 5135 15932
rect 5077 15923 5135 15929
rect 5552 15904 5580 15932
rect 8294 15920 8300 15972
rect 8352 15960 8358 15972
rect 8726 15963 8784 15969
rect 8726 15960 8738 15963
rect 8352 15932 8738 15960
rect 8352 15920 8358 15932
rect 8726 15929 8738 15932
rect 8772 15960 8784 15963
rect 9030 15960 9036 15972
rect 8772 15932 9036 15960
rect 8772 15929 8784 15932
rect 8726 15923 8784 15929
rect 9030 15920 9036 15932
rect 9088 15920 9094 15972
rect 11606 15920 11612 15972
rect 11664 15960 11670 15972
rect 12621 15963 12679 15969
rect 12621 15960 12633 15963
rect 11664 15932 12633 15960
rect 11664 15920 11670 15932
rect 12621 15929 12633 15932
rect 12667 15960 12679 15963
rect 13630 15960 13636 15972
rect 12667 15932 13636 15960
rect 12667 15929 12679 15932
rect 12621 15923 12679 15929
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 15197 15963 15255 15969
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 17034 15960 17040 15972
rect 15243 15932 17040 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 15672 15904 15700 15932
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 17865 15963 17923 15969
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18322 15960 18328 15972
rect 17911 15932 18328 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 18322 15920 18328 15932
rect 18380 15960 18386 15972
rect 18662 15963 18720 15969
rect 18662 15960 18674 15963
rect 18380 15932 18674 15960
rect 18380 15920 18386 15932
rect 18662 15929 18674 15932
rect 18708 15929 18720 15963
rect 18662 15923 18720 15929
rect 19058 15920 19064 15972
rect 19116 15960 19122 15972
rect 20349 15963 20407 15969
rect 20349 15960 20361 15963
rect 19116 15932 20361 15960
rect 19116 15920 19122 15932
rect 20349 15929 20361 15932
rect 20395 15929 20407 15963
rect 20349 15923 20407 15929
rect 23109 15963 23167 15969
rect 23109 15929 23121 15963
rect 23155 15960 23167 15963
rect 23906 15963 23964 15969
rect 23906 15960 23918 15963
rect 23155 15932 23918 15960
rect 23155 15929 23167 15932
rect 23109 15923 23167 15929
rect 23906 15929 23918 15932
rect 23952 15960 23964 15963
rect 24486 15960 24492 15972
rect 23952 15932 24492 15960
rect 23952 15929 23964 15932
rect 23906 15923 23964 15929
rect 24486 15920 24492 15932
rect 24544 15920 24550 15972
rect 25406 15920 25412 15972
rect 25464 15960 25470 15972
rect 25866 15960 25872 15972
rect 25464 15932 25872 15960
rect 25464 15920 25470 15932
rect 25866 15920 25872 15932
rect 25924 15960 25930 15972
rect 25961 15963 26019 15969
rect 25961 15960 25973 15963
rect 25924 15932 25973 15960
rect 25924 15920 25930 15932
rect 25961 15929 25973 15932
rect 26007 15929 26019 15963
rect 25961 15923 26019 15929
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 3605 15895 3663 15901
rect 3605 15892 3617 15895
rect 3292 15864 3617 15892
rect 3292 15852 3298 15864
rect 3605 15861 3617 15864
rect 3651 15861 3663 15895
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 3605 15855 3663 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 6914 15892 6920 15904
rect 5684 15864 5729 15892
rect 6875 15864 6920 15892
rect 5684 15852 5690 15864
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 7340 15864 7389 15892
rect 7340 15852 7346 15864
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 7377 15855 7435 15861
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15892 8171 15895
rect 8570 15892 8576 15904
rect 8159 15864 8576 15892
rect 8159 15861 8171 15864
rect 8113 15855 8171 15861
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 10134 15852 10140 15904
rect 10192 15892 10198 15904
rect 10594 15892 10600 15904
rect 10192 15864 10600 15892
rect 10192 15852 10198 15864
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11330 15892 11336 15904
rect 11291 15864 11336 15892
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 15286 15892 15292 15904
rect 15247 15864 15292 15892
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15654 15852 15660 15904
rect 15712 15852 15718 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19797 15895 19855 15901
rect 19797 15892 19809 15895
rect 19392 15864 19809 15892
rect 19392 15852 19398 15864
rect 19797 15861 19809 15864
rect 19843 15861 19855 15895
rect 19797 15855 19855 15861
rect 21729 15895 21787 15901
rect 21729 15861 21741 15895
rect 21775 15892 21787 15895
rect 21910 15892 21916 15904
rect 21775 15864 21916 15892
rect 21775 15861 21787 15864
rect 21729 15855 21787 15861
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 22281 15895 22339 15901
rect 22281 15892 22293 15895
rect 22244 15864 22293 15892
rect 22244 15852 22250 15864
rect 22281 15861 22293 15864
rect 22327 15861 22339 15895
rect 25590 15892 25596 15904
rect 25551 15864 25596 15892
rect 22281 15855 22339 15861
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 1946 15688 1952 15700
rect 1719 15660 1952 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 4614 15688 4620 15700
rect 4575 15660 4620 15688
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 5408 15660 6285 15688
rect 5408 15648 5414 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7558 15688 7564 15700
rect 7423 15660 7564 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7558 15648 7564 15660
rect 7616 15688 7622 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7616 15660 7849 15688
rect 7616 15648 7622 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8478 15688 8484 15700
rect 8067 15660 8484 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8478 15648 8484 15660
rect 8536 15688 8542 15700
rect 9401 15691 9459 15697
rect 9401 15688 9413 15691
rect 8536 15660 9413 15688
rect 8536 15648 8542 15660
rect 9401 15657 9413 15660
rect 9447 15657 9459 15691
rect 9401 15651 9459 15657
rect 10597 15691 10655 15697
rect 10597 15657 10609 15691
rect 10643 15688 10655 15691
rect 10778 15688 10784 15700
rect 10643 15660 10784 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 12342 15648 12348 15700
rect 12400 15688 12406 15700
rect 13722 15688 13728 15700
rect 12400 15660 13728 15688
rect 12400 15648 12406 15660
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 13872 15660 14657 15688
rect 13872 15648 13878 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 15105 15691 15163 15697
rect 15105 15657 15117 15691
rect 15151 15688 15163 15691
rect 15838 15688 15844 15700
rect 15151 15660 15844 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 2225 15623 2283 15629
rect 2225 15620 2237 15623
rect 1964 15592 2237 15620
rect 1964 15564 1992 15592
rect 2225 15589 2237 15592
rect 2271 15589 2283 15623
rect 2225 15583 2283 15589
rect 2590 15580 2596 15632
rect 2648 15620 2654 15632
rect 6917 15623 6975 15629
rect 6917 15620 6929 15623
rect 2648 15592 6929 15620
rect 2648 15580 2654 15592
rect 6917 15589 6929 15592
rect 6963 15620 6975 15623
rect 7282 15620 7288 15632
rect 6963 15592 7288 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 7282 15580 7288 15592
rect 7340 15620 7346 15632
rect 8570 15620 8576 15632
rect 7340 15592 8576 15620
rect 7340 15580 7346 15592
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 10137 15623 10195 15629
rect 10137 15589 10149 15623
rect 10183 15620 10195 15623
rect 10686 15620 10692 15632
rect 10183 15592 10692 15620
rect 10183 15589 10195 15592
rect 10137 15583 10195 15589
rect 10686 15580 10692 15592
rect 10744 15620 10750 15632
rect 10744 15592 10824 15620
rect 10744 15580 10750 15592
rect 1946 15512 1952 15564
rect 2004 15512 2010 15564
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 2179 15524 2789 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 2777 15521 2789 15524
rect 2823 15552 2835 15555
rect 4062 15552 4068 15564
rect 2823 15524 4068 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4893 15555 4951 15561
rect 4893 15552 4905 15555
rect 4387 15524 4905 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4893 15521 4905 15524
rect 4939 15552 4951 15555
rect 4982 15552 4988 15564
rect 4939 15524 4988 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5160 15555 5218 15561
rect 5160 15521 5172 15555
rect 5206 15552 5218 15555
rect 5442 15552 5448 15564
rect 5206 15524 5448 15552
rect 5206 15521 5218 15524
rect 5160 15515 5218 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 7708 15524 8401 15552
rect 7708 15512 7714 15524
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 2866 15484 2872 15496
rect 2372 15456 2872 15484
rect 2372 15444 2378 15456
rect 2866 15444 2872 15456
rect 2924 15484 2930 15496
rect 3513 15487 3571 15493
rect 3513 15484 3525 15487
rect 2924 15456 3525 15484
rect 2924 15444 2930 15456
rect 3513 15453 3525 15456
rect 3559 15453 3571 15487
rect 8478 15484 8484 15496
rect 8439 15456 8484 15484
rect 3513 15447 3571 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15416 1823 15419
rect 2038 15416 2044 15428
rect 1811 15388 2044 15416
rect 1811 15385 1823 15388
rect 1765 15379 1823 15385
rect 2038 15376 2044 15388
rect 2096 15376 2102 15428
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 8588 15416 8616 15447
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10796 15493 10824 15592
rect 12060 15555 12118 15561
rect 12060 15521 12072 15555
rect 12106 15552 12118 15555
rect 12342 15552 12348 15564
rect 12106 15524 12348 15552
rect 12106 15521 12118 15524
rect 12060 15515 12118 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10652 15456 10701 15484
rect 10652 15444 10658 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 10781 15487 10839 15493
rect 10781 15453 10793 15487
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11609 15487 11667 15493
rect 11609 15484 11621 15487
rect 11296 15456 11621 15484
rect 11296 15444 11302 15456
rect 11609 15453 11621 15456
rect 11655 15453 11667 15487
rect 11790 15484 11796 15496
rect 11751 15456 11796 15484
rect 11609 15447 11667 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 9582 15416 9588 15428
rect 8352 15388 9588 15416
rect 8352 15376 8358 15388
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 10229 15419 10287 15425
rect 10229 15416 10241 15419
rect 9692 15388 10241 15416
rect 3234 15348 3240 15360
rect 3195 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 8386 15308 8392 15360
rect 8444 15348 8450 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8444 15320 9045 15348
rect 8444 15308 8450 15320
rect 9033 15317 9045 15320
rect 9079 15317 9091 15351
rect 9033 15311 9091 15317
rect 9490 15308 9496 15360
rect 9548 15348 9554 15360
rect 9692 15348 9720 15388
rect 10229 15385 10241 15388
rect 10275 15385 10287 15419
rect 10229 15379 10287 15385
rect 13173 15419 13231 15425
rect 13173 15385 13185 15419
rect 13219 15416 13231 15419
rect 13446 15416 13452 15428
rect 13219 15388 13452 15416
rect 13219 15385 13231 15388
rect 13173 15379 13231 15385
rect 13446 15376 13452 15388
rect 13504 15416 13510 15428
rect 15120 15416 15148 15651
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16298 15648 16304 15700
rect 16356 15688 16362 15700
rect 16669 15691 16727 15697
rect 16669 15688 16681 15691
rect 16356 15660 16681 15688
rect 16356 15648 16362 15660
rect 16669 15657 16681 15660
rect 16715 15688 16727 15691
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 16715 15660 17233 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 17221 15657 17233 15660
rect 17267 15688 17279 15691
rect 17402 15688 17408 15700
rect 17267 15660 17408 15688
rect 17267 15657 17279 15660
rect 17221 15651 17279 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 18414 15688 18420 15700
rect 18375 15660 18420 15688
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 21358 15648 21364 15700
rect 21416 15688 21422 15700
rect 21821 15691 21879 15697
rect 21821 15688 21833 15691
rect 21416 15660 21833 15688
rect 21416 15648 21422 15660
rect 21821 15657 21833 15660
rect 21867 15688 21879 15691
rect 22370 15688 22376 15700
rect 21867 15660 22376 15688
rect 21867 15657 21879 15660
rect 21821 15651 21879 15657
rect 22370 15648 22376 15660
rect 22428 15648 22434 15700
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 23293 15691 23351 15697
rect 23293 15688 23305 15691
rect 22704 15660 23305 15688
rect 22704 15648 22710 15660
rect 23293 15657 23305 15660
rect 23339 15688 23351 15691
rect 23382 15688 23388 15700
rect 23339 15660 23388 15688
rect 23339 15657 23351 15660
rect 23293 15651 23351 15657
rect 23382 15648 23388 15660
rect 23440 15648 23446 15700
rect 24854 15688 24860 15700
rect 24815 15660 24860 15688
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 26142 15688 26148 15700
rect 26103 15660 26148 15688
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 26510 15648 26516 15700
rect 26568 15688 26574 15700
rect 26881 15691 26939 15697
rect 26881 15688 26893 15691
rect 26568 15660 26893 15688
rect 26568 15648 26574 15660
rect 26881 15657 26893 15660
rect 26927 15688 26939 15691
rect 27614 15688 27620 15700
rect 26927 15660 27620 15688
rect 26927 15657 26939 15660
rect 26881 15651 26939 15657
rect 27614 15648 27620 15660
rect 27672 15648 27678 15700
rect 15562 15629 15568 15632
rect 15556 15620 15568 15629
rect 15523 15592 15568 15620
rect 15556 15583 15568 15592
rect 15562 15580 15568 15583
rect 15620 15580 15626 15632
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18877 15623 18935 15629
rect 18877 15620 18889 15623
rect 18012 15592 18889 15620
rect 18012 15580 18018 15592
rect 18877 15589 18889 15592
rect 18923 15589 18935 15623
rect 18877 15583 18935 15589
rect 24765 15623 24823 15629
rect 24765 15589 24777 15623
rect 24811 15620 24823 15623
rect 25314 15620 25320 15632
rect 24811 15592 25320 15620
rect 24811 15589 24823 15592
rect 24765 15583 24823 15589
rect 25314 15580 25320 15592
rect 25372 15580 25378 15632
rect 25590 15580 25596 15632
rect 25648 15620 25654 15632
rect 26160 15620 26188 15648
rect 25648 15592 26188 15620
rect 25648 15580 25654 15592
rect 18782 15552 18788 15564
rect 18743 15524 18788 15552
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 22186 15561 22192 15564
rect 22180 15552 22192 15561
rect 22147 15524 22192 15552
rect 22180 15515 22192 15524
rect 22186 15512 22192 15515
rect 22244 15512 22250 15564
rect 25130 15512 25136 15564
rect 25188 15552 25194 15564
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 25188 15524 25237 15552
rect 25188 15512 25194 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25682 15552 25688 15564
rect 25225 15515 25283 15521
rect 25516 15524 25688 15552
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 18966 15484 18972 15496
rect 18927 15456 18972 15484
rect 15289 15447 15347 15453
rect 13504 15388 15148 15416
rect 13504 15376 13510 15388
rect 9548 15320 9720 15348
rect 11333 15351 11391 15357
rect 9548 15308 9554 15320
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11514 15348 11520 15360
rect 11379 15320 11520 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 15304 15348 15332 15447
rect 18966 15444 18972 15456
rect 19024 15484 19030 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19024 15456 19441 15484
rect 19024 15444 19030 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 21910 15484 21916 15496
rect 21871 15456 21916 15484
rect 19429 15447 19487 15453
rect 21910 15444 21916 15456
rect 21968 15444 21974 15496
rect 25038 15444 25044 15496
rect 25096 15484 25102 15496
rect 25516 15493 25544 15524
rect 25682 15512 25688 15524
rect 25740 15552 25746 15564
rect 26418 15552 26424 15564
rect 25740 15524 26424 15552
rect 25740 15512 25746 15524
rect 26418 15512 26424 15524
rect 26476 15512 26482 15564
rect 25317 15487 25375 15493
rect 25317 15484 25329 15487
rect 25096 15456 25329 15484
rect 25096 15444 25102 15456
rect 25317 15453 25329 15456
rect 25363 15453 25375 15487
rect 25317 15447 25375 15453
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26973 15487 27031 15493
rect 26973 15484 26985 15487
rect 26384 15456 26985 15484
rect 26384 15444 26390 15456
rect 26973 15453 26985 15456
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 27522 15484 27528 15496
rect 27203 15456 27528 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 24026 15376 24032 15428
rect 24084 15416 24090 15428
rect 24213 15419 24271 15425
rect 24213 15416 24225 15419
rect 24084 15388 24225 15416
rect 24084 15376 24090 15388
rect 24213 15385 24225 15388
rect 24259 15385 24271 15419
rect 24213 15379 24271 15385
rect 25774 15376 25780 15428
rect 25832 15416 25838 15428
rect 26418 15416 26424 15428
rect 25832 15388 26424 15416
rect 25832 15376 25838 15388
rect 26418 15376 26424 15388
rect 26476 15376 26482 15428
rect 21450 15348 21456 15360
rect 14700 15320 15332 15348
rect 21411 15320 21456 15348
rect 14700 15308 14706 15320
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 23937 15351 23995 15357
rect 23937 15317 23949 15351
rect 23983 15348 23995 15351
rect 24118 15348 24124 15360
rect 23983 15320 24124 15348
rect 23983 15317 23995 15320
rect 23937 15311 23995 15317
rect 24118 15308 24124 15320
rect 24176 15308 24182 15360
rect 26510 15348 26516 15360
rect 26471 15320 26516 15348
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 3145 15147 3203 15153
rect 3145 15113 3157 15147
rect 3191 15144 3203 15147
rect 3510 15144 3516 15156
rect 3191 15116 3516 15144
rect 3191 15113 3203 15116
rect 3145 15107 3203 15113
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7377 15147 7435 15153
rect 7377 15113 7389 15147
rect 7423 15144 7435 15147
rect 8294 15144 8300 15156
rect 7423 15116 8300 15144
rect 7423 15113 7435 15116
rect 7377 15107 7435 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9674 15144 9680 15156
rect 9635 15116 9680 15144
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10781 15147 10839 15153
rect 10781 15144 10793 15147
rect 10008 15116 10793 15144
rect 10008 15104 10014 15116
rect 10781 15113 10793 15116
rect 10827 15113 10839 15147
rect 10781 15107 10839 15113
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 16209 15147 16267 15153
rect 16209 15144 16221 15147
rect 15804 15116 16221 15144
rect 15804 15104 15810 15116
rect 16209 15113 16221 15116
rect 16255 15144 16267 15147
rect 16255 15116 16528 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 10321 15079 10379 15085
rect 10321 15045 10333 15079
rect 10367 15076 10379 15079
rect 10594 15076 10600 15088
rect 10367 15048 10600 15076
rect 10367 15045 10379 15048
rect 10321 15039 10379 15045
rect 10594 15036 10600 15048
rect 10652 15036 10658 15088
rect 14369 15079 14427 15085
rect 14369 15045 14381 15079
rect 14415 15076 14427 15079
rect 15654 15076 15660 15088
rect 14415 15048 15660 15076
rect 14415 15045 14427 15048
rect 14369 15039 14427 15045
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 3988 14980 4261 15008
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 1854 14940 1860 14952
rect 1811 14912 1860 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 2032 14943 2090 14949
rect 2032 14909 2044 14943
rect 2078 14940 2090 14943
rect 2314 14940 2320 14952
rect 2078 14912 2320 14940
rect 2078 14909 2090 14912
rect 2032 14903 2090 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 1946 14804 1952 14816
rect 1719 14776 1952 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 3988 14804 4016 14980
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 4249 14971 4307 14977
rect 9508 14980 11345 15008
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 6914 14940 6920 14952
rect 4120 14912 6920 14940
rect 4120 14900 4126 14912
rect 6914 14900 6920 14912
rect 6972 14940 6978 14952
rect 7650 14940 7656 14952
rect 6972 14912 7656 14940
rect 6972 14900 6978 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 8294 14940 8300 14952
rect 8255 14912 8300 14940
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 4516 14875 4574 14881
rect 4516 14841 4528 14875
rect 4562 14872 4574 14875
rect 4706 14872 4712 14884
rect 4562 14844 4712 14872
rect 4562 14841 4574 14844
rect 4516 14835 4574 14841
rect 4706 14832 4712 14844
rect 4764 14832 4770 14884
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 8542 14875 8600 14881
rect 8542 14872 8554 14875
rect 7984 14844 8554 14872
rect 7984 14832 7990 14844
rect 8542 14841 8554 14844
rect 8588 14872 8600 14875
rect 9508 14872 9536 14980
rect 11333 14977 11345 14980
rect 11379 15008 11391 15011
rect 11514 15008 11520 15020
rect 11379 14980 11520 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 15488 15017 15516 15048
rect 15654 15036 15660 15048
rect 15712 15076 15718 15088
rect 16298 15076 16304 15088
rect 15712 15048 16304 15076
rect 15712 15036 15718 15048
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 16393 15079 16451 15085
rect 16393 15045 16405 15079
rect 16439 15045 16451 15079
rect 16393 15039 16451 15045
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12768 14980 13001 15008
rect 12768 14968 12774 14980
rect 12989 14977 13001 14980
rect 13035 15008 13047 15011
rect 13449 15011 13507 15017
rect 13449 15008 13461 15011
rect 13035 14980 13461 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13449 14977 13461 14980
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 16408 15008 16436 15039
rect 15473 14971 15531 14977
rect 16316 14980 16436 15008
rect 11146 14940 11152 14952
rect 11107 14912 11152 14940
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 11848 14912 11897 14940
rect 11848 14900 11854 14912
rect 11885 14909 11897 14912
rect 11931 14940 11943 14943
rect 12618 14940 12624 14952
rect 11931 14912 12624 14940
rect 11931 14909 11943 14912
rect 11885 14903 11943 14909
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 11238 14872 11244 14884
rect 8588 14844 9536 14872
rect 11199 14844 11244 14872
rect 8588 14841 8600 14844
rect 8542 14835 8600 14841
rect 11238 14832 11244 14844
rect 11296 14832 11302 14884
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 12176 14844 12817 14872
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 3835 14776 4169 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 4157 14773 4169 14776
rect 4203 14804 4215 14807
rect 4982 14804 4988 14816
rect 4203 14776 4988 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5500 14776 5641 14804
rect 5500 14764 5506 14776
rect 5629 14773 5641 14776
rect 5675 14804 5687 14807
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5675 14776 6193 14804
rect 5675 14773 5687 14776
rect 5629 14767 5687 14773
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6181 14767 6239 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7800 14776 8033 14804
rect 7800 14764 7806 14776
rect 8021 14773 8033 14776
rect 8067 14804 8079 14807
rect 8386 14804 8392 14816
rect 8067 14776 8392 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 10778 14804 10784 14816
rect 10735 14776 10784 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 12176 14813 12204 14844
rect 12805 14841 12817 14844
rect 12851 14872 12863 14875
rect 12986 14872 12992 14884
rect 12851 14844 12992 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 14001 14875 14059 14881
rect 14001 14841 14013 14875
rect 14047 14872 14059 14875
rect 15289 14875 15347 14881
rect 15289 14872 15301 14875
rect 14047 14844 15301 14872
rect 14047 14841 14059 14844
rect 14001 14835 14059 14841
rect 15289 14841 15301 14844
rect 15335 14872 15347 14875
rect 16316 14872 16344 14980
rect 16500 14940 16528 15116
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 17773 15147 17831 15153
rect 17773 15144 17785 15147
rect 16632 15116 17785 15144
rect 16632 15104 16638 15116
rect 17773 15113 17785 15116
rect 17819 15144 17831 15147
rect 17862 15144 17868 15156
rect 17819 15116 17868 15144
rect 17819 15113 17831 15116
rect 17773 15107 17831 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 18601 15147 18659 15153
rect 18601 15113 18613 15147
rect 18647 15144 18659 15147
rect 18966 15144 18972 15156
rect 18647 15116 18972 15144
rect 18647 15113 18659 15116
rect 18601 15107 18659 15113
rect 18966 15104 18972 15116
rect 19024 15104 19030 15156
rect 21634 15104 21640 15156
rect 21692 15144 21698 15156
rect 21729 15147 21787 15153
rect 21729 15144 21741 15147
rect 21692 15116 21741 15144
rect 21692 15104 21698 15116
rect 21729 15113 21741 15116
rect 21775 15113 21787 15147
rect 23382 15144 23388 15156
rect 23343 15116 23388 15144
rect 21729 15107 21787 15113
rect 23382 15104 23388 15116
rect 23440 15144 23446 15156
rect 25682 15144 25688 15156
rect 23440 15116 23796 15144
rect 25643 15116 25688 15144
rect 23440 15104 23446 15116
rect 18230 15036 18236 15088
rect 18288 15076 18294 15088
rect 18877 15079 18935 15085
rect 18877 15076 18889 15079
rect 18288 15048 18889 15076
rect 18288 15036 18294 15048
rect 18877 15045 18889 15048
rect 18923 15076 18935 15079
rect 21542 15076 21548 15088
rect 18923 15048 19104 15076
rect 18923 15045 18935 15048
rect 18877 15039 18935 15045
rect 16942 15008 16948 15020
rect 16903 14980 16948 15008
rect 16942 14968 16948 14980
rect 17000 15008 17006 15020
rect 19076 15017 19104 15048
rect 20732 15048 21548 15076
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 17000 14980 17417 15008
rect 17000 14968 17006 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 16850 14940 16856 14952
rect 16500 14912 16856 14940
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 19076 14940 19104 14971
rect 20732 14940 20760 15048
rect 21542 15036 21548 15048
rect 21600 15076 21606 15088
rect 21910 15076 21916 15088
rect 21600 15048 21916 15076
rect 21600 15036 21606 15048
rect 21910 15036 21916 15048
rect 21968 15036 21974 15088
rect 23661 15079 23719 15085
rect 23661 15076 23673 15079
rect 22204 15048 23673 15076
rect 22204 15017 22232 15048
rect 23661 15045 23673 15048
rect 23707 15045 23719 15079
rect 23661 15039 23719 15045
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21315 14980 22201 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22370 15008 22376 15020
rect 22331 14980 22376 15008
rect 22189 14971 22247 14977
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 23768 15008 23796 15116
rect 25682 15104 25688 15116
rect 25740 15104 25746 15156
rect 27522 15104 27528 15156
rect 27580 15144 27586 15156
rect 28077 15147 28135 15153
rect 28077 15144 28089 15147
rect 27580 15116 28089 15144
rect 27580 15104 27586 15116
rect 28077 15113 28089 15116
rect 28123 15113 28135 15147
rect 28077 15107 28135 15113
rect 25590 15036 25596 15088
rect 25648 15076 25654 15088
rect 25961 15079 26019 15085
rect 25961 15076 25973 15079
rect 25648 15048 25973 15076
rect 25648 15036 25654 15048
rect 25961 15045 25973 15048
rect 26007 15076 26019 15079
rect 26007 15048 26188 15076
rect 26007 15045 26019 15048
rect 25961 15039 26019 15045
rect 26160 15017 26188 15048
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23768 14980 24225 15008
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 19076 14912 20760 14940
rect 21450 14900 21456 14952
rect 21508 14940 21514 14952
rect 21818 14940 21824 14952
rect 21508 14912 21824 14940
rect 21508 14900 21514 14912
rect 21818 14900 21824 14912
rect 21876 14940 21882 14952
rect 26418 14949 26424 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 21876 14912 22109 14940
rect 21876 14900 21882 14912
rect 22097 14909 22109 14912
rect 22143 14909 22155 14943
rect 26412 14940 26424 14949
rect 26379 14912 26424 14940
rect 22097 14903 22155 14909
rect 26412 14903 26424 14912
rect 26418 14900 26424 14903
rect 26476 14900 26482 14952
rect 19334 14881 19340 14884
rect 19328 14872 19340 14881
rect 15335 14844 16344 14872
rect 19295 14844 19340 14872
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 19328 14835 19340 14844
rect 19334 14832 19340 14835
rect 19392 14832 19398 14884
rect 20346 14832 20352 14884
rect 20404 14872 20410 14884
rect 21637 14875 21695 14881
rect 21637 14872 21649 14875
rect 20404 14844 21649 14872
rect 20404 14832 20410 14844
rect 21637 14841 21649 14844
rect 21683 14872 21695 14875
rect 21683 14844 21864 14872
rect 21683 14841 21695 14844
rect 21637 14835 21695 14841
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 11940 14776 12173 14804
rect 11940 14764 11946 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12897 14807 12955 14813
rect 12492 14776 12537 14804
rect 12492 14764 12498 14776
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13262 14804 13268 14816
rect 12943 14776 13268 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 14642 14804 14648 14816
rect 14603 14776 14648 14804
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 14829 14807 14887 14813
rect 14829 14773 14841 14807
rect 14875 14804 14887 14807
rect 15010 14804 15016 14816
rect 14875 14776 15016 14804
rect 14875 14773 14887 14776
rect 14829 14767 14887 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15194 14804 15200 14816
rect 15155 14776 15200 14804
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15804 14776 15853 14804
rect 15804 14764 15810 14776
rect 15841 14773 15853 14776
rect 15887 14804 15899 14807
rect 16758 14804 16764 14816
rect 15887 14776 16764 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18230 14804 18236 14816
rect 18095 14776 18236 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 20438 14804 20444 14816
rect 20399 14776 20444 14804
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21836 14804 21864 14844
rect 21910 14832 21916 14884
rect 21968 14872 21974 14884
rect 22741 14875 22799 14881
rect 22741 14872 22753 14875
rect 21968 14844 22753 14872
rect 21968 14832 21974 14844
rect 22741 14841 22753 14844
rect 22787 14841 22799 14875
rect 24026 14872 24032 14884
rect 23987 14844 24032 14872
rect 22741 14835 22799 14841
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 22186 14804 22192 14816
rect 21836 14776 22192 14804
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 24118 14804 24124 14816
rect 24079 14776 24124 14804
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 24949 14807 25007 14813
rect 24949 14773 24961 14807
rect 24995 14804 25007 14807
rect 25038 14804 25044 14816
rect 24995 14776 25044 14804
rect 24995 14773 25007 14776
rect 24949 14767 25007 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 25130 14764 25136 14816
rect 25188 14804 25194 14816
rect 25225 14807 25283 14813
rect 25225 14804 25237 14807
rect 25188 14776 25237 14804
rect 25188 14764 25194 14776
rect 25225 14773 25237 14776
rect 25271 14773 25283 14807
rect 25225 14767 25283 14773
rect 27338 14764 27344 14816
rect 27396 14804 27402 14816
rect 27525 14807 27583 14813
rect 27525 14804 27537 14807
rect 27396 14776 27537 14804
rect 27396 14764 27402 14776
rect 27525 14773 27537 14776
rect 27571 14804 27583 14807
rect 27706 14804 27712 14816
rect 27571 14776 27712 14804
rect 27571 14773 27583 14776
rect 27525 14767 27583 14773
rect 27706 14764 27712 14776
rect 27764 14764 27770 14816
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 2866 14600 2872 14612
rect 2827 14572 2872 14600
rect 2866 14560 2872 14572
rect 2924 14600 2930 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 2924 14572 3801 14600
rect 2924 14560 2930 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 4706 14600 4712 14612
rect 4619 14572 4712 14600
rect 3789 14563 3847 14569
rect 4706 14560 4712 14572
rect 4764 14600 4770 14612
rect 5810 14600 5816 14612
rect 4764 14572 5816 14600
rect 4764 14560 4770 14572
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 8389 14603 8447 14609
rect 8076 14572 8121 14600
rect 8076 14560 8082 14572
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 9490 14600 9496 14612
rect 8435 14572 9496 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 11514 14600 11520 14612
rect 11475 14572 11520 14600
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12342 14600 12348 14612
rect 12207 14572 12348 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 14737 14603 14795 14609
rect 14737 14569 14749 14603
rect 14783 14600 14795 14603
rect 15194 14600 15200 14612
rect 14783 14572 15200 14600
rect 14783 14569 14795 14572
rect 14737 14563 14795 14569
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 15562 14600 15568 14612
rect 15523 14572 15568 14600
rect 15562 14560 15568 14572
rect 15620 14600 15626 14612
rect 16942 14600 16948 14612
rect 15620 14572 16948 14600
rect 15620 14560 15626 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 18417 14603 18475 14609
rect 18417 14569 18429 14603
rect 18463 14600 18475 14603
rect 18782 14600 18788 14612
rect 18463 14572 18788 14600
rect 18463 14569 18475 14572
rect 18417 14563 18475 14569
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19702 14600 19708 14612
rect 19663 14572 19708 14600
rect 19702 14560 19708 14572
rect 19760 14560 19766 14612
rect 20346 14600 20352 14612
rect 20307 14572 20352 14600
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 21266 14560 21272 14612
rect 21324 14600 21330 14612
rect 21361 14603 21419 14609
rect 21361 14600 21373 14603
rect 21324 14572 21373 14600
rect 21324 14560 21330 14572
rect 21361 14569 21373 14572
rect 21407 14569 21419 14603
rect 21361 14563 21419 14569
rect 23474 14560 23480 14612
rect 23532 14600 23538 14612
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 23532 14572 24409 14600
rect 23532 14560 23538 14572
rect 24397 14569 24409 14572
rect 24443 14600 24455 14603
rect 24946 14600 24952 14612
rect 24443 14572 24952 14600
rect 24443 14569 24455 14572
rect 24397 14563 24455 14569
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 25222 14560 25228 14612
rect 25280 14600 25286 14612
rect 25409 14603 25467 14609
rect 25409 14600 25421 14603
rect 25280 14572 25421 14600
rect 25280 14560 25286 14572
rect 25409 14569 25421 14572
rect 25455 14569 25467 14603
rect 25409 14563 25467 14569
rect 26237 14603 26295 14609
rect 26237 14569 26249 14603
rect 26283 14600 26295 14603
rect 26418 14600 26424 14612
rect 26283 14572 26424 14600
rect 26283 14569 26295 14572
rect 26237 14563 26295 14569
rect 26418 14560 26424 14572
rect 26476 14560 26482 14612
rect 26510 14560 26516 14612
rect 26568 14600 26574 14612
rect 26973 14603 27031 14609
rect 26973 14600 26985 14603
rect 26568 14572 26985 14600
rect 26568 14560 26574 14572
rect 26973 14569 26985 14572
rect 27019 14600 27031 14603
rect 28258 14600 28264 14612
rect 27019 14572 28264 14600
rect 27019 14569 27031 14572
rect 26973 14563 27031 14569
rect 28258 14560 28264 14572
rect 28316 14560 28322 14612
rect 1854 14532 1860 14544
rect 1504 14504 1860 14532
rect 1504 14473 1532 14504
rect 1854 14492 1860 14504
rect 1912 14492 1918 14544
rect 5350 14492 5356 14544
rect 5408 14532 5414 14544
rect 5690 14535 5748 14541
rect 5690 14532 5702 14535
rect 5408 14504 5702 14532
rect 5408 14492 5414 14504
rect 5690 14501 5702 14504
rect 5736 14501 5748 14535
rect 5690 14495 5748 14501
rect 7282 14492 7288 14544
rect 7340 14532 7346 14544
rect 10594 14532 10600 14544
rect 7340 14504 10600 14532
rect 7340 14492 7346 14504
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 12529 14535 12587 14541
rect 12529 14501 12541 14535
rect 12575 14532 12587 14535
rect 15105 14535 15163 14541
rect 12575 14504 13308 14532
rect 12575 14501 12587 14504
rect 12529 14495 12587 14501
rect 13280 14476 13308 14504
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 15580 14532 15608 14560
rect 16666 14541 16672 14544
rect 16660 14532 16672 14541
rect 15151 14504 15608 14532
rect 16627 14504 16672 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 16660 14495 16672 14504
rect 16666 14492 16672 14495
rect 16724 14492 16730 14544
rect 24026 14492 24032 14544
rect 24084 14532 24090 14544
rect 24489 14535 24547 14541
rect 24489 14532 24501 14535
rect 24084 14504 24501 14532
rect 24084 14492 24090 14504
rect 24489 14501 24501 14504
rect 24535 14501 24547 14535
rect 24489 14495 24547 14501
rect 25133 14535 25191 14541
rect 25133 14501 25145 14535
rect 25179 14532 25191 14535
rect 25498 14532 25504 14544
rect 25179 14504 25504 14532
rect 25179 14501 25191 14504
rect 25133 14495 25191 14501
rect 25498 14492 25504 14504
rect 25556 14492 25562 14544
rect 27614 14532 27620 14544
rect 27575 14504 27620 14532
rect 27614 14492 27620 14504
rect 27672 14492 27678 14544
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14433 1547 14467
rect 1489 14427 1547 14433
rect 1756 14467 1814 14473
rect 1756 14433 1768 14467
rect 1802 14464 1814 14467
rect 2774 14464 2780 14476
rect 1802 14436 2780 14464
rect 1802 14433 1814 14436
rect 1756 14427 1814 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4246 14464 4252 14476
rect 4111 14436 4252 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9490 14464 9496 14476
rect 8527 14436 9496 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 10410 14473 10416 14476
rect 10404 14464 10416 14473
rect 10371 14436 10416 14464
rect 10404 14427 10416 14436
rect 10410 14424 10416 14427
rect 10468 14424 10474 14476
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 12877 14467 12935 14473
rect 12877 14464 12889 14467
rect 12768 14436 12889 14464
rect 12768 14424 12774 14436
rect 12877 14433 12889 14436
rect 12923 14433 12935 14467
rect 12877 14427 12935 14433
rect 13262 14424 13268 14476
rect 13320 14424 13326 14476
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 18966 14464 18972 14476
rect 18831 14436 18972 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 18966 14424 18972 14436
rect 19024 14464 19030 14476
rect 19426 14464 19432 14476
rect 19024 14436 19432 14464
rect 19024 14424 19030 14436
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19576 14436 19625 14464
rect 19576 14424 19582 14436
rect 19613 14433 19625 14436
rect 19659 14433 19671 14467
rect 19613 14427 19671 14433
rect 21812 14467 21870 14473
rect 21812 14433 21824 14467
rect 21858 14464 21870 14467
rect 22094 14464 22100 14476
rect 21858 14436 22100 14464
rect 21858 14433 21870 14436
rect 21812 14427 21870 14433
rect 22094 14424 22100 14436
rect 22152 14424 22158 14476
rect 26510 14424 26516 14476
rect 26568 14464 26574 14476
rect 26881 14467 26939 14473
rect 26881 14464 26893 14467
rect 26568 14436 26893 14464
rect 26568 14424 26574 14436
rect 26881 14433 26893 14436
rect 26927 14433 26939 14467
rect 26881 14427 26939 14433
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5040 14368 5457 14396
rect 5040 14356 5046 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 8662 14396 8668 14408
rect 8623 14368 8668 14396
rect 5445 14359 5503 14365
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 2924 14232 3433 14260
rect 2924 14220 2930 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 3421 14223 3479 14229
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4249 14263 4307 14269
rect 4249 14260 4261 14263
rect 4120 14232 4261 14260
rect 4120 14220 4126 14232
rect 4249 14229 4261 14232
rect 4295 14229 4307 14263
rect 4249 14223 4307 14229
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5169 14263 5227 14269
rect 5169 14260 5181 14263
rect 5040 14232 5181 14260
rect 5040 14220 5046 14232
rect 5169 14229 5181 14232
rect 5215 14229 5227 14263
rect 5460 14260 5488 14359
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 10134 14396 10140 14408
rect 9048 14368 10140 14396
rect 8294 14328 8300 14340
rect 6380 14300 8300 14328
rect 6380 14272 6408 14300
rect 8294 14288 8300 14300
rect 8352 14328 8358 14340
rect 9048 14337 9076 14368
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 12618 14396 12624 14408
rect 12579 14368 12624 14396
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 16390 14396 16396 14408
rect 14700 14368 16396 14396
rect 14700 14356 14706 14368
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 19886 14396 19892 14408
rect 19847 14368 19892 14396
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 21266 14356 21272 14408
rect 21324 14396 21330 14408
rect 21542 14396 21548 14408
rect 21324 14368 21548 14396
rect 21324 14356 21330 14368
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 27154 14396 27160 14408
rect 27115 14368 27160 14396
rect 24581 14359 24639 14365
rect 9033 14331 9091 14337
rect 9033 14328 9045 14331
rect 8352 14300 9045 14328
rect 8352 14288 8358 14300
rect 9033 14297 9045 14300
rect 9079 14297 9091 14331
rect 13998 14328 14004 14340
rect 13959 14300 14004 14328
rect 9033 14291 9091 14297
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 19153 14331 19211 14337
rect 19153 14297 19165 14331
rect 19199 14328 19211 14331
rect 19334 14328 19340 14340
rect 19199 14300 19340 14328
rect 19199 14297 19211 14300
rect 19153 14291 19211 14297
rect 19334 14288 19340 14300
rect 19392 14328 19398 14340
rect 19392 14300 19748 14328
rect 19392 14288 19398 14300
rect 19720 14272 19748 14300
rect 23198 14288 23204 14340
rect 23256 14328 23262 14340
rect 24029 14331 24087 14337
rect 24029 14328 24041 14331
rect 23256 14300 24041 14328
rect 23256 14288 23262 14300
rect 24029 14297 24041 14300
rect 24075 14297 24087 14331
rect 24596 14328 24624 14359
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 26326 14328 26332 14340
rect 24029 14291 24087 14297
rect 24504 14300 24624 14328
rect 25792 14300 26332 14328
rect 6362 14260 6368 14272
rect 5460 14232 6368 14260
rect 5169 14223 5227 14229
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6788 14232 6837 14260
rect 6788 14220 6794 14232
rect 6825 14229 6837 14232
rect 6871 14229 6883 14263
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 6825 14223 6883 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 19702 14220 19708 14272
rect 19760 14220 19766 14272
rect 22186 14220 22192 14272
rect 22244 14260 22250 14272
rect 22925 14263 22983 14269
rect 22925 14260 22937 14263
rect 22244 14232 22937 14260
rect 22244 14220 22250 14232
rect 22925 14229 22937 14232
rect 22971 14260 22983 14263
rect 23845 14263 23903 14269
rect 23845 14260 23857 14263
rect 22971 14232 23857 14260
rect 22971 14229 22983 14232
rect 22925 14223 22983 14229
rect 23845 14229 23857 14232
rect 23891 14260 23903 14263
rect 24504 14260 24532 14300
rect 25792 14272 25820 14300
rect 26326 14288 26332 14300
rect 26384 14288 26390 14340
rect 26513 14331 26571 14337
rect 26513 14297 26525 14331
rect 26559 14328 26571 14331
rect 26602 14328 26608 14340
rect 26559 14300 26608 14328
rect 26559 14297 26571 14300
rect 26513 14291 26571 14297
rect 26602 14288 26608 14300
rect 26660 14288 26666 14340
rect 25774 14260 25780 14272
rect 23891 14232 24532 14260
rect 25735 14232 25780 14260
rect 23891 14229 23903 14232
rect 23845 14223 23903 14229
rect 25774 14220 25780 14232
rect 25832 14220 25838 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4246 14056 4252 14068
rect 4203 14028 4252 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 5350 14056 5356 14068
rect 4755 14028 5356 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 6638 14056 6644 14068
rect 6551 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14056 6702 14068
rect 7282 14056 7288 14068
rect 6696 14028 7288 14056
rect 6696 14016 6702 14028
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 10686 14056 10692 14068
rect 10647 14028 10692 14056
rect 10686 14016 10692 14028
rect 10744 14056 10750 14068
rect 10744 14028 11192 14056
rect 10744 14016 10750 14028
rect 4338 13948 4344 14000
rect 4396 13988 4402 14000
rect 4985 13991 5043 13997
rect 4985 13988 4997 13991
rect 4396 13960 4997 13988
rect 4396 13948 4402 13960
rect 4985 13957 4997 13960
rect 5031 13988 5043 13991
rect 5534 13988 5540 14000
rect 5031 13960 5540 13988
rect 5031 13957 5043 13960
rect 4985 13951 5043 13957
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 9692 13960 10793 13988
rect 5810 13920 5816 13932
rect 5771 13892 5816 13920
rect 5810 13880 5816 13892
rect 5868 13920 5874 13932
rect 7374 13920 7380 13932
rect 5868 13892 7380 13920
rect 5868 13880 5874 13892
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9692 13929 9720 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9364 13892 9689 13920
rect 9364 13880 9370 13892
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 10410 13920 10416 13932
rect 9907 13892 10416 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 1854 13852 1860 13864
rect 1719 13824 1860 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5040 13824 5641 13852
rect 5040 13812 5046 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6880 13824 7205 13852
rect 6880 13812 6886 13824
rect 7193 13821 7205 13824
rect 7239 13852 7251 13855
rect 7837 13855 7895 13861
rect 7837 13852 7849 13855
rect 7239 13824 7849 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7837 13821 7849 13824
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8662 13852 8668 13864
rect 8343 13824 8668 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8662 13812 8668 13824
rect 8720 13852 8726 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8720 13824 9137 13852
rect 8720 13812 8726 13824
rect 9125 13821 9137 13824
rect 9171 13852 9183 13855
rect 9876 13852 9904 13883
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 11164 13920 11192 14028
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 12124 14028 12173 14056
rect 12124 14016 12130 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 12676 14028 13553 14056
rect 12676 14016 12682 14028
rect 13541 14025 13553 14028
rect 13587 14056 13599 14059
rect 14642 14056 14648 14068
rect 13587 14028 14648 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15013 14059 15071 14065
rect 15013 14025 15025 14059
rect 15059 14056 15071 14059
rect 15194 14056 15200 14068
rect 15059 14028 15200 14056
rect 15059 14025 15071 14028
rect 15013 14019 15071 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 16761 14059 16819 14065
rect 16761 14056 16773 14059
rect 16724 14028 16773 14056
rect 16724 14016 16730 14028
rect 16761 14025 16773 14028
rect 16807 14025 16819 14059
rect 16761 14019 16819 14025
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 18506 14056 18512 14068
rect 17911 14028 18512 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19058 14056 19064 14068
rect 18739 14028 19064 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 20070 14056 20076 14068
rect 20031 14028 20076 14056
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 20254 14056 20260 14068
rect 20215 14028 20260 14056
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 21818 14056 21824 14068
rect 21779 14028 21824 14056
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 24210 14016 24216 14068
rect 24268 14056 24274 14068
rect 24394 14056 24400 14068
rect 24268 14028 24400 14056
rect 24268 14016 24274 14028
rect 24394 14016 24400 14028
rect 24452 14016 24458 14068
rect 26694 14056 26700 14068
rect 26655 14028 26700 14056
rect 26694 14016 26700 14028
rect 26752 14016 26758 14068
rect 27154 14016 27160 14068
rect 27212 14056 27218 14068
rect 27893 14059 27951 14065
rect 27893 14056 27905 14059
rect 27212 14028 27905 14056
rect 27212 14016 27218 14028
rect 27893 14025 27905 14028
rect 27939 14025 27951 14059
rect 28258 14056 28264 14068
rect 28219 14028 28264 14056
rect 27893 14019 27951 14025
rect 28258 14016 28264 14028
rect 28316 14016 28322 14068
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 11164 13892 11345 13920
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11379 13892 11805 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11793 13889 11805 13892
rect 11839 13920 11851 13923
rect 12710 13920 12716 13932
rect 11839 13892 12716 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 12710 13880 12716 13892
rect 12768 13920 12774 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12768 13892 13001 13920
rect 12768 13880 12774 13892
rect 12989 13889 13001 13892
rect 13035 13920 13047 13923
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 13035 13892 13829 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 13817 13883 13875 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 18524 13920 18552 14016
rect 25777 13991 25835 13997
rect 25777 13957 25789 13991
rect 25823 13988 25835 13991
rect 26050 13988 26056 14000
rect 25823 13960 26056 13988
rect 25823 13957 25835 13960
rect 25777 13951 25835 13957
rect 26050 13948 26056 13960
rect 26108 13948 26114 14000
rect 26142 13948 26148 14000
rect 26200 13988 26206 14000
rect 27172 13988 27200 14016
rect 26200 13960 27200 13988
rect 26200 13948 26206 13960
rect 19150 13920 19156 13932
rect 18524 13892 19156 13920
rect 19150 13880 19156 13892
rect 19208 13920 19214 13932
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 19208 13892 19257 13920
rect 19208 13880 19214 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20404 13892 20821 13920
rect 20404 13880 20410 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13920 22523 13923
rect 22646 13920 22652 13932
rect 22511 13892 22652 13920
rect 22511 13889 22523 13892
rect 22465 13883 22523 13889
rect 22646 13880 22652 13892
rect 22704 13880 22710 13932
rect 27338 13880 27344 13932
rect 27396 13920 27402 13932
rect 27525 13923 27583 13929
rect 27525 13920 27537 13923
rect 27396 13892 27537 13920
rect 27396 13880 27402 13892
rect 27525 13889 27537 13892
rect 27571 13920 27583 13923
rect 27614 13920 27620 13932
rect 27571 13892 27620 13920
rect 27571 13889 27583 13892
rect 27525 13883 27583 13889
rect 27614 13880 27620 13892
rect 27672 13880 27678 13932
rect 9171 13824 9904 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10100 13824 11008 13852
rect 10100 13812 10106 13824
rect 2124 13787 2182 13793
rect 2124 13753 2136 13787
rect 2170 13784 2182 13787
rect 2866 13784 2872 13796
rect 2170 13756 2872 13784
rect 2170 13753 2182 13756
rect 2124 13747 2182 13753
rect 2866 13744 2872 13756
rect 2924 13744 2930 13796
rect 5534 13784 5540 13796
rect 5495 13756 5540 13784
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 7282 13784 7288 13796
rect 7243 13756 7288 13784
rect 7282 13744 7288 13756
rect 7340 13744 7346 13796
rect 8757 13787 8815 13793
rect 8757 13753 8769 13787
rect 8803 13784 8815 13787
rect 10980 13784 11008 13824
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 14826 13852 14832 13864
rect 12124 13824 12480 13852
rect 14787 13824 14832 13852
rect 12124 13812 12130 13824
rect 11149 13787 11207 13793
rect 11149 13784 11161 13787
rect 8803 13756 9628 13784
rect 10980 13756 11161 13784
rect 8803 13753 8815 13756
rect 8757 13747 8815 13753
rect 9600 13728 9628 13756
rect 11149 13753 11161 13756
rect 11195 13784 11207 13787
rect 11422 13784 11428 13796
rect 11195 13756 11428 13784
rect 11195 13753 11207 13756
rect 11149 13747 11207 13753
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 12452 13784 12480 13824
rect 14826 13812 14832 13824
rect 14884 13852 14890 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 14884 13824 15485 13852
rect 14884 13812 14890 13824
rect 15473 13821 15485 13824
rect 15519 13852 15531 13855
rect 18506 13852 18512 13864
rect 15519 13824 15608 13852
rect 18467 13824 18512 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 15580 13796 15608 13824
rect 18506 13812 18512 13824
rect 18564 13852 18570 13864
rect 18966 13852 18972 13864
rect 18564 13824 18972 13852
rect 18564 13812 18570 13824
rect 18966 13812 18972 13824
rect 19024 13852 19030 13864
rect 19024 13824 19196 13852
rect 19024 13812 19030 13824
rect 12802 13784 12808 13796
rect 12452 13756 12808 13784
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 15562 13744 15568 13796
rect 15620 13744 15626 13796
rect 19058 13784 19064 13796
rect 19019 13756 19064 13784
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 19168 13793 19196 13824
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19576 13824 19717 13852
rect 19576 13812 19582 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 20070 13812 20076 13864
rect 20128 13852 20134 13864
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 20128 13824 20729 13852
rect 20128 13812 20134 13824
rect 20717 13821 20729 13824
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22152 13824 22845 13852
rect 22152 13812 22158 13824
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 24026 13852 24032 13864
rect 23987 13824 24032 13852
rect 22833 13815 22891 13821
rect 24026 13812 24032 13824
rect 24084 13812 24090 13864
rect 24394 13852 24400 13864
rect 24307 13824 24400 13852
rect 24394 13812 24400 13824
rect 24452 13852 24458 13864
rect 25498 13852 25504 13864
rect 24452 13824 25504 13852
rect 24452 13812 24458 13824
rect 25498 13812 25504 13824
rect 25556 13812 25562 13864
rect 26694 13812 26700 13864
rect 26752 13852 26758 13864
rect 26752 13824 27384 13852
rect 26752 13812 26758 13824
rect 19153 13787 19211 13793
rect 19153 13753 19165 13787
rect 19199 13753 19211 13787
rect 19153 13747 19211 13753
rect 20162 13744 20168 13796
rect 20220 13784 20226 13796
rect 20625 13787 20683 13793
rect 20625 13784 20637 13787
rect 20220 13756 20637 13784
rect 20220 13744 20226 13756
rect 20625 13753 20637 13756
rect 20671 13753 20683 13787
rect 20625 13747 20683 13753
rect 21729 13787 21787 13793
rect 21729 13753 21741 13787
rect 21775 13784 21787 13787
rect 22281 13787 22339 13793
rect 21775 13756 22232 13784
rect 21775 13753 21787 13756
rect 21729 13747 21787 13753
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3237 13719 3295 13725
rect 3237 13716 3249 13719
rect 2832 13688 3249 13716
rect 2832 13676 2838 13688
rect 3237 13685 3249 13688
rect 3283 13685 3295 13719
rect 3237 13679 3295 13685
rect 5169 13719 5227 13725
rect 5169 13685 5181 13719
rect 5215 13716 5227 13719
rect 5350 13716 5356 13728
rect 5215 13688 5356 13716
rect 5215 13685 5227 13688
rect 5169 13679 5227 13685
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 6273 13719 6331 13725
rect 6273 13685 6285 13719
rect 6319 13716 6331 13719
rect 6362 13716 6368 13728
rect 6319 13688 6368 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 9582 13716 9588 13728
rect 9543 13688 9588 13716
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 10192 13688 10333 13716
rect 10192 13676 10198 13688
rect 10321 13685 10333 13688
rect 10367 13716 10379 13719
rect 10502 13716 10508 13728
rect 10367 13688 10508 13716
rect 10367 13685 10379 13688
rect 10321 13679 10379 13685
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 11241 13719 11299 13725
rect 11241 13685 11253 13719
rect 11287 13716 11299 13719
rect 11330 13716 11336 13728
rect 11287 13688 11336 13716
rect 11287 13685 11299 13688
rect 11241 13679 11299 13685
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12492 13688 12537 13716
rect 12492 13676 12498 13688
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 13998 13716 14004 13728
rect 12952 13688 12997 13716
rect 13959 13688 14004 13716
rect 12952 13676 12958 13688
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 14918 13676 14924 13728
rect 14976 13716 14982 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 14976 13688 15393 13716
rect 14976 13676 14982 13688
rect 15381 13685 15393 13688
rect 15427 13685 15439 13719
rect 15381 13679 15439 13685
rect 16390 13676 16396 13728
rect 16448 13716 16454 13728
rect 16485 13719 16543 13725
rect 16485 13716 16497 13719
rect 16448 13688 16497 13716
rect 16448 13676 16454 13688
rect 16485 13685 16497 13688
rect 16531 13716 16543 13719
rect 17126 13716 17132 13728
rect 16531 13688 17132 13716
rect 16531 13685 16543 13688
rect 16485 13679 16543 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 21266 13716 21272 13728
rect 21227 13688 21272 13716
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 22204 13725 22232 13756
rect 22281 13753 22293 13787
rect 22327 13784 22339 13787
rect 23198 13784 23204 13796
rect 22327 13756 23204 13784
rect 22327 13753 22339 13756
rect 22281 13747 22339 13753
rect 23198 13744 23204 13756
rect 23256 13744 23262 13796
rect 23658 13744 23664 13796
rect 23716 13784 23722 13796
rect 24642 13787 24700 13793
rect 24642 13784 24654 13787
rect 23716 13756 24654 13784
rect 23716 13744 23722 13756
rect 24642 13753 24654 13756
rect 24688 13784 24700 13787
rect 24762 13784 24768 13796
rect 24688 13756 24768 13784
rect 24688 13753 24700 13756
rect 24642 13747 24700 13753
rect 24762 13744 24768 13756
rect 24820 13744 24826 13796
rect 26421 13787 26479 13793
rect 26421 13753 26433 13787
rect 26467 13784 26479 13787
rect 27154 13784 27160 13796
rect 26467 13756 27160 13784
rect 26467 13753 26479 13756
rect 26421 13747 26479 13753
rect 27154 13744 27160 13756
rect 27212 13784 27218 13796
rect 27356 13793 27384 13824
rect 27249 13787 27307 13793
rect 27249 13784 27261 13787
rect 27212 13756 27261 13784
rect 27212 13744 27218 13756
rect 27249 13753 27261 13756
rect 27295 13753 27307 13787
rect 27249 13747 27307 13753
rect 27341 13787 27399 13793
rect 27341 13753 27353 13787
rect 27387 13753 27399 13787
rect 27341 13747 27399 13753
rect 22189 13719 22247 13725
rect 22189 13685 22201 13719
rect 22235 13716 22247 13719
rect 22462 13716 22468 13728
rect 22235 13688 22468 13716
rect 22235 13685 22247 13688
rect 22189 13679 22247 13685
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 26878 13716 26884 13728
rect 26839 13688 26884 13716
rect 26878 13676 26884 13688
rect 26936 13676 26942 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 5166 13512 5172 13524
rect 4847 13484 5172 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 5166 13472 5172 13484
rect 5224 13512 5230 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 5224 13484 5273 13512
rect 5224 13472 5230 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 5261 13475 5319 13481
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 5868 13484 5917 13512
rect 5868 13472 5874 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 9306 13512 9312 13524
rect 9267 13484 9312 13512
rect 5905 13475 5963 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 10321 13515 10379 13521
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 10410 13512 10416 13524
rect 10367 13484 10416 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 10735 13484 11161 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 11149 13481 11161 13484
rect 11195 13512 11207 13515
rect 11330 13512 11336 13524
rect 11195 13484 11336 13512
rect 11195 13481 11207 13484
rect 11149 13475 11207 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12308 13484 12633 13512
rect 12308 13472 12314 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13170 13512 13176 13524
rect 13127 13484 13176 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15252 13484 15761 13512
rect 15252 13472 15258 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19886 13512 19892 13524
rect 19383 13484 19892 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20162 13512 20168 13524
rect 20036 13484 20168 13512
rect 20036 13472 20042 13484
rect 20162 13472 20168 13484
rect 20220 13512 20226 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 20220 13484 20269 13512
rect 20220 13472 20226 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 23198 13512 23204 13524
rect 23159 13484 23204 13512
rect 20257 13475 20315 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 23753 13515 23811 13521
rect 23753 13512 23765 13515
rect 23716 13484 23765 13512
rect 23716 13472 23722 13484
rect 23753 13481 23765 13484
rect 23799 13481 23811 13515
rect 25314 13512 25320 13524
rect 25227 13484 25320 13512
rect 23753 13475 23811 13481
rect 25314 13472 25320 13484
rect 25372 13512 25378 13524
rect 26142 13512 26148 13524
rect 25372 13484 26148 13512
rect 25372 13472 25378 13484
rect 26142 13472 26148 13484
rect 26200 13472 26206 13524
rect 26329 13515 26387 13521
rect 26329 13481 26341 13515
rect 26375 13512 26387 13515
rect 26878 13512 26884 13524
rect 26375 13484 26884 13512
rect 26375 13481 26387 13484
rect 26329 13475 26387 13481
rect 26878 13472 26884 13484
rect 26936 13472 26942 13524
rect 27614 13512 27620 13524
rect 27575 13484 27620 13512
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 5408 13416 6285 13444
rect 5408 13404 5414 13416
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 6273 13407 6331 13413
rect 14737 13447 14795 13453
rect 14737 13413 14749 13447
rect 14783 13444 14795 13447
rect 15286 13444 15292 13456
rect 14783 13416 15292 13444
rect 14783 13413 14795 13416
rect 14737 13407 14795 13413
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 16850 13404 16856 13456
rect 16908 13444 16914 13456
rect 17396 13447 17454 13453
rect 17396 13444 17408 13447
rect 16908 13416 17408 13444
rect 16908 13404 16914 13416
rect 17396 13413 17408 13416
rect 17442 13444 17454 13447
rect 17770 13444 17776 13456
rect 17442 13416 17776 13444
rect 17442 13413 17454 13416
rect 17396 13407 17454 13413
rect 17770 13404 17776 13416
rect 17828 13404 17834 13456
rect 19610 13444 19616 13456
rect 19571 13416 19616 13444
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 24394 13444 24400 13456
rect 23952 13416 24400 13444
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 6730 13385 6736 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2464 13348 2513 13376
rect 2464 13336 2470 13348
rect 2501 13345 2513 13348
rect 2547 13376 2559 13379
rect 3513 13379 3571 13385
rect 3513 13376 3525 13379
rect 2547 13348 3525 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3513 13345 3525 13348
rect 3559 13345 3571 13379
rect 6724 13376 6736 13385
rect 6691 13348 6736 13376
rect 3513 13339 3571 13345
rect 6724 13339 6736 13348
rect 6730 13336 6736 13339
rect 6788 13336 6794 13388
rect 11330 13336 11336 13388
rect 11388 13376 11394 13388
rect 11517 13379 11575 13385
rect 11517 13376 11529 13379
rect 11388 13348 11529 13376
rect 11388 13336 11394 13348
rect 11517 13345 11529 13348
rect 11563 13376 11575 13379
rect 12158 13376 12164 13388
rect 11563 13348 12164 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 15010 13336 15016 13388
rect 15068 13376 15074 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15068 13348 15669 13376
rect 15068 13336 15074 13348
rect 15657 13345 15669 13348
rect 15703 13376 15715 13379
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15703 13348 16313 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 21433 13379 21491 13385
rect 21433 13376 21445 13379
rect 20864 13348 21445 13376
rect 20864 13336 20870 13348
rect 21433 13345 21445 13348
rect 21479 13345 21491 13379
rect 21433 13339 21491 13345
rect 23014 13336 23020 13388
rect 23072 13376 23078 13388
rect 23952 13385 23980 13416
rect 24394 13404 24400 13416
rect 24452 13404 24458 13456
rect 23937 13379 23995 13385
rect 23937 13376 23949 13379
rect 23072 13348 23949 13376
rect 23072 13336 23078 13348
rect 23937 13345 23949 13348
rect 23983 13345 23995 13379
rect 23937 13339 23995 13345
rect 24204 13379 24262 13385
rect 24204 13345 24216 13379
rect 24250 13376 24262 13379
rect 24670 13376 24676 13388
rect 24250 13348 24676 13376
rect 24250 13345 24262 13348
rect 24204 13339 24262 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 26050 13336 26056 13388
rect 26108 13376 26114 13388
rect 26108 13348 27200 13376
rect 26108 13336 26114 13348
rect 2590 13308 2596 13320
rect 2551 13280 2596 13308
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13308 2835 13311
rect 2958 13308 2964 13320
rect 2823 13280 2964 13308
rect 2823 13277 2835 13280
rect 2777 13271 2835 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 5258 13268 5264 13320
rect 5316 13308 5322 13320
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5316 13280 5365 13308
rect 5316 13268 5322 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5500 13280 5545 13308
rect 5500 13268 5506 13280
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6420 13280 6469 13308
rect 6420 13268 6426 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 6457 13271 6515 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 13170 13308 13176 13320
rect 13131 13280 13176 13308
rect 11701 13271 11759 13277
rect 4890 13240 4896 13252
rect 4851 13212 4896 13240
rect 4890 13200 4896 13212
rect 4948 13200 4954 13252
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 8757 13243 8815 13249
rect 8757 13240 8769 13243
rect 8260 13212 8769 13240
rect 8260 13200 8266 13212
rect 8757 13209 8769 13212
rect 8803 13209 8815 13243
rect 11514 13240 11520 13252
rect 8757 13203 8815 13209
rect 11072 13212 11520 13240
rect 11072 13184 11100 13212
rect 11514 13200 11520 13212
rect 11572 13240 11578 13252
rect 11716 13240 11744 13271
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20438 13308 20444 13320
rect 19843 13280 20444 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 21174 13308 21180 13320
rect 21135 13280 21180 13308
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 26970 13308 26976 13320
rect 26931 13280 26976 13308
rect 26970 13268 26976 13280
rect 27028 13268 27034 13320
rect 27172 13317 27200 13348
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13308 27215 13311
rect 27522 13308 27528 13320
rect 27203 13280 27528 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 11572 13212 11744 13240
rect 12713 13243 12771 13249
rect 11572 13200 11578 13212
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 12894 13240 12900 13252
rect 12759 13212 12900 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 12894 13200 12900 13212
rect 12952 13240 12958 13252
rect 13725 13243 13783 13249
rect 13725 13240 13737 13243
rect 12952 13212 13737 13240
rect 12952 13200 12958 13212
rect 13725 13209 13737 13212
rect 13771 13209 13783 13243
rect 13725 13203 13783 13209
rect 15289 13243 15347 13249
rect 15289 13209 15301 13243
rect 15335 13240 15347 13243
rect 15378 13240 15384 13252
rect 15335 13212 15384 13240
rect 15335 13209 15347 13212
rect 15289 13203 15347 13209
rect 15378 13200 15384 13212
rect 15436 13200 15442 13252
rect 25961 13243 26019 13249
rect 25961 13209 25973 13243
rect 26007 13240 26019 13243
rect 26510 13240 26516 13252
rect 26007 13212 26516 13240
rect 26007 13209 26019 13212
rect 25961 13203 26019 13209
rect 26510 13200 26516 13212
rect 26568 13200 26574 13252
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2130 13172 2136 13184
rect 2091 13144 2136 13172
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 2832 13144 3157 13172
rect 2832 13132 2838 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 4246 13172 4252 13184
rect 4207 13144 4252 13172
rect 3145 13135 3203 13141
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7248 13144 7849 13172
rect 7248 13132 7254 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 7837 13135 7895 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 9950 13172 9956 13184
rect 9911 13144 9956 13172
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 11054 13172 11060 13184
rect 11015 13144 11060 13172
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 12575 13144 12633 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12621 13141 12633 13144
rect 12667 13172 12679 13175
rect 12802 13172 12808 13184
rect 12667 13144 12808 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 14918 13172 14924 13184
rect 14608 13144 14924 13172
rect 14608 13132 14614 13144
rect 14918 13132 14924 13144
rect 14976 13172 14982 13184
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14976 13144 15025 13172
rect 14976 13132 14982 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 18506 13172 18512 13184
rect 18467 13144 18512 13172
rect 15013 13135 15071 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 22094 13172 22100 13184
rect 21048 13144 22100 13172
rect 21048 13132 21054 13144
rect 22094 13132 22100 13144
rect 22152 13172 22158 13184
rect 22557 13175 22615 13181
rect 22557 13172 22569 13175
rect 22152 13144 22569 13172
rect 22152 13132 22158 13144
rect 22557 13141 22569 13144
rect 22603 13141 22615 13175
rect 22557 13135 22615 13141
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 2648 12940 3985 12968
rect 2648 12928 2654 12940
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 3973 12931 4031 12937
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5074 12968 5080 12980
rect 5031 12940 5080 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5316 12940 6009 12968
rect 5316 12928 5322 12940
rect 5997 12937 6009 12940
rect 6043 12937 6055 12971
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 5997 12931 6055 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 11112 12940 11253 12968
rect 11112 12928 11118 12940
rect 11241 12937 11253 12940
rect 11287 12937 11299 12971
rect 11241 12931 11299 12937
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 12437 12971 12495 12977
rect 12437 12968 12449 12971
rect 11480 12940 12449 12968
rect 11480 12928 11486 12940
rect 12437 12937 12449 12940
rect 12483 12937 12495 12971
rect 12437 12931 12495 12937
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13446 12968 13452 12980
rect 13228 12940 13452 12968
rect 13228 12928 13234 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 14516 12940 14841 12968
rect 14516 12928 14522 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 15010 12968 15016 12980
rect 14971 12940 15016 12968
rect 14829 12931 14887 12937
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3053 12903 3111 12909
rect 3053 12900 3065 12903
rect 2924 12872 3065 12900
rect 2924 12860 2930 12872
rect 3053 12869 3065 12872
rect 3099 12869 3111 12903
rect 3053 12863 3111 12869
rect 4525 12903 4583 12909
rect 4525 12869 4537 12903
rect 4571 12900 4583 12903
rect 4893 12903 4951 12909
rect 4893 12900 4905 12903
rect 4571 12872 4905 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 4893 12869 4905 12872
rect 4939 12900 4951 12903
rect 5442 12900 5448 12912
rect 4939 12872 5448 12900
rect 4939 12869 4951 12872
rect 4893 12863 4951 12869
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 5460 12832 5488 12860
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5460 12804 5549 12832
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 5537 12795 5595 12801
rect 7926 12792 7932 12804
rect 7984 12832 7990 12844
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 7984 12804 8309 12832
rect 7984 12792 7990 12804
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 11572 12804 13093 12832
rect 11572 12792 11578 12804
rect 13081 12801 13093 12804
rect 13127 12832 13139 12835
rect 13354 12832 13360 12844
rect 13127 12804 13360 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13354 12792 13360 12804
rect 13412 12832 13418 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13412 12804 13921 12832
rect 13412 12792 13418 12804
rect 13909 12801 13921 12804
rect 13955 12832 13967 12835
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13955 12804 14197 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 1762 12764 1768 12776
rect 1719 12736 1768 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12764 5411 12767
rect 6822 12764 6828 12776
rect 5399 12736 6828 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7650 12764 7656 12776
rect 7563 12736 7656 12764
rect 7650 12724 7656 12736
rect 7708 12764 7714 12776
rect 8386 12764 8392 12776
rect 7708 12736 8392 12764
rect 7708 12724 7714 12736
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 9861 12767 9919 12773
rect 9861 12764 9873 12767
rect 9815 12736 9873 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 9861 12733 9873 12736
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 1940 12699 1998 12705
rect 1940 12665 1952 12699
rect 1986 12696 1998 12699
rect 2774 12696 2780 12708
rect 1986 12668 2780 12696
rect 1986 12665 1998 12668
rect 1940 12659 1998 12665
rect 2774 12656 2780 12668
rect 2832 12696 2838 12708
rect 2958 12696 2964 12708
rect 2832 12668 2964 12696
rect 2832 12656 2838 12668
rect 2958 12656 2964 12668
rect 3016 12696 3022 12708
rect 3605 12699 3663 12705
rect 3605 12696 3617 12699
rect 3016 12668 3617 12696
rect 3016 12656 3022 12668
rect 3605 12665 3617 12668
rect 3651 12696 3663 12699
rect 3694 12696 3700 12708
rect 3651 12668 3700 12696
rect 3651 12665 3663 12668
rect 3605 12659 3663 12665
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7101 12699 7159 12705
rect 7101 12696 7113 12699
rect 6788 12668 7113 12696
rect 6788 12656 6794 12668
rect 7101 12665 7113 12668
rect 7147 12696 7159 12699
rect 8110 12696 8116 12708
rect 7147 12668 8116 12696
rect 7147 12665 7159 12668
rect 7101 12659 7159 12665
rect 8110 12656 8116 12668
rect 8168 12656 8174 12708
rect 9876 12696 9904 12727
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10117 12767 10175 12773
rect 10117 12764 10129 12767
rect 10008 12736 10129 12764
rect 10008 12724 10014 12736
rect 10117 12733 10129 12736
rect 10163 12733 10175 12767
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 10117 12727 10175 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12764 12955 12767
rect 14274 12764 14280 12776
rect 12943 12736 14280 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 10502 12696 10508 12708
rect 9876 12668 10508 12696
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 12250 12696 12256 12708
rect 12163 12668 12256 12696
rect 12250 12656 12256 12668
rect 12308 12696 12314 12708
rect 12912 12696 12940 12727
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14844 12764 14872 12931
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15896 12940 16037 12968
rect 15896 12928 15902 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16025 12931 16083 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 18782 12968 18788 12980
rect 18647 12940 18788 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 20349 12971 20407 12977
rect 20349 12937 20361 12971
rect 20395 12968 20407 12971
rect 20530 12968 20536 12980
rect 20395 12940 20536 12968
rect 20395 12937 20407 12940
rect 20349 12931 20407 12937
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 21637 12971 21695 12977
rect 21637 12968 21649 12971
rect 20956 12940 21649 12968
rect 20956 12928 20962 12940
rect 21637 12937 21649 12940
rect 21683 12968 21695 12971
rect 21729 12971 21787 12977
rect 21729 12968 21741 12971
rect 21683 12940 21741 12968
rect 21683 12937 21695 12940
rect 21637 12931 21695 12937
rect 21729 12937 21741 12940
rect 21775 12937 21787 12971
rect 21910 12968 21916 12980
rect 21871 12940 21916 12968
rect 21729 12931 21787 12937
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 23014 12968 23020 12980
rect 22975 12940 23020 12968
rect 23014 12928 23020 12940
rect 23072 12968 23078 12980
rect 23385 12971 23443 12977
rect 23385 12968 23397 12971
rect 23072 12940 23397 12968
rect 23072 12928 23078 12940
rect 23385 12937 23397 12940
rect 23431 12968 23443 12971
rect 23566 12968 23572 12980
rect 23431 12940 23572 12968
rect 23431 12937 23443 12940
rect 23385 12931 23443 12937
rect 23566 12928 23572 12940
rect 23624 12928 23630 12980
rect 24394 12928 24400 12980
rect 24452 12968 24458 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 24452 12940 24869 12968
rect 24452 12928 24458 12940
rect 24857 12937 24869 12940
rect 24903 12968 24915 12971
rect 24903 12940 25084 12968
rect 24903 12937 24915 12940
rect 24857 12931 24915 12937
rect 20257 12903 20315 12909
rect 20257 12869 20269 12903
rect 20303 12900 20315 12903
rect 21358 12900 21364 12912
rect 20303 12872 21036 12900
rect 21319 12872 21364 12900
rect 20303 12869 20315 12872
rect 20257 12863 20315 12869
rect 21008 12844 21036 12872
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 24121 12903 24179 12909
rect 24121 12869 24133 12903
rect 24167 12900 24179 12903
rect 24946 12900 24952 12912
rect 24167 12872 24952 12900
rect 24167 12869 24179 12872
rect 24121 12863 24179 12869
rect 24946 12860 24952 12872
rect 25004 12860 25010 12912
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15344 12804 15485 12832
rect 15344 12792 15350 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15654 12832 15660 12844
rect 15615 12804 15660 12832
rect 15473 12795 15531 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 19150 12832 19156 12844
rect 19111 12804 19156 12832
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19208 12804 19625 12832
rect 19208 12792 19214 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 20809 12835 20867 12841
rect 20809 12832 20821 12835
rect 20772 12804 20821 12832
rect 20772 12792 20778 12804
rect 20809 12801 20821 12804
rect 20855 12801 20867 12835
rect 20990 12832 20996 12844
rect 20951 12804 20996 12832
rect 20809 12795 20867 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 14844 12736 15393 12764
rect 15381 12733 15393 12736
rect 15427 12764 15439 12767
rect 16390 12764 16396 12776
rect 15427 12736 16396 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 21376 12764 21404 12860
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 25056 12841 25084 12940
rect 26970 12928 26976 12980
rect 27028 12968 27034 12980
rect 27338 12968 27344 12980
rect 27028 12940 27344 12968
rect 27028 12928 27034 12940
rect 27338 12928 27344 12940
rect 27396 12928 27402 12980
rect 27065 12903 27123 12909
rect 27065 12869 27077 12903
rect 27111 12900 27123 12903
rect 27522 12900 27528 12912
rect 27111 12872 27528 12900
rect 27111 12869 27123 12872
rect 27065 12863 27123 12869
rect 27522 12860 27528 12872
rect 27580 12860 27586 12912
rect 22465 12835 22523 12841
rect 22465 12832 22477 12835
rect 22244 12804 22477 12832
rect 22244 12792 22250 12804
rect 22465 12801 22477 12804
rect 22511 12801 22523 12835
rect 22465 12795 22523 12801
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 22002 12764 22008 12776
rect 21376 12736 22008 12764
rect 22002 12724 22008 12736
rect 22060 12764 22066 12776
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 22060 12736 22293 12764
rect 22060 12724 22066 12736
rect 22281 12733 22293 12736
rect 22327 12733 22339 12767
rect 23934 12764 23940 12776
rect 23895 12736 23940 12764
rect 22281 12727 22339 12733
rect 23934 12724 23940 12736
rect 23992 12764 23998 12776
rect 24489 12767 24547 12773
rect 24489 12764 24501 12767
rect 23992 12736 24501 12764
rect 23992 12724 23998 12736
rect 24489 12733 24501 12736
rect 24535 12764 24547 12767
rect 24854 12764 24860 12776
rect 24535 12736 24860 12764
rect 24535 12733 24547 12736
rect 24489 12727 24547 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25314 12773 25320 12776
rect 25308 12764 25320 12773
rect 25275 12736 25320 12764
rect 25308 12727 25320 12736
rect 25314 12724 25320 12727
rect 25372 12724 25378 12776
rect 27522 12764 27528 12776
rect 27483 12736 27528 12764
rect 27522 12724 27528 12736
rect 27580 12764 27586 12776
rect 28077 12767 28135 12773
rect 28077 12764 28089 12767
rect 27580 12736 28089 12764
rect 27580 12724 27586 12736
rect 28077 12733 28089 12736
rect 28123 12733 28135 12767
rect 28077 12727 28135 12733
rect 12308 12668 12940 12696
rect 12308 12656 12314 12668
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 13538 12696 13544 12708
rect 13412 12668 13544 12696
rect 13412 12656 13418 12668
rect 13538 12656 13544 12668
rect 13596 12656 13602 12708
rect 16758 12696 16764 12708
rect 14568 12668 16764 12696
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 4338 12628 4344 12640
rect 2556 12600 4344 12628
rect 2556 12588 2562 12600
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5445 12631 5503 12637
rect 5445 12628 5457 12631
rect 5408 12600 5457 12628
rect 5408 12588 5414 12600
rect 5445 12597 5457 12600
rect 5491 12597 5503 12631
rect 5445 12591 5503 12597
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 6457 12631 6515 12637
rect 6457 12628 6469 12631
rect 6420 12600 6469 12628
rect 6420 12588 6426 12600
rect 6457 12597 6469 12600
rect 6503 12597 6515 12631
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 6457 12591 6515 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 7742 12628 7748 12640
rect 7703 12600 7748 12628
rect 7742 12588 7748 12600
rect 7800 12628 7806 12640
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 7800 12600 8677 12628
rect 7800 12588 7806 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8665 12591 8723 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11664 12600 11897 12628
rect 11664 12588 11670 12600
rect 11885 12597 11897 12600
rect 11931 12628 11943 12631
rect 14568 12628 14596 12668
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 17862 12696 17868 12708
rect 17775 12668 17868 12696
rect 17862 12656 17868 12668
rect 17920 12696 17926 12708
rect 18969 12699 19027 12705
rect 18969 12696 18981 12699
rect 17920 12668 18981 12696
rect 17920 12656 17926 12668
rect 18969 12665 18981 12668
rect 19015 12696 19027 12699
rect 19794 12696 19800 12708
rect 19015 12668 19800 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 16482 12628 16488 12640
rect 11931 12600 14596 12628
rect 16443 12600 16488 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 17184 12600 17233 12628
rect 17184 12588 17190 12600
rect 17221 12597 17233 12600
rect 17267 12628 17279 12631
rect 17770 12628 17776 12640
rect 17267 12600 17776 12628
rect 17267 12597 17279 12600
rect 17221 12591 17279 12597
rect 17770 12588 17776 12600
rect 17828 12588 17834 12640
rect 18509 12631 18567 12637
rect 18509 12597 18521 12631
rect 18555 12628 18567 12631
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 18555 12600 19073 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 19061 12597 19073 12600
rect 19107 12628 19119 12631
rect 19242 12628 19248 12640
rect 19107 12600 19248 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 20622 12588 20628 12640
rect 20680 12628 20686 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 20680 12600 20729 12628
rect 20680 12588 20686 12600
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 21637 12631 21695 12637
rect 21637 12597 21649 12631
rect 21683 12628 21695 12631
rect 22370 12628 22376 12640
rect 21683 12600 22376 12628
rect 21683 12597 21695 12600
rect 21637 12591 21695 12597
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 26418 12628 26424 12640
rect 26379 12600 26424 12628
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 27709 12631 27767 12637
rect 27709 12597 27721 12631
rect 27755 12628 27767 12631
rect 27798 12628 27804 12640
rect 27755 12600 27804 12628
rect 27755 12597 27767 12600
rect 27709 12591 27767 12597
rect 27798 12588 27804 12600
rect 27856 12588 27862 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 2498 12384 2504 12436
rect 2556 12424 2562 12436
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2556 12396 2789 12424
rect 2556 12384 2562 12396
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 2777 12387 2835 12393
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 6822 12424 6828 12436
rect 6595 12396 6828 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7156 12396 7205 12424
rect 7156 12384 7162 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7558 12424 7564 12436
rect 7471 12396 7564 12424
rect 7193 12387 7251 12393
rect 7558 12384 7564 12396
rect 7616 12424 7622 12436
rect 8202 12424 8208 12436
rect 7616 12396 8208 12424
rect 7616 12384 7622 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 10100 12396 10149 12424
rect 10100 12384 10106 12396
rect 10137 12393 10149 12396
rect 10183 12393 10195 12427
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 10137 12387 10195 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 13265 12427 13323 12433
rect 13265 12424 13277 12427
rect 13136 12396 13277 12424
rect 13136 12384 13142 12396
rect 13265 12393 13277 12396
rect 13311 12393 13323 12427
rect 13265 12387 13323 12393
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 15102 12424 15108 12436
rect 14599 12396 15108 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15565 12427 15623 12433
rect 15565 12393 15577 12427
rect 15611 12424 15623 12427
rect 15654 12424 15660 12436
rect 15611 12396 15660 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16666 12424 16672 12436
rect 16408 12396 16672 12424
rect 1854 12316 1860 12368
rect 1912 12356 1918 12368
rect 1949 12359 2007 12365
rect 1949 12356 1961 12359
rect 1912 12328 1961 12356
rect 1912 12316 1918 12328
rect 1949 12325 1961 12328
rect 1995 12356 2007 12359
rect 6362 12356 6368 12368
rect 1995 12328 6368 12356
rect 1995 12325 2007 12328
rect 1949 12319 2007 12325
rect 6362 12316 6368 12328
rect 6420 12316 6426 12368
rect 11330 12316 11336 12368
rect 11388 12316 11394 12368
rect 11514 12316 11520 12368
rect 11572 12365 11578 12368
rect 11572 12359 11636 12365
rect 11572 12325 11590 12359
rect 11624 12325 11636 12359
rect 11572 12319 11636 12325
rect 11572 12316 11578 12319
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 16408 12356 16436 12396
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20806 12424 20812 12436
rect 20763 12396 20812 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20806 12384 20812 12396
rect 20864 12424 20870 12436
rect 22002 12424 22008 12436
rect 20864 12396 22008 12424
rect 20864 12384 20870 12396
rect 22002 12384 22008 12396
rect 22060 12424 22066 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 22060 12396 22293 12424
rect 22060 12384 22066 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 22281 12387 22339 12393
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24305 12427 24363 12433
rect 24305 12424 24317 12427
rect 24268 12396 24317 12424
rect 24268 12384 24274 12396
rect 24305 12393 24317 12396
rect 24351 12393 24363 12427
rect 24670 12424 24676 12436
rect 24631 12396 24676 12424
rect 24305 12387 24363 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 25314 12384 25320 12436
rect 25372 12424 25378 12436
rect 25869 12427 25927 12433
rect 25869 12424 25881 12427
rect 25372 12396 25881 12424
rect 25372 12384 25378 12396
rect 25869 12393 25881 12396
rect 25915 12393 25927 12427
rect 25869 12387 25927 12393
rect 26513 12427 26571 12433
rect 26513 12393 26525 12427
rect 26559 12424 26571 12427
rect 27338 12424 27344 12436
rect 26559 12396 27344 12424
rect 26559 12393 26571 12396
rect 26513 12387 26571 12393
rect 27338 12384 27344 12396
rect 27396 12384 27402 12436
rect 16758 12356 16764 12368
rect 15436 12328 16436 12356
rect 16719 12328 16764 12356
rect 15436 12316 15442 12328
rect 16758 12316 16764 12328
rect 16816 12316 16822 12368
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 18132 12359 18190 12365
rect 18132 12356 18144 12359
rect 17920 12328 18144 12356
rect 17920 12316 17926 12328
rect 18132 12325 18144 12328
rect 18178 12356 18190 12359
rect 18506 12356 18512 12368
rect 18178 12328 18512 12356
rect 18178 12325 18190 12328
rect 18132 12319 18190 12325
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 21266 12356 21272 12368
rect 20916 12328 21272 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1578 12288 1584 12300
rect 1443 12260 1584 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 4792 12291 4850 12297
rect 4792 12288 4804 12291
rect 2792 12260 4804 12288
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2792 12220 2820 12260
rect 3068 12232 3096 12260
rect 4792 12257 4804 12260
rect 4838 12288 4850 12291
rect 5810 12288 5816 12300
rect 4838 12260 5816 12288
rect 4838 12257 4850 12260
rect 4792 12251 4850 12257
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7340 12260 7665 12288
rect 7340 12248 7346 12260
rect 7653 12257 7665 12260
rect 7699 12288 7711 12291
rect 8202 12288 8208 12300
rect 7699 12260 8208 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10870 12288 10876 12300
rect 10091 12260 10876 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 11348 12288 11376 12316
rect 16666 12288 16672 12300
rect 11287 12260 16672 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 20916 12297 20944 12328
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 22186 12316 22192 12368
rect 22244 12356 22250 12368
rect 22833 12359 22891 12365
rect 22833 12356 22845 12359
rect 22244 12328 22845 12356
rect 22244 12316 22250 12328
rect 22833 12325 22845 12328
rect 22879 12325 22891 12359
rect 22833 12319 22891 12325
rect 23934 12316 23940 12368
rect 23992 12356 23998 12368
rect 24578 12356 24584 12368
rect 23992 12328 24584 12356
rect 23992 12316 23998 12328
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 25406 12356 25412 12368
rect 24780 12328 25412 12356
rect 21174 12297 21180 12300
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12257 20959 12291
rect 21168 12288 21180 12297
rect 21135 12260 21180 12288
rect 20901 12251 20959 12257
rect 21168 12251 21180 12260
rect 21174 12248 21180 12251
rect 21232 12248 21238 12300
rect 23474 12248 23480 12300
rect 23532 12288 23538 12300
rect 23753 12291 23811 12297
rect 23753 12288 23765 12291
rect 23532 12260 23765 12288
rect 23532 12248 23538 12260
rect 23753 12257 23765 12260
rect 23799 12288 23811 12291
rect 24780 12288 24808 12328
rect 25406 12316 25412 12328
rect 25464 12316 25470 12368
rect 23799 12260 24808 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 25130 12248 25136 12300
rect 25188 12288 25194 12300
rect 25225 12291 25283 12297
rect 25225 12288 25237 12291
rect 25188 12260 25237 12288
rect 25188 12248 25194 12260
rect 25225 12257 25237 12260
rect 25271 12257 25283 12291
rect 25225 12251 25283 12257
rect 26510 12248 26516 12300
rect 26568 12288 26574 12300
rect 26881 12291 26939 12297
rect 26881 12288 26893 12291
rect 26568 12260 26893 12288
rect 26568 12248 26574 12260
rect 26881 12257 26893 12260
rect 26927 12257 26939 12291
rect 26881 12251 26939 12257
rect 2363 12192 2820 12220
rect 2869 12223 2927 12229
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 3050 12220 3056 12232
rect 2963 12192 3056 12220
rect 2869 12183 2927 12189
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 2222 12152 2228 12164
rect 1627 12124 2228 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 2884 12152 2912 12183
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 4522 12220 4528 12232
rect 4483 12192 4528 12220
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 7834 12220 7840 12232
rect 7795 12192 7840 12220
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 8573 12223 8631 12229
rect 8573 12220 8585 12223
rect 7984 12192 8585 12220
rect 7984 12180 7990 12192
rect 8573 12189 8585 12192
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10284 12192 10329 12220
rect 10284 12180 10290 12192
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 11330 12220 11336 12232
rect 10560 12192 11336 12220
rect 10560 12180 10566 12192
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 16942 12220 16948 12232
rect 16903 12192 16948 12220
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 17828 12192 17877 12220
rect 17828 12180 17834 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12220 20407 12223
rect 20622 12220 20628 12232
rect 20395 12192 20628 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 25038 12180 25044 12232
rect 25096 12220 25102 12232
rect 25317 12223 25375 12229
rect 25317 12220 25329 12223
rect 25096 12192 25329 12220
rect 25096 12180 25102 12192
rect 25317 12189 25329 12192
rect 25363 12189 25375 12223
rect 25317 12183 25375 12189
rect 25406 12180 25412 12232
rect 25464 12220 25470 12232
rect 25464 12192 25509 12220
rect 25464 12180 25470 12192
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 26973 12223 27031 12229
rect 26973 12220 26985 12223
rect 25740 12192 26985 12220
rect 25740 12180 25746 12192
rect 26973 12189 26985 12192
rect 27019 12189 27031 12223
rect 26973 12183 27031 12189
rect 27157 12223 27215 12229
rect 27157 12189 27169 12223
rect 27203 12220 27215 12223
rect 27614 12220 27620 12232
rect 27203 12192 27620 12220
rect 27203 12189 27215 12192
rect 27157 12183 27215 12189
rect 27614 12180 27620 12192
rect 27672 12220 27678 12232
rect 28074 12220 28080 12232
rect 27672 12192 28080 12220
rect 27672 12180 27678 12192
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 3418 12152 3424 12164
rect 2332 12124 3424 12152
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2332 12084 2360 12124
rect 3418 12112 3424 12124
rect 3476 12112 3482 12164
rect 3513 12155 3571 12161
rect 3513 12121 3525 12155
rect 3559 12152 3571 12155
rect 3694 12152 3700 12164
rect 3559 12124 3700 12152
rect 3559 12121 3571 12124
rect 3513 12115 3571 12121
rect 3694 12112 3700 12124
rect 3752 12152 3758 12164
rect 3752 12124 4476 12152
rect 3752 12112 3758 12124
rect 2096 12056 2360 12084
rect 2409 12087 2467 12093
rect 2096 12044 2102 12056
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 2498 12084 2504 12096
rect 2455 12056 2504 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 4212 12056 4261 12084
rect 4212 12044 4218 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4448 12084 4476 12124
rect 7374 12112 7380 12164
rect 7432 12152 7438 12164
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 7432 12124 9321 12152
rect 7432 12112 7438 12124
rect 9309 12121 9321 12124
rect 9355 12121 9367 12155
rect 9309 12115 9367 12121
rect 16209 12155 16267 12161
rect 16209 12121 16221 12155
rect 16255 12152 16267 12155
rect 16850 12152 16856 12164
rect 16255 12124 16856 12152
rect 16255 12121 16267 12124
rect 16209 12115 16267 12121
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 23661 12155 23719 12161
rect 23661 12121 23673 12155
rect 23707 12152 23719 12155
rect 24578 12152 24584 12164
rect 23707 12124 24584 12152
rect 23707 12121 23719 12124
rect 23661 12115 23719 12121
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 25424 12152 25452 12180
rect 26237 12155 26295 12161
rect 26237 12152 26249 12155
rect 25424 12124 26249 12152
rect 26237 12121 26249 12124
rect 26283 12152 26295 12155
rect 26418 12152 26424 12164
rect 26283 12124 26424 12152
rect 26283 12121 26295 12124
rect 26237 12115 26295 12121
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 5905 12087 5963 12093
rect 5905 12084 5917 12087
rect 4448 12056 5917 12084
rect 4249 12047 4307 12053
rect 5905 12053 5917 12056
rect 5951 12053 5963 12087
rect 7098 12084 7104 12096
rect 7059 12056 7104 12084
rect 5905 12047 5963 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 8938 12084 8944 12096
rect 8899 12056 8944 12084
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9674 12084 9680 12096
rect 9635 12056 9680 12084
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15378 12084 15384 12096
rect 14967 12056 15384 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 16298 12084 16304 12096
rect 16259 12056 16304 12084
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 19208 12056 19257 12084
rect 19208 12044 19214 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 19245 12047 19303 12053
rect 23937 12087 23995 12093
rect 23937 12053 23949 12087
rect 23983 12084 23995 12087
rect 24670 12084 24676 12096
rect 23983 12056 24676 12084
rect 23983 12053 23995 12056
rect 23937 12047 23995 12053
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 24857 12087 24915 12093
rect 24857 12053 24869 12087
rect 24903 12084 24915 12087
rect 26970 12084 26976 12096
rect 24903 12056 26976 12084
rect 24903 12053 24915 12056
rect 24857 12047 24915 12053
rect 26970 12044 26976 12056
rect 27028 12044 27034 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2590 11880 2596 11892
rect 2547 11852 2596 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 4430 11880 4436 11892
rect 4019 11852 4436 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4430 11840 4436 11852
rect 4488 11880 4494 11892
rect 4614 11880 4620 11892
rect 4488 11852 4620 11880
rect 4488 11840 4494 11852
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5166 11880 5172 11892
rect 5127 11852 5172 11880
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7558 11880 7564 11892
rect 7055 11852 7564 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 8113 11883 8171 11889
rect 8113 11880 8125 11883
rect 7892 11852 8125 11880
rect 7892 11840 7898 11852
rect 8113 11849 8125 11852
rect 8159 11880 8171 11883
rect 9950 11880 9956 11892
rect 8159 11852 9956 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10505 11883 10563 11889
rect 10505 11880 10517 11883
rect 10100 11852 10517 11880
rect 10100 11840 10106 11852
rect 10505 11849 10517 11852
rect 10551 11849 10563 11883
rect 10870 11880 10876 11892
rect 10831 11852 10876 11880
rect 10505 11843 10563 11849
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 11572 11852 11713 11880
rect 11572 11840 11578 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 11701 11843 11759 11849
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 12584 11852 14657 11880
rect 12584 11840 12590 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 15933 11883 15991 11889
rect 15933 11849 15945 11883
rect 15979 11880 15991 11883
rect 16666 11880 16672 11892
rect 15979 11852 16672 11880
rect 15979 11849 15991 11852
rect 15933 11843 15991 11849
rect 3234 11812 3240 11824
rect 2976 11784 3240 11812
rect 2976 11753 3004 11784
rect 3234 11772 3240 11784
rect 3292 11772 3298 11824
rect 3694 11772 3700 11824
rect 3752 11812 3758 11824
rect 4249 11815 4307 11821
rect 4249 11812 4261 11815
rect 3752 11784 4261 11812
rect 3752 11772 3758 11784
rect 4249 11781 4261 11784
rect 4295 11781 4307 11815
rect 4249 11775 4307 11781
rect 4709 11815 4767 11821
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 4982 11812 4988 11824
rect 4755 11784 4988 11812
rect 4755 11781 4767 11784
rect 4709 11775 4767 11781
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2961 11747 3019 11753
rect 2961 11744 2973 11747
rect 2455 11716 2973 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2961 11713 2973 11716
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 3050 11704 3056 11756
rect 3108 11744 3114 11756
rect 3108 11716 3153 11744
rect 3108 11704 3114 11716
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4724 11676 4752 11775
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 6420 11784 8309 11812
rect 6420 11772 6426 11784
rect 8297 11781 8309 11784
rect 8343 11812 8355 11815
rect 8389 11815 8447 11821
rect 8389 11812 8401 11815
rect 8343 11784 8401 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 8389 11781 8401 11784
rect 8435 11781 8447 11815
rect 8389 11775 8447 11781
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 11425 11815 11483 11821
rect 11425 11812 11437 11815
rect 11388 11784 11437 11812
rect 11388 11772 11394 11784
rect 11425 11781 11437 11784
rect 11471 11812 11483 11815
rect 12618 11812 12624 11824
rect 11471 11784 12624 11812
rect 11471 11781 11483 11784
rect 11425 11775 11483 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6638 11744 6644 11756
rect 5859 11716 6644 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7156 11716 7573 11744
rect 7156 11704 7162 11716
rect 7561 11713 7573 11716
rect 7607 11744 7619 11747
rect 7926 11744 7932 11756
rect 7607 11716 7932 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 7926 11704 7932 11716
rect 7984 11744 7990 11756
rect 8478 11744 8484 11756
rect 7984 11716 8484 11744
rect 7984 11704 7990 11716
rect 8478 11704 8484 11716
rect 8536 11744 8542 11756
rect 8536 11716 8708 11744
rect 8536 11704 8542 11716
rect 5534 11676 5540 11688
rect 4111 11648 4752 11676
rect 5495 11648 5540 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 8343 11648 8585 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8680 11676 8708 11716
rect 8829 11679 8887 11685
rect 8829 11676 8841 11679
rect 8680 11648 8841 11676
rect 8573 11639 8631 11645
rect 8829 11645 8841 11648
rect 8875 11645 8887 11679
rect 14660 11676 14688 11843
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 17862 11880 17868 11892
rect 17823 11852 17868 11880
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 20772 11852 21465 11880
rect 20772 11840 20778 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 23474 11880 23480 11892
rect 23435 11852 23480 11880
rect 21453 11843 21511 11849
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 25038 11880 25044 11892
rect 24999 11852 25044 11880
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 25682 11880 25688 11892
rect 25643 11852 25688 11880
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 26510 11880 26516 11892
rect 25976 11852 26516 11880
rect 16301 11815 16359 11821
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 16758 11812 16764 11824
rect 16347 11784 16764 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 16758 11772 16764 11784
rect 16816 11772 16822 11824
rect 17696 11784 17908 11812
rect 15378 11744 15384 11756
rect 15339 11716 15384 11744
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 17034 11744 17040 11756
rect 16947 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11744 17098 11756
rect 17402 11744 17408 11756
rect 17092 11716 17408 11744
rect 17092 11704 17098 11716
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14660 11648 15209 11676
rect 8829 11639 8887 11645
rect 15197 11645 15209 11648
rect 15243 11676 15255 11679
rect 17696 11676 17724 11784
rect 17770 11704 17776 11756
rect 17828 11704 17834 11756
rect 17880 11744 17908 11784
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18322 11812 18328 11824
rect 18012 11784 18328 11812
rect 18012 11772 18018 11784
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 20993 11815 21051 11821
rect 20993 11781 21005 11815
rect 21039 11812 21051 11815
rect 21266 11812 21272 11824
rect 21039 11784 21272 11812
rect 21039 11781 21051 11784
rect 20993 11775 21051 11781
rect 18414 11744 18420 11756
rect 17880 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 21008 11744 21036 11775
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 24854 11772 24860 11824
rect 24912 11812 24918 11824
rect 25976 11821 26004 11852
rect 26510 11840 26516 11852
rect 26568 11840 26574 11892
rect 28074 11880 28080 11892
rect 28035 11852 28080 11880
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 25961 11815 26019 11821
rect 25961 11812 25973 11815
rect 24912 11784 25973 11812
rect 24912 11772 24918 11784
rect 25961 11781 25973 11784
rect 26007 11781 26019 11815
rect 25961 11775 26019 11781
rect 22002 11744 22008 11756
rect 19996 11716 21036 11744
rect 21963 11716 22008 11744
rect 15243 11648 17724 11676
rect 17788 11676 17816 11704
rect 18325 11679 18383 11685
rect 18325 11676 18337 11679
rect 17788 11648 18337 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 18325 11645 18337 11648
rect 18371 11676 18383 11679
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18371 11648 18889 11676
rect 18371 11645 18383 11648
rect 18325 11639 18383 11645
rect 18877 11645 18889 11648
rect 18923 11676 18935 11679
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18923 11648 18981 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 18969 11645 18981 11648
rect 19015 11676 19027 11679
rect 19996 11676 20024 11716
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 23750 11704 23756 11756
rect 23808 11744 23814 11756
rect 23845 11747 23903 11753
rect 23845 11744 23857 11747
rect 23808 11716 23857 11744
rect 23808 11704 23814 11716
rect 23845 11713 23857 11716
rect 23891 11713 23903 11747
rect 23845 11707 23903 11713
rect 19015 11648 20024 11676
rect 19015 11645 19027 11648
rect 18969 11639 19027 11645
rect 20530 11636 20536 11688
rect 20588 11676 20594 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 20588 11648 21925 11676
rect 20588 11636 20594 11648
rect 21913 11645 21925 11648
rect 21959 11676 21971 11679
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 21959 11648 22477 11676
rect 21959 11645 21971 11648
rect 21913 11639 21971 11645
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 23860 11676 23888 11707
rect 24210 11704 24216 11756
rect 24268 11744 24274 11756
rect 24489 11747 24547 11753
rect 24489 11744 24501 11747
rect 24268 11716 24501 11744
rect 24268 11704 24274 11716
rect 24489 11713 24501 11716
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 24578 11704 24584 11756
rect 24636 11744 24642 11756
rect 24636 11716 24681 11744
rect 24636 11704 24642 11716
rect 24397 11679 24455 11685
rect 24397 11676 24409 11679
rect 23860 11648 24409 11676
rect 22465 11639 22523 11645
rect 24397 11645 24409 11648
rect 24443 11645 24455 11679
rect 26142 11676 26148 11688
rect 26103 11648 26148 11676
rect 24397 11639 24455 11645
rect 26142 11636 26148 11648
rect 26200 11636 26206 11688
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 2915 11580 3617 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 3605 11577 3617 11580
rect 3651 11608 3663 11611
rect 4246 11608 4252 11620
rect 3651 11580 4252 11608
rect 3651 11577 3663 11580
rect 3605 11571 3663 11577
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 5629 11611 5687 11617
rect 5629 11577 5641 11611
rect 5675 11608 5687 11611
rect 6270 11608 6276 11620
rect 5675 11580 6276 11608
rect 5675 11577 5687 11580
rect 5629 11571 5687 11577
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 8938 11608 8944 11620
rect 7484 11580 8944 11608
rect 7484 11552 7512 11580
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 15289 11611 15347 11617
rect 15289 11608 15301 11611
rect 14608 11580 15301 11608
rect 14608 11568 14614 11580
rect 15289 11577 15301 11580
rect 15335 11577 15347 11611
rect 16850 11608 16856 11620
rect 16763 11580 16856 11608
rect 15289 11571 15347 11577
rect 16850 11568 16856 11580
rect 16908 11608 16914 11620
rect 17770 11608 17776 11620
rect 16908 11580 17776 11608
rect 16908 11568 16914 11580
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 19150 11568 19156 11620
rect 19208 11617 19214 11620
rect 19208 11611 19272 11617
rect 19208 11577 19226 11611
rect 19260 11577 19272 11611
rect 19208 11571 19272 11577
rect 19208 11568 19214 11571
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 21821 11611 21879 11617
rect 21821 11608 21833 11611
rect 20864 11580 21833 11608
rect 20864 11568 20870 11580
rect 21821 11577 21833 11580
rect 21867 11608 21879 11611
rect 22186 11608 22192 11620
rect 21867 11580 22192 11608
rect 21867 11577 21879 11580
rect 21821 11571 21879 11577
rect 22186 11568 22192 11580
rect 22244 11568 22250 11620
rect 25406 11568 25412 11620
rect 25464 11608 25470 11620
rect 26390 11611 26448 11617
rect 26390 11608 26402 11611
rect 25464 11580 26402 11608
rect 25464 11568 25470 11580
rect 26390 11577 26402 11580
rect 26436 11577 26448 11611
rect 26390 11571 26448 11577
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 1544 11512 1593 11540
rect 1544 11500 1550 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1581 11503 1639 11509
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4798 11540 4804 11552
rect 4580 11512 4804 11540
rect 4580 11500 4586 11512
rect 4798 11500 4804 11512
rect 4856 11540 4862 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4856 11512 4997 11540
rect 4856 11500 4862 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 6181 11543 6239 11549
rect 6181 11540 6193 11543
rect 5868 11512 6193 11540
rect 5868 11500 5874 11512
rect 6181 11509 6193 11512
rect 6227 11509 6239 11543
rect 6638 11540 6644 11552
rect 6599 11512 6644 11540
rect 6181 11503 6239 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 7466 11540 7472 11552
rect 7427 11512 7472 11540
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 14826 11540 14832 11552
rect 14787 11512 14832 11540
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 16390 11540 16396 11552
rect 16351 11512 16396 11540
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 16758 11540 16764 11552
rect 16540 11512 16764 11540
rect 16540 11500 16546 11512
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 20349 11543 20407 11549
rect 20349 11540 20361 11543
rect 20220 11512 20361 11540
rect 20220 11500 20226 11512
rect 20349 11509 20361 11512
rect 20395 11540 20407 11543
rect 21266 11540 21272 11552
rect 20395 11512 21272 11540
rect 20395 11509 20407 11512
rect 20349 11503 20407 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 24026 11540 24032 11552
rect 23987 11512 24032 11540
rect 24026 11500 24032 11512
rect 24084 11500 24090 11552
rect 27062 11500 27068 11552
rect 27120 11540 27126 11552
rect 27525 11543 27583 11549
rect 27525 11540 27537 11543
rect 27120 11512 27537 11540
rect 27120 11500 27126 11512
rect 27525 11509 27537 11512
rect 27571 11509 27583 11543
rect 27525 11503 27583 11509
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 1452 11308 1593 11336
rect 1452 11296 1458 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 2406 11336 2412 11348
rect 2367 11308 2412 11336
rect 1581 11299 1639 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 2958 11336 2964 11348
rect 2915 11308 2964 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 4338 11336 4344 11348
rect 3568 11308 4344 11336
rect 3568 11296 3574 11308
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 5629 11339 5687 11345
rect 5629 11305 5641 11339
rect 5675 11336 5687 11339
rect 5810 11336 5816 11348
rect 5675 11308 5816 11336
rect 5675 11305 5687 11308
rect 5629 11299 5687 11305
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 6270 11336 6276 11348
rect 6231 11308 6276 11336
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11336 10103 11339
rect 10410 11336 10416 11348
rect 10091 11308 10416 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14608 11308 14841 11336
rect 14608 11296 14614 11308
rect 14829 11305 14841 11308
rect 14875 11305 14887 11339
rect 14829 11299 14887 11305
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15620 11308 16313 11336
rect 15620 11296 15626 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 16390 11296 16396 11348
rect 16448 11336 16454 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 16448 11308 17325 11336
rect 16448 11296 16454 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 17313 11299 17371 11305
rect 17497 11339 17555 11345
rect 17497 11305 17509 11339
rect 17543 11336 17555 11339
rect 17586 11336 17592 11348
rect 17543 11308 17592 11336
rect 17543 11305 17555 11308
rect 17497 11299 17555 11305
rect 3697 11271 3755 11277
rect 3697 11237 3709 11271
rect 3743 11268 3755 11271
rect 4246 11268 4252 11280
rect 3743 11240 4252 11268
rect 3743 11237 3755 11240
rect 3697 11231 3755 11237
rect 4246 11228 4252 11240
rect 4304 11268 4310 11280
rect 4494 11271 4552 11277
rect 4494 11268 4506 11271
rect 4304 11240 4506 11268
rect 4304 11228 4310 11240
rect 4494 11237 4506 11240
rect 4540 11237 4552 11271
rect 6638 11268 6644 11280
rect 6551 11240 6644 11268
rect 4494 11231 4552 11237
rect 6638 11228 6644 11240
rect 6696 11268 6702 11280
rect 7009 11271 7067 11277
rect 7009 11268 7021 11271
rect 6696 11240 7021 11268
rect 6696 11228 6702 11240
rect 7009 11237 7021 11240
rect 7055 11268 7067 11271
rect 7190 11268 7196 11280
rect 7055 11240 7196 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7190 11228 7196 11240
rect 7248 11268 7254 11280
rect 7368 11271 7426 11277
rect 7368 11268 7380 11271
rect 7248 11240 7380 11268
rect 7248 11228 7254 11240
rect 7368 11237 7380 11240
rect 7414 11268 7426 11271
rect 8018 11268 8024 11280
rect 7414 11240 8024 11268
rect 7414 11237 7426 11240
rect 7368 11231 7426 11237
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 9033 11271 9091 11277
rect 9033 11268 9045 11271
rect 8168 11240 9045 11268
rect 8168 11228 8174 11240
rect 9033 11237 9045 11240
rect 9079 11268 9091 11271
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 9079 11240 9413 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 9401 11237 9413 11240
rect 9447 11268 9459 11271
rect 9582 11268 9588 11280
rect 9447 11240 9588 11268
rect 9447 11237 9459 11240
rect 9401 11231 9459 11237
rect 9582 11228 9588 11240
rect 9640 11268 9646 11280
rect 10226 11268 10232 11280
rect 9640 11240 10232 11268
rect 9640 11228 9646 11240
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 15378 11228 15384 11280
rect 15436 11268 15442 11280
rect 16482 11268 16488 11280
rect 15436 11240 16488 11268
rect 15436 11228 15442 11240
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 16942 11268 16948 11280
rect 16903 11240 16948 11268
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 17328 11268 17356 11299
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 19242 11336 19248 11348
rect 19203 11308 19248 11336
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19610 11336 19616 11348
rect 19571 11308 19616 11336
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 21450 11336 21456 11348
rect 21411 11308 21456 11336
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 21913 11339 21971 11345
rect 21913 11305 21925 11339
rect 21959 11336 21971 11339
rect 22002 11336 22008 11348
rect 21959 11308 22008 11336
rect 21959 11305 21971 11308
rect 21913 11299 21971 11305
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22186 11336 22192 11348
rect 22147 11308 22192 11336
rect 22186 11296 22192 11308
rect 22244 11296 22250 11348
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 23014 11336 23020 11348
rect 22787 11308 23020 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 23014 11296 23020 11308
rect 23072 11336 23078 11348
rect 23937 11339 23995 11345
rect 23937 11336 23949 11339
rect 23072 11308 23949 11336
rect 23072 11296 23078 11308
rect 23937 11305 23949 11308
rect 23983 11305 23995 11339
rect 24394 11336 24400 11348
rect 24355 11308 24400 11336
rect 23937 11299 23995 11305
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 25041 11339 25099 11345
rect 25041 11305 25053 11339
rect 25087 11336 25099 11339
rect 25130 11336 25136 11348
rect 25087 11308 25136 11336
rect 25087 11305 25099 11308
rect 25041 11299 25099 11305
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 25406 11336 25412 11348
rect 25367 11308 25412 11336
rect 25406 11296 25412 11308
rect 25464 11296 25470 11348
rect 26694 11296 26700 11348
rect 26752 11336 26758 11348
rect 26881 11339 26939 11345
rect 26881 11336 26893 11339
rect 26752 11308 26893 11336
rect 26752 11296 26758 11308
rect 26881 11305 26893 11308
rect 26927 11305 26939 11339
rect 26881 11299 26939 11305
rect 26970 11296 26976 11348
rect 27028 11336 27034 11348
rect 27614 11336 27620 11348
rect 27028 11308 27620 11336
rect 27028 11296 27034 11308
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 17865 11271 17923 11277
rect 17865 11268 17877 11271
rect 17328 11240 17877 11268
rect 17865 11237 17877 11240
rect 17911 11237 17923 11271
rect 17865 11231 17923 11237
rect 17954 11228 17960 11280
rect 18012 11268 18018 11280
rect 18012 11240 18057 11268
rect 18012 11228 18018 11240
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3510 11200 3516 11212
rect 2823 11172 3516 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 4798 11200 4804 11212
rect 4264 11172 4804 11200
rect 2314 11132 2320 11144
rect 2227 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 3050 11132 3056 11144
rect 2372 11104 3056 11132
rect 2372 11092 2378 11104
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4264 11141 4292 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 6730 11132 6736 11144
rect 6420 11104 6736 11132
rect 6420 11092 6426 11104
rect 6730 11092 6736 11104
rect 6788 11132 6794 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6788 11104 7113 11132
rect 6788 11092 6794 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10244 11141 10272 11228
rect 18506 11200 18512 11212
rect 15948 11172 18512 11200
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9824 11104 10149 11132
rect 9824 11092 9830 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 9674 11064 9680 11076
rect 9635 11036 9680 11064
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 15948 11073 15976 11172
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19628 11200 19656 11296
rect 19705 11271 19763 11277
rect 19705 11237 19717 11271
rect 19751 11268 19763 11271
rect 19794 11268 19800 11280
rect 19751 11240 19800 11268
rect 19751 11237 19763 11240
rect 19705 11231 19763 11237
rect 19794 11228 19800 11240
rect 19852 11268 19858 11280
rect 19852 11240 22600 11268
rect 19852 11228 19858 11240
rect 19300 11172 19656 11200
rect 21269 11203 21327 11209
rect 19300 11160 19306 11172
rect 21269 11169 21281 11203
rect 21315 11200 21327 11203
rect 21358 11200 21364 11212
rect 21315 11172 21364 11200
rect 21315 11169 21327 11172
rect 21269 11163 21327 11169
rect 21358 11160 21364 11172
rect 21416 11160 21422 11212
rect 22572 11200 22600 11240
rect 22646 11228 22652 11280
rect 22704 11268 22710 11280
rect 22833 11271 22891 11277
rect 22833 11268 22845 11271
rect 22704 11240 22845 11268
rect 22704 11228 22710 11240
rect 22833 11237 22845 11240
rect 22879 11268 22891 11271
rect 24026 11268 24032 11280
rect 22879 11240 24032 11268
rect 22879 11237 22891 11240
rect 22833 11231 22891 11237
rect 24026 11228 24032 11240
rect 24084 11228 24090 11280
rect 26142 11268 26148 11280
rect 24228 11240 26148 11268
rect 22572 11172 23520 11200
rect 16393 11135 16451 11141
rect 16393 11101 16405 11135
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11033 15991 11067
rect 16408 11064 16436 11095
rect 16482 11092 16488 11144
rect 16540 11132 16546 11144
rect 18046 11132 18052 11144
rect 16540 11104 16585 11132
rect 18007 11104 18052 11132
rect 16540 11092 16546 11104
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 20162 11132 20168 11144
rect 19935 11104 20168 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20162 11092 20168 11104
rect 20220 11092 20226 11144
rect 22922 11132 22928 11144
rect 22883 11104 22928 11132
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 23492 11132 23520 11172
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 23661 11203 23719 11209
rect 23661 11200 23673 11203
rect 23624 11172 23673 11200
rect 23624 11160 23630 11172
rect 23661 11169 23673 11172
rect 23707 11200 23719 11203
rect 24228 11200 24256 11240
rect 26142 11228 26148 11240
rect 26200 11228 26206 11280
rect 23707 11172 24256 11200
rect 24305 11203 24363 11209
rect 23707 11169 23719 11172
rect 23661 11163 23719 11169
rect 24305 11169 24317 11203
rect 24351 11200 24363 11203
rect 24762 11200 24768 11212
rect 24351 11172 24768 11200
rect 24351 11169 24363 11172
rect 24305 11163 24363 11169
rect 23845 11135 23903 11141
rect 23845 11132 23857 11135
rect 23492 11104 23857 11132
rect 23845 11101 23857 11104
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 16408 11036 16528 11064
rect 15933 11027 15991 11033
rect 16500 10996 16528 11036
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 18969 11067 19027 11073
rect 18969 11064 18981 11067
rect 17000 11036 18981 11064
rect 17000 11024 17006 11036
rect 18969 11033 18981 11036
rect 19015 11064 19027 11067
rect 19150 11064 19156 11076
rect 19015 11036 19156 11064
rect 19015 11033 19027 11036
rect 18969 11027 19027 11033
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 22373 11067 22431 11073
rect 22373 11033 22385 11067
rect 22419 11064 22431 11067
rect 23382 11064 23388 11076
rect 22419 11036 23388 11064
rect 22419 11033 22431 11036
rect 22373 11027 22431 11033
rect 23382 11024 23388 11036
rect 23440 11024 23446 11076
rect 24320 11064 24348 11163
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 24578 11132 24584 11144
rect 24539 11104 24584 11132
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 27062 11132 27068 11144
rect 27023 11104 27068 11132
rect 27062 11092 27068 11104
rect 27120 11092 27126 11144
rect 23492 11036 24348 11064
rect 16850 10996 16856 11008
rect 16500 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 21174 10996 21180 11008
rect 21135 10968 21180 10996
rect 21174 10956 21180 10968
rect 21232 10956 21238 11008
rect 23106 10956 23112 11008
rect 23164 10996 23170 11008
rect 23492 10996 23520 11036
rect 26326 11024 26332 11076
rect 26384 11064 26390 11076
rect 26513 11067 26571 11073
rect 26513 11064 26525 11067
rect 26384 11036 26525 11064
rect 26384 11024 26390 11036
rect 26513 11033 26525 11036
rect 26559 11033 26571 11067
rect 26513 11027 26571 11033
rect 23164 10968 23520 10996
rect 23845 10999 23903 11005
rect 23164 10956 23170 10968
rect 23845 10965 23857 10999
rect 23891 10996 23903 10999
rect 26602 10996 26608 11008
rect 23891 10968 26608 10996
rect 23891 10965 23903 10968
rect 23845 10959 23903 10965
rect 26602 10956 26608 10968
rect 26660 10956 26666 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 3016 10764 3065 10792
rect 3016 10752 3022 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 3605 10795 3663 10801
rect 3605 10761 3617 10795
rect 3651 10792 3663 10795
rect 3786 10792 3792 10804
rect 3651 10764 3792 10792
rect 3651 10761 3663 10764
rect 3605 10755 3663 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 5166 10792 5172 10804
rect 5127 10764 5172 10792
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6638 10792 6644 10804
rect 6319 10764 6644 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 4614 10724 4620 10736
rect 3804 10696 4620 10724
rect 3804 10668 3832 10696
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 6089 10727 6147 10733
rect 6089 10724 6101 10727
rect 4764 10696 6101 10724
rect 4764 10684 4770 10696
rect 6089 10693 6101 10696
rect 6135 10693 6147 10727
rect 6089 10687 6147 10693
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2774 10656 2780 10668
rect 2731 10628 2780 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3936 10628 4077 10656
rect 3936 10616 3942 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4246 10656 4252 10668
rect 4207 10628 4252 10656
rect 4065 10619 4123 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 5442 10656 5448 10668
rect 4540 10628 5448 10656
rect 3510 10588 3516 10600
rect 3423 10560 3516 10588
rect 3510 10548 3516 10560
rect 3568 10588 3574 10600
rect 4540 10588 4568 10628
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6288 10656 6316 10755
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7432 10764 7481 10792
rect 7432 10752 7438 10764
rect 7469 10761 7481 10764
rect 7515 10761 7527 10795
rect 7469 10755 7527 10761
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8812 10764 8861 10792
rect 8812 10752 8818 10764
rect 8849 10761 8861 10764
rect 8895 10792 8907 10795
rect 8895 10764 9168 10792
rect 8895 10761 8907 10764
rect 8849 10755 8907 10761
rect 8294 10684 8300 10736
rect 8352 10724 8358 10736
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 8352 10696 9045 10724
rect 8352 10684 8358 10696
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 9033 10687 9091 10693
rect 8018 10656 8024 10668
rect 5859 10628 6316 10656
rect 7979 10628 8024 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 3568 10560 4568 10588
rect 3568 10548 3574 10560
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4672 10560 4721 10588
rect 4672 10548 4678 10560
rect 4709 10557 4721 10560
rect 4755 10588 4767 10591
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 4755 10560 5641 10588
rect 4755 10557 4767 10560
rect 4709 10551 4767 10557
rect 5629 10557 5641 10560
rect 5675 10588 5687 10591
rect 6362 10588 6368 10600
rect 5675 10560 6368 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7926 10588 7932 10600
rect 7300 10560 7932 10588
rect 1949 10523 2007 10529
rect 1949 10489 1961 10523
rect 1995 10520 2007 10523
rect 2409 10523 2467 10529
rect 2409 10520 2421 10523
rect 1995 10492 2421 10520
rect 1995 10489 2007 10492
rect 1949 10483 2007 10489
rect 2409 10489 2421 10492
rect 2455 10520 2467 10523
rect 3973 10523 4031 10529
rect 2455 10492 3924 10520
rect 2455 10489 2467 10492
rect 2409 10483 2467 10489
rect 2041 10455 2099 10461
rect 2041 10421 2053 10455
rect 2087 10452 2099 10455
rect 2222 10452 2228 10464
rect 2087 10424 2228 10452
rect 2087 10421 2099 10424
rect 2041 10415 2099 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 3896 10452 3924 10492
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4062 10520 4068 10532
rect 4019 10492 4068 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 7300 10529 7328 10560
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 9140 10588 9168 10764
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15620 10764 15945 10792
rect 15620 10752 15626 10764
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 16482 10792 16488 10804
rect 16439 10764 16488 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 17589 10795 17647 10801
rect 17589 10761 17601 10795
rect 17635 10792 17647 10795
rect 17862 10792 17868 10804
rect 17635 10764 17868 10792
rect 17635 10761 17647 10764
rect 17589 10755 17647 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 18012 10764 18061 10792
rect 18012 10752 18018 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 19153 10795 19211 10801
rect 19153 10761 19165 10795
rect 19199 10792 19211 10795
rect 19242 10792 19248 10804
rect 19199 10764 19248 10792
rect 19199 10761 19211 10764
rect 19153 10755 19211 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 19392 10764 19441 10792
rect 19392 10752 19398 10764
rect 19429 10761 19441 10764
rect 19475 10792 19487 10795
rect 19475 10764 20024 10792
rect 19475 10761 19487 10764
rect 19429 10755 19487 10761
rect 17221 10727 17279 10733
rect 17221 10693 17233 10727
rect 17267 10724 17279 10727
rect 17402 10724 17408 10736
rect 17267 10696 17408 10724
rect 17267 10693 17279 10696
rect 17221 10687 17279 10693
rect 17402 10684 17408 10696
rect 17460 10724 17466 10736
rect 17460 10696 18644 10724
rect 17460 10684 17466 10696
rect 9582 10656 9588 10668
rect 9543 10628 9588 10656
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 18506 10656 18512 10668
rect 18467 10628 18512 10656
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 18616 10665 18644 10696
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9140 10560 9505 10588
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 9493 10551 9551 10557
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 19996 10597 20024 10764
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 20772 10764 21189 10792
rect 20772 10752 20778 10764
rect 21177 10761 21189 10764
rect 21223 10761 21235 10795
rect 21177 10755 21235 10761
rect 22465 10795 22523 10801
rect 22465 10761 22477 10795
rect 22511 10792 22523 10795
rect 22922 10792 22928 10804
rect 22511 10764 22928 10792
rect 22511 10761 22523 10764
rect 22465 10755 22523 10761
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 23106 10792 23112 10804
rect 23067 10764 23112 10792
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 24394 10792 24400 10804
rect 23523 10764 24400 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 26694 10752 26700 10804
rect 26752 10792 26758 10804
rect 27157 10795 27215 10801
rect 27157 10792 27169 10795
rect 26752 10764 27169 10792
rect 26752 10752 26758 10764
rect 27157 10761 27169 10764
rect 27203 10761 27215 10795
rect 27157 10755 27215 10761
rect 27614 10752 27620 10804
rect 27672 10792 27678 10804
rect 27893 10795 27951 10801
rect 27893 10792 27905 10795
rect 27672 10764 27905 10792
rect 27672 10752 27678 10764
rect 27893 10761 27905 10764
rect 27939 10761 27951 10795
rect 27893 10755 27951 10761
rect 21085 10727 21143 10733
rect 21085 10693 21097 10727
rect 21131 10724 21143 10727
rect 21358 10724 21364 10736
rect 21131 10696 21364 10724
rect 21131 10693 21143 10696
rect 21085 10687 21143 10693
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 25314 10684 25320 10736
rect 25372 10724 25378 10736
rect 26145 10727 26203 10733
rect 26145 10724 26157 10727
rect 25372 10696 26157 10724
rect 25372 10684 25378 10696
rect 26145 10693 26157 10696
rect 26191 10693 26203 10727
rect 26145 10687 26203 10693
rect 20162 10656 20168 10668
rect 20075 10628 20168 10656
rect 20162 10616 20168 10628
rect 20220 10656 20226 10668
rect 20714 10656 20720 10668
rect 20220 10628 20720 10656
rect 20220 10616 20226 10628
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 21450 10656 21456 10668
rect 21232 10628 21456 10656
rect 21232 10616 21238 10628
rect 21450 10616 21456 10628
rect 21508 10656 21514 10668
rect 21637 10659 21695 10665
rect 21637 10656 21649 10659
rect 21508 10628 21649 10656
rect 21508 10616 21514 10628
rect 21637 10625 21649 10628
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 21821 10659 21879 10665
rect 21821 10625 21833 10659
rect 21867 10656 21879 10659
rect 22002 10656 22008 10668
rect 21867 10628 22008 10656
rect 21867 10625 21879 10628
rect 21821 10619 21879 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 23566 10616 23572 10668
rect 23624 10656 23630 10668
rect 23661 10659 23719 10665
rect 23661 10656 23673 10659
rect 23624 10628 23673 10656
rect 23624 10616 23630 10628
rect 23661 10625 23673 10628
rect 23707 10625 23719 10659
rect 26697 10659 26755 10665
rect 26697 10656 26709 10659
rect 23661 10619 23719 10625
rect 25608 10628 26709 10656
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 20073 10591 20131 10597
rect 20073 10557 20085 10591
rect 20119 10588 20131 10591
rect 20254 10588 20260 10600
rect 20119 10560 20260 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 6089 10523 6147 10529
rect 4396 10492 5120 10520
rect 4396 10480 4402 10492
rect 4430 10452 4436 10464
rect 2556 10424 2601 10452
rect 3896 10424 4436 10452
rect 2556 10412 2562 10424
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 5092 10461 5120 10492
rect 6089 10489 6101 10523
rect 6135 10520 6147 10523
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 6135 10492 7297 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 7285 10489 7297 10492
rect 7331 10489 7343 10523
rect 7285 10483 7343 10489
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10520 7895 10523
rect 7883 10492 8616 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8588 10464 8616 10492
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 9364 10492 9413 10520
rect 9364 10480 9370 10492
rect 9401 10489 9413 10492
rect 9447 10489 9459 10523
rect 20530 10520 20536 10532
rect 9401 10483 9459 10489
rect 19628 10492 20536 10520
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5534 10452 5540 10464
rect 5123 10424 5540 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 6730 10452 6736 10464
rect 6687 10424 6736 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 8570 10452 8576 10464
rect 8531 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10045 10455 10103 10461
rect 10045 10452 10057 10455
rect 9824 10424 10057 10452
rect 9824 10412 9830 10424
rect 10045 10421 10057 10424
rect 10091 10421 10103 10455
rect 10410 10452 10416 10464
rect 10371 10424 10416 10452
rect 10045 10415 10103 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 16761 10455 16819 10461
rect 16761 10421 16773 10455
rect 16807 10452 16819 10455
rect 16850 10452 16856 10464
rect 16807 10424 16856 10452
rect 16807 10421 16819 10424
rect 16761 10415 16819 10421
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 19628 10461 19656 10492
rect 20530 10480 20536 10492
rect 20588 10480 20594 10532
rect 23474 10480 23480 10532
rect 23532 10520 23538 10532
rect 23928 10523 23986 10529
rect 23928 10520 23940 10523
rect 23532 10492 23940 10520
rect 23532 10480 23538 10492
rect 23928 10489 23940 10492
rect 23974 10520 23986 10523
rect 24578 10520 24584 10532
rect 23974 10492 24584 10520
rect 23974 10489 23986 10492
rect 23928 10483 23986 10489
rect 24578 10480 24584 10492
rect 24636 10520 24642 10532
rect 25608 10529 25636 10628
rect 26697 10625 26709 10628
rect 26743 10656 26755 10659
rect 27062 10656 27068 10668
rect 26743 10628 27068 10656
rect 26743 10625 26755 10628
rect 26697 10619 26755 10625
rect 27062 10616 27068 10628
rect 27120 10656 27126 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27120 10628 27537 10656
rect 27120 10616 27126 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 26602 10588 26608 10600
rect 26563 10560 26608 10588
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 25593 10523 25651 10529
rect 25593 10520 25605 10523
rect 24636 10492 25605 10520
rect 24636 10480 24642 10492
rect 25593 10489 25605 10492
rect 25639 10489 25651 10523
rect 25958 10520 25964 10532
rect 25919 10492 25964 10520
rect 25593 10483 25651 10489
rect 25958 10480 25964 10492
rect 26016 10520 26022 10532
rect 26418 10520 26424 10532
rect 26016 10492 26424 10520
rect 26016 10480 26022 10492
rect 26418 10480 26424 10492
rect 26476 10520 26482 10532
rect 26513 10523 26571 10529
rect 26513 10520 26525 10523
rect 26476 10492 26525 10520
rect 26476 10480 26482 10492
rect 26513 10489 26525 10492
rect 26559 10489 26571 10523
rect 26513 10483 26571 10489
rect 19613 10455 19671 10461
rect 19613 10421 19625 10455
rect 19659 10421 19671 10455
rect 20714 10452 20720 10464
rect 20675 10424 20720 10452
rect 19613 10415 19671 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 21542 10452 21548 10464
rect 21503 10424 21548 10452
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 3418 10248 3424 10260
rect 2823 10220 3424 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3513 10251 3571 10257
rect 3513 10217 3525 10251
rect 3559 10248 3571 10251
rect 4246 10248 4252 10260
rect 3559 10220 4252 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 4246 10208 4252 10220
rect 4304 10248 4310 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 4304 10220 5457 10248
rect 4304 10208 4310 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 4338 10189 4344 10192
rect 4332 10180 4344 10189
rect 4251 10152 4344 10180
rect 4332 10143 4344 10152
rect 4396 10180 4402 10192
rect 7944 10180 7972 10211
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 8260 10220 8493 10248
rect 8260 10208 8266 10220
rect 8481 10217 8493 10220
rect 8527 10217 8539 10251
rect 8481 10211 8539 10217
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 8628 10220 9689 10248
rect 8628 10208 8634 10220
rect 9677 10217 9689 10220
rect 9723 10217 9735 10251
rect 10226 10248 10232 10260
rect 10187 10220 10232 10248
rect 9677 10211 9735 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 17589 10251 17647 10257
rect 17589 10217 17601 10251
rect 17635 10248 17647 10251
rect 18046 10248 18052 10260
rect 17635 10220 18052 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18230 10248 18236 10260
rect 18191 10220 18236 10248
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18472 10220 18889 10248
rect 18472 10208 18478 10220
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 18877 10211 18935 10217
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 21542 10248 21548 10260
rect 20763 10220 21548 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 21726 10208 21732 10260
rect 21784 10248 21790 10260
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 21784 10220 22017 10248
rect 21784 10208 21790 10220
rect 22005 10217 22017 10220
rect 22051 10217 22063 10251
rect 22646 10248 22652 10260
rect 22607 10220 22652 10248
rect 22005 10211 22063 10217
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 23014 10248 23020 10260
rect 22975 10220 23020 10248
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 23474 10248 23480 10260
rect 23435 10220 23480 10248
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 26237 10251 26295 10257
rect 26237 10217 26249 10251
rect 26283 10248 26295 10251
rect 26602 10248 26608 10260
rect 26283 10220 26608 10248
rect 26283 10217 26295 10220
rect 26237 10211 26295 10217
rect 26602 10208 26608 10220
rect 26660 10208 26666 10260
rect 27062 10248 27068 10260
rect 27023 10220 27068 10248
rect 27062 10208 27068 10220
rect 27120 10208 27126 10260
rect 27154 10208 27160 10260
rect 27212 10248 27218 10260
rect 27617 10251 27675 10257
rect 27617 10248 27629 10251
rect 27212 10220 27629 10248
rect 27212 10208 27218 10220
rect 27617 10217 27629 10220
rect 27663 10217 27675 10251
rect 27617 10211 27675 10217
rect 4396 10152 7972 10180
rect 4338 10140 4344 10143
rect 4396 10140 4402 10152
rect 9030 10140 9036 10192
rect 9088 10180 9094 10192
rect 9125 10183 9183 10189
rect 9125 10180 9137 10183
rect 9088 10152 9137 10180
rect 9088 10140 9094 10152
rect 9125 10149 9137 10152
rect 9171 10180 9183 10183
rect 9306 10180 9312 10192
rect 9171 10152 9312 10180
rect 9171 10149 9183 10152
rect 9125 10143 9183 10149
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 18322 10180 18328 10192
rect 17460 10152 18328 10180
rect 17460 10140 17466 10152
rect 18322 10140 18328 10152
rect 18380 10140 18386 10192
rect 19337 10183 19395 10189
rect 19337 10149 19349 10183
rect 19383 10180 19395 10183
rect 19794 10180 19800 10192
rect 19383 10152 19800 10180
rect 19383 10149 19395 10152
rect 19337 10143 19395 10149
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 20438 10140 20444 10192
rect 20496 10180 20502 10192
rect 21910 10180 21916 10192
rect 20496 10152 21916 10180
rect 20496 10140 20502 10152
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 22922 10140 22928 10192
rect 22980 10180 22986 10192
rect 23814 10183 23872 10189
rect 23814 10180 23826 10183
rect 22980 10152 23826 10180
rect 22980 10140 22986 10152
rect 23814 10149 23826 10152
rect 23860 10180 23872 10183
rect 24670 10180 24676 10192
rect 23860 10152 24676 10180
rect 23860 10149 23872 10152
rect 23814 10143 23872 10149
rect 24670 10140 24676 10152
rect 24728 10180 24734 10192
rect 25038 10180 25044 10192
rect 24728 10152 25044 10180
rect 24728 10140 24734 10152
rect 25038 10140 25044 10152
rect 25096 10140 25102 10192
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3326 10112 3332 10124
rect 2915 10084 3332 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 6805 10115 6863 10121
rect 6805 10112 6817 10115
rect 6420 10084 6817 10112
rect 6420 10072 6426 10084
rect 6805 10081 6817 10084
rect 6851 10081 6863 10115
rect 6805 10075 6863 10081
rect 20073 10115 20131 10121
rect 20073 10081 20085 10115
rect 20119 10112 20131 10115
rect 20714 10112 20720 10124
rect 20119 10084 20720 10112
rect 20119 10081 20131 10084
rect 20073 10075 20131 10081
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10112 21327 10115
rect 22002 10112 22008 10124
rect 21315 10084 22008 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 23566 10112 23572 10124
rect 23527 10084 23572 10112
rect 23566 10072 23572 10084
rect 23624 10072 23630 10124
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 1949 10047 2007 10053
rect 1949 10044 1961 10047
rect 1820 10016 1961 10044
rect 1820 10004 1826 10016
rect 1949 10013 1961 10016
rect 1995 10044 2007 10047
rect 2961 10047 3019 10053
rect 1995 10016 2820 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2792 9988 2820 10016
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10044 3939 10047
rect 4062 10044 4068 10056
rect 3927 10016 4068 10044
rect 3927 10013 3939 10016
rect 3881 10007 3939 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 2976 9976 3004 10007
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 3050 9976 3056 9988
rect 2832 9948 3056 9976
rect 2832 9936 2838 9948
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2682 9908 2688 9920
rect 2455 9880 2688 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 6089 9911 6147 9917
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6270 9908 6276 9920
rect 6135 9880 6276 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6564 9908 6592 10007
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 18417 10047 18475 10053
rect 18417 10044 18429 10047
rect 16540 10016 18429 10044
rect 16540 10004 16546 10016
rect 18417 10013 18429 10016
rect 18463 10044 18475 10047
rect 18690 10044 18696 10056
rect 18463 10016 18696 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 22186 10044 22192 10056
rect 22147 10016 22192 10044
rect 22186 10004 22192 10016
rect 22244 10004 22250 10056
rect 16758 9936 16764 9988
rect 16816 9976 16822 9988
rect 17865 9979 17923 9985
rect 17865 9976 17877 9979
rect 16816 9948 17877 9976
rect 16816 9936 16822 9948
rect 17865 9945 17877 9948
rect 17911 9945 17923 9979
rect 17865 9939 17923 9945
rect 6730 9908 6736 9920
rect 6420 9880 6465 9908
rect 6564 9880 6736 9908
rect 6420 9868 6426 9880
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 24946 9908 24952 9920
rect 24907 9880 24952 9908
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 26697 9911 26755 9917
rect 26697 9877 26709 9911
rect 26743 9908 26755 9911
rect 26878 9908 26884 9920
rect 26743 9880 26884 9908
rect 26743 9877 26755 9880
rect 26697 9871 26755 9877
rect 26878 9868 26884 9880
rect 26936 9868 26942 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 1762 9704 1768 9716
rect 1723 9676 1768 9704
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 3326 9704 3332 9716
rect 3287 9676 3332 9704
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 3605 9707 3663 9713
rect 3605 9673 3617 9707
rect 3651 9704 3663 9707
rect 3878 9704 3884 9716
rect 3651 9676 3884 9704
rect 3651 9673 3663 9676
rect 3605 9667 3663 9673
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4062 9664 4068 9716
rect 4120 9664 4126 9716
rect 6454 9704 6460 9716
rect 6380 9676 6460 9704
rect 1857 9639 1915 9645
rect 1857 9605 1869 9639
rect 1903 9636 1915 9639
rect 2406 9636 2412 9648
rect 1903 9608 2412 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 3418 9636 3424 9648
rect 2915 9608 3424 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 4080 9636 4108 9664
rect 4080 9608 4200 9636
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 2188 9540 2329 9568
rect 2188 9528 2194 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2958 9568 2964 9580
rect 2547 9540 2964 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 4172 9500 4200 9608
rect 5258 9596 5264 9648
rect 5316 9636 5322 9648
rect 6380 9636 6408 9676
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 18230 9704 18236 9716
rect 17880 9676 18236 9704
rect 5316 9608 6408 9636
rect 7469 9639 7527 9645
rect 5316 9596 5322 9608
rect 7469 9605 7481 9639
rect 7515 9636 7527 9639
rect 7650 9636 7656 9648
rect 7515 9608 7656 9636
rect 7515 9605 7527 9608
rect 7469 9599 7527 9605
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 7944 9608 8585 9636
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 4338 9568 4344 9580
rect 4295 9540 4344 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4338 9528 4344 9540
rect 4396 9568 4402 9580
rect 4890 9568 4896 9580
rect 4396 9540 4896 9568
rect 4396 9528 4402 9540
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 5810 9568 5816 9580
rect 5771 9540 5816 9568
rect 5810 9528 5816 9540
rect 5868 9568 5874 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5868 9540 6193 9568
rect 5868 9528 5874 9540
rect 6181 9537 6193 9540
rect 6227 9568 6239 9571
rect 6362 9568 6368 9580
rect 6227 9540 6368 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 7944 9577 7972 9608
rect 8573 9605 8585 9608
rect 8619 9636 8631 9639
rect 9582 9636 9588 9648
rect 8619 9608 9588 9636
rect 8619 9605 8631 9608
rect 8573 9599 8631 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17880 9636 17908 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 21450 9664 21456 9716
rect 21508 9704 21514 9716
rect 21545 9707 21603 9713
rect 21545 9704 21557 9707
rect 21508 9676 21557 9704
rect 21508 9664 21514 9676
rect 21545 9673 21557 9676
rect 21591 9673 21603 9707
rect 21545 9667 21603 9673
rect 22922 9664 22928 9716
rect 22980 9704 22986 9716
rect 23017 9707 23075 9713
rect 23017 9704 23029 9707
rect 22980 9676 23029 9704
rect 22980 9664 22986 9676
rect 23017 9673 23029 9676
rect 23063 9673 23075 9707
rect 23017 9667 23075 9673
rect 24762 9664 24768 9716
rect 24820 9664 24826 9716
rect 26329 9707 26387 9713
rect 26329 9673 26341 9707
rect 26375 9704 26387 9707
rect 26694 9704 26700 9716
rect 26375 9676 26700 9704
rect 26375 9673 26387 9676
rect 26329 9667 26387 9673
rect 17175 9608 17908 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 18012 9608 18061 9636
rect 18012 9596 18018 9608
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 18049 9599 18107 9605
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 19610 9636 19616 9648
rect 18196 9608 18552 9636
rect 19571 9608 19616 9636
rect 18196 9596 18202 9608
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 8018 9528 8024 9580
rect 8076 9568 8082 9580
rect 17402 9568 17408 9580
rect 8076 9540 8121 9568
rect 17363 9540 17408 9568
rect 8076 9528 8082 9540
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 17770 9568 17776 9580
rect 17731 9540 17776 9568
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18524 9577 18552 9608
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 21085 9639 21143 9645
rect 21085 9605 21097 9639
rect 21131 9636 21143 9639
rect 21818 9636 21824 9648
rect 21131 9608 21824 9636
rect 21131 9605 21143 9608
rect 21085 9599 21143 9605
rect 21818 9596 21824 9608
rect 21876 9596 21882 9648
rect 23842 9636 23848 9648
rect 23803 9608 23848 9636
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 24780 9636 24808 9664
rect 24780 9608 25452 9636
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9537 18567 9571
rect 18690 9568 18696 9580
rect 18651 9540 18696 9568
rect 18509 9531 18567 9537
rect 18690 9528 18696 9540
rect 18748 9568 18754 9580
rect 19061 9571 19119 9577
rect 19061 9568 19073 9571
rect 18748 9540 19073 9568
rect 18748 9528 18754 9540
rect 19061 9537 19073 9540
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 19702 9528 19708 9580
rect 19760 9568 19766 9580
rect 20165 9571 20223 9577
rect 20165 9568 20177 9571
rect 19760 9540 20177 9568
rect 19760 9528 19766 9540
rect 20165 9537 20177 9540
rect 20211 9537 20223 9571
rect 20714 9568 20720 9580
rect 20627 9540 20720 9568
rect 20165 9531 20223 9537
rect 20714 9528 20720 9540
rect 20772 9568 20778 9580
rect 22186 9568 22192 9580
rect 20772 9540 22192 9568
rect 20772 9528 20778 9540
rect 22186 9528 22192 9540
rect 22244 9568 22250 9580
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22244 9540 22569 9568
rect 22244 9528 22250 9540
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9568 23535 9571
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 23523 9540 24501 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 24489 9537 24501 9540
rect 24535 9568 24547 9571
rect 24762 9568 24768 9580
rect 24535 9540 24768 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 24762 9528 24768 9540
rect 24820 9528 24826 9580
rect 25424 9577 25452 9608
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 4172 9472 4721 9500
rect 4709 9469 4721 9472
rect 4755 9500 4767 9503
rect 4798 9500 4804 9512
rect 4755 9472 4804 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4798 9460 4804 9472
rect 4856 9500 4862 9512
rect 5350 9500 5356 9512
rect 4856 9472 5356 9500
rect 4856 9460 4862 9472
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5500 9472 5549 9500
rect 5500 9460 5506 9472
rect 5537 9469 5549 9472
rect 5583 9500 5595 9503
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 5583 9472 9045 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 9033 9469 9045 9472
rect 9079 9469 9091 9503
rect 17788 9500 17816 9528
rect 18414 9500 18420 9512
rect 17788 9472 18420 9500
rect 9033 9463 9091 9469
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 20070 9500 20076 9512
rect 20031 9472 20076 9500
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 21358 9500 21364 9512
rect 21319 9472 21364 9500
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 21818 9460 21824 9512
rect 21876 9500 21882 9512
rect 26436 9509 26464 9676
rect 26694 9664 26700 9676
rect 26752 9664 26758 9716
rect 26605 9639 26663 9645
rect 26605 9605 26617 9639
rect 26651 9636 26663 9639
rect 26970 9636 26976 9648
rect 26651 9608 26976 9636
rect 26651 9605 26663 9608
rect 26605 9599 26663 9605
rect 26970 9596 26976 9608
rect 27028 9596 27034 9648
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 21876 9472 22017 9500
rect 21876 9460 21882 9472
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9469 26479 9503
rect 26421 9463 26479 9469
rect 26510 9460 26516 9512
rect 26568 9500 26574 9512
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 26568 9472 26985 9500
rect 26568 9460 26574 9472
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 27522 9500 27528 9512
rect 27483 9472 27528 9500
rect 26973 9463 27031 9469
rect 27522 9460 27528 9472
rect 27580 9500 27586 9512
rect 28077 9503 28135 9509
rect 28077 9500 28089 9503
rect 27580 9472 28089 9500
rect 27580 9460 27586 9472
rect 28077 9469 28089 9472
rect 28123 9469 28135 9503
rect 28077 9463 28135 9469
rect 2038 9392 2044 9444
rect 2096 9432 2102 9444
rect 2590 9432 2596 9444
rect 2096 9404 2596 9432
rect 2096 9392 2102 9404
rect 2590 9392 2596 9404
rect 2648 9392 2654 9444
rect 3973 9435 4031 9441
rect 3973 9401 3985 9435
rect 4019 9432 4031 9435
rect 4246 9432 4252 9444
rect 4019 9404 4252 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 4246 9392 4252 9404
rect 4304 9392 4310 9444
rect 4430 9392 4436 9444
rect 4488 9432 4494 9444
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 4488 9404 4997 9432
rect 4488 9392 4494 9404
rect 4985 9401 4997 9404
rect 5031 9432 5043 9435
rect 19521 9435 19579 9441
rect 5031 9404 5672 9432
rect 5031 9401 5043 9404
rect 4985 9395 5043 9401
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5644 9373 5672 9404
rect 19521 9401 19533 9435
rect 19567 9432 19579 9435
rect 20088 9432 20116 9460
rect 19567 9404 20116 9432
rect 21376 9432 21404 9460
rect 21913 9435 21971 9441
rect 21913 9432 21925 9435
rect 21376 9404 21925 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 21913 9401 21925 9404
rect 21959 9401 21971 9435
rect 21913 9395 21971 9401
rect 23474 9392 23480 9444
rect 23532 9432 23538 9444
rect 24213 9435 24271 9441
rect 24213 9432 24225 9435
rect 23532 9404 24225 9432
rect 23532 9392 23538 9404
rect 24213 9401 24225 9404
rect 24259 9432 24271 9435
rect 24857 9435 24915 9441
rect 24857 9432 24869 9435
rect 24259 9404 24869 9432
rect 24259 9401 24271 9404
rect 24213 9395 24271 9401
rect 24857 9401 24869 9404
rect 24903 9401 24915 9435
rect 24857 9395 24915 9401
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 5132 9336 5181 9364
rect 5132 9324 5138 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 5629 9367 5687 9373
rect 5629 9333 5641 9367
rect 5675 9364 5687 9367
rect 5902 9364 5908 9376
rect 5675 9336 5908 9364
rect 5675 9333 5687 9336
rect 5629 9327 5687 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6052 9336 6561 9364
rect 6052 9324 6058 9336
rect 6549 9333 6561 9336
rect 6595 9364 6607 9367
rect 6730 9364 6736 9376
rect 6595 9336 6736 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 7377 9367 7435 9373
rect 7377 9333 7389 9367
rect 7423 9364 7435 9367
rect 7834 9364 7840 9376
rect 7423 9336 7840 9364
rect 7423 9333 7435 9336
rect 7377 9327 7435 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 14734 9364 14740 9376
rect 10836 9336 14740 9364
rect 10836 9324 10842 9336
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 19978 9364 19984 9376
rect 19939 9336 19984 9364
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 24305 9367 24363 9373
rect 24305 9333 24317 9367
rect 24351 9364 24363 9367
rect 24394 9364 24400 9376
rect 24351 9336 24400 9364
rect 24351 9333 24363 9336
rect 24305 9327 24363 9333
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 27706 9364 27712 9376
rect 27667 9336 27712 9364
rect 27706 9324 27712 9336
rect 27764 9324 27770 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2958 9160 2964 9172
rect 1995 9132 2964 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 4212 9132 4353 9160
rect 4212 9120 4218 9132
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 4341 9123 4399 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8018 9160 8024 9172
rect 7975 9132 8024 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 18138 9160 18144 9172
rect 18099 9132 18144 9160
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18509 9163 18567 9169
rect 18509 9129 18521 9163
rect 18555 9160 18567 9163
rect 18690 9160 18696 9172
rect 18555 9132 18696 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 19705 9163 19763 9169
rect 19705 9129 19717 9163
rect 19751 9160 19763 9163
rect 19978 9160 19984 9172
rect 19751 9132 19984 9160
rect 19751 9129 19763 9132
rect 19705 9123 19763 9129
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 21637 9163 21695 9169
rect 21637 9129 21649 9163
rect 21683 9160 21695 9163
rect 21726 9160 21732 9172
rect 21683 9132 21732 9160
rect 21683 9129 21695 9132
rect 21637 9123 21695 9129
rect 21726 9120 21732 9132
rect 21784 9120 21790 9172
rect 21910 9160 21916 9172
rect 21871 9132 21916 9160
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 23566 9160 23572 9172
rect 23527 9132 23572 9160
rect 23566 9120 23572 9132
rect 23624 9120 23630 9172
rect 24029 9163 24087 9169
rect 24029 9129 24041 9163
rect 24075 9160 24087 9163
rect 24394 9160 24400 9172
rect 24075 9132 24400 9160
rect 24075 9129 24087 9132
rect 24029 9123 24087 9129
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 24765 9163 24823 9169
rect 24765 9129 24777 9163
rect 24811 9160 24823 9163
rect 25314 9160 25320 9172
rect 24811 9132 25320 9160
rect 24811 9129 24823 9132
rect 24765 9123 24823 9129
rect 25314 9120 25320 9132
rect 25372 9120 25378 9172
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9092 2375 9095
rect 6172 9095 6230 9101
rect 2363 9064 3740 9092
rect 2363 9061 2375 9064
rect 2317 9055 2375 9061
rect 2777 9027 2835 9033
rect 2777 8993 2789 9027
rect 2823 9024 2835 9027
rect 3142 9024 3148 9036
rect 2823 8996 3148 9024
rect 2823 8993 2835 8996
rect 2777 8987 2835 8993
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 3712 9033 3740 9064
rect 6172 9061 6184 9095
rect 6218 9092 6230 9095
rect 6362 9092 6368 9104
rect 6218 9064 6368 9092
rect 6218 9061 6230 9064
rect 6172 9055 6230 9061
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 24854 9092 24860 9104
rect 24767 9064 24860 9092
rect 24854 9052 24860 9064
rect 24912 9092 24918 9104
rect 26142 9092 26148 9104
rect 24912 9064 26148 9092
rect 24912 9052 24918 9064
rect 26142 9052 26148 9064
rect 26200 9052 26206 9104
rect 3697 9027 3755 9033
rect 3697 8993 3709 9027
rect 3743 9024 3755 9027
rect 4338 9024 4344 9036
rect 3743 8996 4344 9024
rect 3743 8993 3755 8996
rect 3697 8987 3755 8993
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 4982 9024 4988 9036
rect 4755 8996 4988 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5994 9024 6000 9036
rect 5920 8996 6000 9024
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2976 8928 3065 8956
rect 2976 8900 3004 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 2958 8848 2964 8900
rect 3016 8848 3022 8900
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 4816 8888 4844 8919
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 4948 8928 4993 8956
rect 4948 8916 4954 8928
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5920 8965 5948 8996
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5500 8928 5917 8956
rect 5500 8916 5506 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 24670 8916 24676 8968
rect 24728 8956 24734 8968
rect 24949 8959 25007 8965
rect 24949 8956 24961 8959
rect 24728 8928 24961 8956
rect 24728 8916 24734 8928
rect 24949 8925 24961 8928
rect 24995 8925 25007 8959
rect 24949 8919 25007 8925
rect 4764 8860 4844 8888
rect 4764 8848 4770 8860
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2409 8823 2467 8829
rect 2409 8820 2421 8823
rect 2372 8792 2421 8820
rect 2372 8780 2378 8792
rect 2409 8789 2421 8792
rect 2455 8789 2467 8823
rect 5810 8820 5816 8832
rect 5771 8792 5816 8820
rect 2409 8783 2467 8789
rect 5810 8780 5816 8792
rect 5868 8820 5874 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 5868 8792 7297 8820
rect 5868 8780 5874 8792
rect 7285 8789 7297 8792
rect 7331 8820 7343 8823
rect 7374 8820 7380 8832
rect 7331 8792 7380 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8352 8792 8401 8820
rect 8352 8780 8358 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 26694 8820 26700 8832
rect 26655 8792 26700 8820
rect 8389 8783 8447 8789
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1636 8588 1961 8616
rect 1636 8576 1642 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 1949 8579 2007 8585
rect 3050 8576 3056 8588
rect 3108 8616 3114 8628
rect 3108 8588 3832 8616
rect 3108 8576 3114 8588
rect 3142 8508 3148 8560
rect 3200 8548 3206 8560
rect 3605 8551 3663 8557
rect 3605 8548 3617 8551
rect 3200 8520 3617 8548
rect 3200 8508 3206 8520
rect 3605 8517 3617 8520
rect 3651 8517 3663 8551
rect 3804 8548 3832 8588
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6328 8588 6837 8616
rect 6328 8576 6334 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 24489 8619 24547 8625
rect 24489 8585 24501 8619
rect 24535 8616 24547 8619
rect 24670 8616 24676 8628
rect 24535 8588 24676 8616
rect 24535 8585 24547 8588
rect 24489 8579 24547 8585
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25225 8619 25283 8625
rect 25225 8585 25237 8619
rect 25271 8616 25283 8619
rect 25314 8616 25320 8628
rect 25271 8588 25320 8616
rect 25271 8585 25283 8588
rect 25225 8579 25283 8585
rect 25314 8576 25320 8588
rect 25372 8576 25378 8628
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26568 8588 27353 8616
rect 26568 8576 26574 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27706 8616 27712 8628
rect 27667 8588 27712 8616
rect 27341 8579 27399 8585
rect 27706 8576 27712 8588
rect 27764 8576 27770 8628
rect 3804 8520 4200 8548
rect 3605 8511 3663 8517
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2038 8480 2044 8492
rect 1903 8452 2044 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2038 8440 2044 8452
rect 2096 8480 2102 8492
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2096 8452 2513 8480
rect 2096 8440 2102 8452
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 4062 8480 4068 8492
rect 3559 8452 4068 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4172 8489 4200 8520
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 4764 8520 5181 8548
rect 4764 8508 4770 8520
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 5442 8508 5448 8560
rect 5500 8548 5506 8560
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 5500 8520 6193 8548
rect 5500 8508 5506 8520
rect 6181 8517 6193 8520
rect 6227 8517 6239 8551
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 6181 8511 6239 8517
rect 7208 8520 8401 8548
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 4157 8443 4215 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 2314 8412 2320 8424
rect 2275 8384 2320 8412
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 3602 8372 3608 8424
rect 3660 8412 3666 8424
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3660 8384 3985 8412
rect 3660 8372 3666 8384
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 4396 8384 4721 8412
rect 4396 8372 4402 8384
rect 4709 8381 4721 8384
rect 4755 8412 4767 8415
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 4755 8384 5641 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5629 8381 5641 8384
rect 5675 8412 5687 8415
rect 5902 8412 5908 8424
rect 5675 8384 5908 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 7208 8421 7236 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 26602 8548 26608 8560
rect 26563 8520 26608 8548
rect 8389 8511 8447 8517
rect 26602 8508 26608 8520
rect 26660 8508 26666 8560
rect 26786 8508 26792 8560
rect 26844 8548 26850 8560
rect 26973 8551 27031 8557
rect 26973 8548 26985 8551
rect 26844 8520 26985 8548
rect 26844 8508 26850 8520
rect 26973 8517 26985 8520
rect 27019 8517 27031 8551
rect 26973 8511 27031 8517
rect 7374 8480 7380 8492
rect 7335 8452 7380 8480
rect 7374 8440 7380 8452
rect 7432 8480 7438 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7432 8452 7849 8480
rect 7432 8440 7438 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8754 8480 8760 8492
rect 8343 8452 8760 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8754 8440 8760 8452
rect 8812 8480 8818 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8812 8452 8861 8480
rect 8812 8440 8818 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 6880 8384 7205 8412
rect 6880 8372 6886 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8956 8412 8984 8443
rect 8444 8384 8984 8412
rect 8444 8372 8450 8384
rect 25222 8372 25228 8424
rect 25280 8412 25286 8424
rect 25317 8415 25375 8421
rect 25317 8412 25329 8415
rect 25280 8384 25329 8412
rect 25280 8372 25286 8384
rect 25317 8381 25329 8384
rect 25363 8412 25375 8415
rect 25869 8415 25927 8421
rect 25869 8412 25881 8415
rect 25363 8384 25881 8412
rect 25363 8381 25375 8384
rect 25317 8375 25375 8381
rect 25869 8381 25881 8384
rect 25915 8381 25927 8415
rect 25869 8375 25927 8381
rect 26421 8415 26479 8421
rect 26421 8381 26433 8415
rect 26467 8412 26479 8415
rect 26804 8412 26832 8508
rect 27522 8412 27528 8424
rect 26467 8384 26832 8412
rect 27483 8384 27528 8412
rect 26467 8381 26479 8384
rect 26421 8375 26479 8381
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27580 8384 28089 8412
rect 27580 8372 27586 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 2406 8344 2412 8356
rect 2367 8316 2412 8344
rect 2406 8304 2412 8316
rect 2464 8304 2470 8356
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5537 8347 5595 8353
rect 5537 8344 5549 8347
rect 5123 8316 5549 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5537 8313 5549 8316
rect 5583 8344 5595 8347
rect 5718 8344 5724 8356
rect 5583 8316 5724 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6972 8316 7297 8344
rect 6972 8304 6978 8316
rect 7285 8313 7297 8316
rect 7331 8313 7343 8347
rect 7285 8307 7343 8313
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6420 8248 6561 8276
rect 6420 8236 6426 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 8757 8279 8815 8285
rect 8757 8276 8769 8279
rect 8444 8248 8769 8276
rect 8444 8236 8450 8248
rect 8757 8245 8769 8248
rect 8803 8276 8815 8279
rect 9030 8276 9036 8288
rect 8803 8248 9036 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2498 8072 2504 8084
rect 2179 8044 2504 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 2958 8032 2964 8084
rect 3016 8072 3022 8084
rect 3053 8075 3111 8081
rect 3053 8072 3065 8075
rect 3016 8044 3065 8072
rect 3016 8032 3022 8044
rect 3053 8041 3065 8044
rect 3099 8041 3111 8075
rect 3602 8072 3608 8084
rect 3563 8044 3608 8072
rect 3053 8035 3111 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 4304 8044 4997 8072
rect 4304 8032 4310 8044
rect 4985 8041 4997 8044
rect 5031 8072 5043 8075
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 5031 8044 5181 8072
rect 5031 8041 5043 8044
rect 4985 8035 5043 8041
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5316 8044 5549 8072
rect 5316 8032 5322 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 5629 8075 5687 8081
rect 5629 8041 5641 8075
rect 5675 8072 5687 8075
rect 6270 8072 6276 8084
rect 5675 8044 6276 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 6270 8032 6276 8044
rect 6328 8072 6334 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6328 8044 6745 8072
rect 6328 8032 6334 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 25501 8075 25559 8081
rect 25501 8041 25513 8075
rect 25547 8072 25559 8075
rect 25866 8072 25872 8084
rect 25547 8044 25872 8072
rect 25547 8041 25559 8044
rect 25501 8035 25559 8041
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 4890 8004 4896 8016
rect 4755 7976 4896 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 2958 7936 2964 7948
rect 2547 7908 2964 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 4062 7936 4068 7948
rect 4023 7908 4068 7936
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 6822 7936 6828 7948
rect 6319 7908 6828 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7374 7936 7380 7948
rect 7147 7908 7380 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7936 25375 7939
rect 25406 7936 25412 7948
rect 25363 7908 25412 7936
rect 25363 7905 25375 7908
rect 25317 7899 25375 7905
rect 25406 7896 25412 7908
rect 25464 7896 25470 7948
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 27246 7936 27252 7948
rect 26559 7908 27252 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 27246 7896 27252 7908
rect 27304 7896 27310 7948
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 8294 7868 8300 7880
rect 7331 7840 8300 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 4028 7772 4261 7800
rect 4028 7760 4034 7772
rect 4249 7769 4261 7772
rect 4295 7769 4307 7803
rect 4249 7763 4307 7769
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 7300 7800 7328 7831
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 6420 7772 7328 7800
rect 6420 7760 6426 7772
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7732 6610 7744
rect 6914 7732 6920 7744
rect 6604 7704 6920 7732
rect 6604 7692 6610 7704
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 26326 7692 26332 7744
rect 26384 7732 26390 7744
rect 26697 7735 26755 7741
rect 26697 7732 26709 7735
rect 26384 7704 26709 7732
rect 26384 7692 26390 7704
rect 26697 7701 26709 7704
rect 26743 7701 26755 7735
rect 26697 7695 26755 7701
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 1452 7500 2329 7528
rect 1452 7488 1458 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2648 7500 2697 7528
rect 2648 7488 2654 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 2685 7491 2743 7497
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3789 7531 3847 7537
rect 3789 7528 3801 7531
rect 3292 7500 3801 7528
rect 3292 7488 3298 7500
rect 3789 7497 3801 7500
rect 3835 7497 3847 7531
rect 3789 7491 3847 7497
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 4120 7500 4169 7528
rect 4120 7488 4126 7500
rect 4157 7497 4169 7500
rect 4203 7497 4215 7531
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 4157 7491 4215 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6089 7531 6147 7537
rect 6089 7497 6101 7531
rect 6135 7528 6147 7531
rect 6270 7528 6276 7540
rect 6135 7500 6276 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 25406 7528 25412 7540
rect 25367 7500 25412 7528
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 27246 7488 27252 7540
rect 27304 7528 27310 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 27304 7500 27353 7528
rect 27304 7488 27310 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 1578 7460 1584 7472
rect 1539 7432 1584 7460
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4893 7463 4951 7469
rect 4893 7460 4905 7463
rect 4028 7432 4905 7460
rect 4028 7420 4034 7432
rect 4893 7429 4905 7432
rect 4939 7429 4951 7463
rect 27706 7460 27712 7472
rect 27667 7432 27712 7460
rect 4893 7423 4951 7429
rect 27706 7420 27712 7432
rect 27764 7420 27770 7472
rect 2038 7392 2044 7404
rect 1412 7364 2044 7392
rect 1412 7333 1440 7364
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2516 7364 3525 7392
rect 2516 7333 2544 7364
rect 3513 7361 3525 7364
rect 3559 7392 3571 7395
rect 6454 7392 6460 7404
rect 3559 7364 6460 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 2501 7287 2559 7293
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 4580 7296 4721 7324
rect 4580 7284 4586 7296
rect 4709 7293 4721 7296
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 26421 7327 26479 7333
rect 26421 7293 26433 7327
rect 26467 7324 26479 7327
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26467 7296 26985 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 26973 7293 26985 7296
rect 27019 7324 27031 7327
rect 27062 7324 27068 7336
rect 27019 7296 27068 7324
rect 27019 7293 27031 7296
rect 26973 7287 27031 7293
rect 27062 7284 27068 7296
rect 27120 7284 27126 7336
rect 27522 7324 27528 7336
rect 27483 7296 27528 7324
rect 27522 7284 27528 7296
rect 27580 7324 27586 7336
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27580 7296 28089 7324
rect 27580 7284 27586 7296
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3145 7259 3203 7265
rect 3145 7256 3157 7259
rect 3016 7228 3157 7256
rect 3016 7216 3022 7228
rect 3145 7225 3157 7228
rect 3191 7256 3203 7259
rect 4798 7256 4804 7268
rect 3191 7228 4804 7256
rect 3191 7225 3203 7228
rect 3145 7219 3203 7225
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 7101 7259 7159 7265
rect 7101 7225 7113 7259
rect 7147 7256 7159 7259
rect 7190 7256 7196 7268
rect 7147 7228 7196 7256
rect 7147 7225 7159 7228
rect 7101 7219 7159 7225
rect 7190 7216 7196 7228
rect 7248 7256 7254 7268
rect 9674 7256 9680 7268
rect 7248 7228 9680 7256
rect 7248 7216 7254 7228
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6420 7160 6561 7188
rect 6420 7148 6426 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 7374 7188 7380 7200
rect 7335 7160 7380 7188
rect 6549 7151 6607 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 26605 7191 26663 7197
rect 26605 7157 26617 7191
rect 26651 7188 26663 7191
rect 26786 7188 26792 7200
rect 26651 7160 26792 7188
rect 26651 7157 26663 7160
rect 26605 7151 26663 7157
rect 26786 7148 26792 7160
rect 26844 7148 26850 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3053 6987 3111 6993
rect 3053 6984 3065 6987
rect 2924 6956 3065 6984
rect 2924 6944 2930 6956
rect 3053 6953 3065 6956
rect 3099 6953 3111 6987
rect 3602 6984 3608 6996
rect 3563 6956 3608 6984
rect 3053 6947 3111 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 5721 6987 5779 6993
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 6546 6984 6552 6996
rect 5767 6956 6552 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 6089 6919 6147 6925
rect 6089 6885 6101 6919
rect 6135 6916 6147 6919
rect 6270 6916 6276 6928
rect 6135 6888 6276 6916
rect 6135 6885 6147 6888
rect 6089 6879 6147 6885
rect 6270 6876 6276 6888
rect 6328 6916 6334 6928
rect 6730 6916 6736 6928
rect 6328 6888 6736 6916
rect 6328 6876 6334 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1854 6848 1860 6860
rect 1443 6820 1860 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2130 6848 2136 6860
rect 2087 6820 2136 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2280 6820 2329 6848
rect 2280 6808 2286 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2516 6780 2544 6811
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 4062 6848 4068 6860
rect 3568 6820 4068 6848
rect 3568 6808 3574 6820
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4706 6848 4712 6860
rect 4667 6820 4712 6848
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 4982 6848 4988 6860
rect 4943 6820 4988 6848
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 5684 6820 6193 6848
rect 5684 6808 5690 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 27430 6848 27436 6860
rect 26559 6820 27436 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 27430 6808 27436 6820
rect 27488 6808 27494 6860
rect 3418 6780 3424 6792
rect 2516 6752 3424 6780
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 6362 6780 6368 6792
rect 6323 6752 6368 6780
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2004 6684 2697 6712
rect 2004 6672 2010 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 4212 6616 4261 6644
rect 4212 6604 4218 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 26694 6644 26700 6656
rect 26655 6616 26700 6644
rect 4249 6607 4307 6613
rect 26694 6604 26700 6616
rect 26752 6604 26758 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1854 6400 1860 6452
rect 1912 6440 1918 6452
rect 1912 6412 2728 6440
rect 1912 6400 1918 6412
rect 1578 6372 1584 6384
rect 1539 6344 1584 6372
rect 1578 6332 1584 6344
rect 1636 6332 1642 6384
rect 2041 6375 2099 6381
rect 2041 6341 2053 6375
rect 2087 6372 2099 6375
rect 2590 6372 2596 6384
rect 2087 6344 2596 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6335
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 2700 6372 2728 6412
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 4120 6412 4169 6440
rect 4120 6400 4126 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 4157 6403 4215 6409
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5684 6412 5733 6440
rect 5684 6400 5690 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6270 6440 6276 6452
rect 6227 6412 6276 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 26329 6443 26387 6449
rect 26329 6409 26341 6443
rect 26375 6440 26387 6443
rect 26418 6440 26424 6452
rect 26375 6412 26424 6440
rect 26375 6409 26387 6412
rect 26329 6403 26387 6409
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 26602 6440 26608 6452
rect 26563 6412 26608 6440
rect 26602 6400 26608 6412
rect 26660 6400 26666 6452
rect 27065 6443 27123 6449
rect 27065 6409 27077 6443
rect 27111 6440 27123 6443
rect 27430 6440 27436 6452
rect 27111 6412 27436 6440
rect 27111 6409 27123 6412
rect 27065 6403 27123 6409
rect 27430 6400 27436 6412
rect 27488 6400 27494 6452
rect 3326 6372 3332 6384
rect 2700 6344 3332 6372
rect 3326 6332 3332 6344
rect 3384 6332 3390 6384
rect 3418 6332 3424 6384
rect 3476 6372 3482 6384
rect 3513 6375 3571 6381
rect 3513 6372 3525 6375
rect 3476 6344 3525 6372
rect 3476 6332 3482 6344
rect 3513 6341 3525 6344
rect 3559 6372 3571 6375
rect 4430 6372 4436 6384
rect 3559 6344 4436 6372
rect 3559 6341 3571 6344
rect 3513 6335 3571 6341
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 3145 6307 3203 6313
rect 3145 6304 3157 6307
rect 2516 6276 3157 6304
rect 2516 6245 2544 6276
rect 3145 6273 3157 6276
rect 3191 6304 3203 6307
rect 3234 6304 3240 6316
rect 3191 6276 3240 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 1443 6208 2084 6236
rect 2501 6239 2559 6245
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 3602 6236 3608 6248
rect 3515 6208 3608 6236
rect 2501 6199 2559 6205
rect 3602 6196 3608 6208
rect 3660 6236 3666 6248
rect 3786 6236 3792 6248
rect 3660 6208 3792 6236
rect 3660 6196 3666 6208
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 26418 6236 26424 6248
rect 26379 6208 26424 6236
rect 26418 6196 26424 6208
rect 26476 6196 26482 6248
rect 1412 6140 2728 6168
rect 1412 6112 1440 6140
rect 1394 6060 1400 6112
rect 1452 6060 1458 6112
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2700 6109 2728 6140
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 1912 6072 2329 6100
rect 1912 6060 1918 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2317 6063 2375 6069
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6069 2743 6103
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 2685 6063 2743 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 6420 6072 6561 6100
rect 6420 6060 6426 6072
rect 6549 6069 6561 6072
rect 6595 6100 6607 6103
rect 8294 6100 8300 6112
rect 6595 6072 8300 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3602 5896 3608 5908
rect 3563 5868 3608 5896
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5828 2099 5831
rect 2406 5828 2412 5840
rect 2087 5800 2412 5828
rect 2087 5797 2099 5800
rect 2041 5791 2099 5797
rect 2406 5788 2412 5800
rect 2464 5788 2470 5840
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1762 5760 1768 5772
rect 1443 5732 1768 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2498 5760 2504 5772
rect 2459 5732 2504 5760
rect 2498 5720 2504 5732
rect 2556 5760 2562 5772
rect 8386 5760 8392 5772
rect 2556 5732 8392 5760
rect 2556 5720 2562 5732
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 26694 5624 26700 5636
rect 26655 5596 26700 5624
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2038 5352 2044 5364
rect 1999 5324 2044 5352
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26568 5324 27353 5352
rect 26568 5312 26574 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2038 5148 2044 5160
rect 1443 5120 2044 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 26326 5108 26332 5160
rect 26384 5148 26390 5160
rect 26421 5151 26479 5157
rect 26421 5148 26433 5151
rect 26384 5120 26433 5148
rect 26384 5108 26390 5120
rect 26421 5117 26433 5120
rect 26467 5148 26479 5151
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26467 5120 26985 5148
rect 26467 5117 26479 5120
rect 26421 5111 26479 5117
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1762 4808 1768 4820
rect 1719 4780 1768 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5592 2604 6285 2632
rect 5592 2592 5598 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 6273 2595 6331 2601
rect 6288 2428 6316 2595
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 7190 2505 7196 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7184 2496 7196 2505
rect 6779 2468 7196 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7184 2459 7196 2468
rect 7190 2456 7196 2459
rect 7248 2456 7254 2508
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6288 2400 6929 2428
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3516 23400 3568 23452
rect 11980 23400 12032 23452
rect 3516 22516 3568 22568
rect 7932 22516 7984 22568
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 27160 21088 27212 21140
rect 29000 21020 29052 21072
rect 23848 20952 23900 21004
rect 4068 20748 4120 20800
rect 5724 20748 5776 20800
rect 19984 20748 20036 20800
rect 21456 20748 21508 20800
rect 25136 20748 25188 20800
rect 25688 20791 25740 20800
rect 25688 20757 25697 20791
rect 25697 20757 25731 20791
rect 25731 20757 25740 20791
rect 25688 20748 25740 20757
rect 26608 20748 26660 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 940 20544 992 20596
rect 8208 20544 8260 20596
rect 10232 20544 10284 20596
rect 14004 20544 14056 20596
rect 15844 20544 15896 20596
rect 17776 20544 17828 20596
rect 19616 20544 19668 20596
rect 21548 20544 21600 20596
rect 25228 20544 25280 20596
rect 19984 20451 20036 20460
rect 19984 20417 19993 20451
rect 19993 20417 20027 20451
rect 20027 20417 20036 20451
rect 19984 20408 20036 20417
rect 25780 20408 25832 20460
rect 7104 20340 7156 20392
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 14832 20340 14884 20392
rect 17592 20340 17644 20392
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 18604 20204 18656 20256
rect 20720 20340 20772 20392
rect 19432 20272 19484 20324
rect 25688 20272 25740 20324
rect 19340 20247 19392 20256
rect 19340 20213 19349 20247
rect 19349 20213 19383 20247
rect 19383 20213 19392 20247
rect 19340 20204 19392 20213
rect 23848 20204 23900 20256
rect 24032 20247 24084 20256
rect 24032 20213 24041 20247
rect 24041 20213 24075 20247
rect 24075 20213 24084 20247
rect 24032 20204 24084 20213
rect 25228 20204 25280 20256
rect 25596 20247 25648 20256
rect 25596 20213 25605 20247
rect 25605 20213 25639 20247
rect 25639 20213 25648 20247
rect 25596 20204 25648 20213
rect 25872 20204 25924 20256
rect 26148 20204 26200 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 12256 20000 12308 20052
rect 17500 20000 17552 20052
rect 25596 19932 25648 19984
rect 11888 19864 11940 19916
rect 15660 19907 15712 19916
rect 15660 19873 15669 19907
rect 15669 19873 15703 19907
rect 15703 19873 15712 19907
rect 15660 19864 15712 19873
rect 15752 19907 15804 19916
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 17960 19864 18012 19916
rect 18696 19864 18748 19916
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 19432 19839 19484 19848
rect 18328 19728 18380 19780
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 25136 19728 25188 19780
rect 1952 19660 2004 19712
rect 5080 19660 5132 19712
rect 10968 19660 11020 19712
rect 12348 19660 12400 19712
rect 12808 19660 12860 19712
rect 15108 19660 15160 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 16396 19703 16448 19712
rect 16396 19669 16405 19703
rect 16405 19669 16439 19703
rect 16439 19669 16448 19703
rect 16396 19660 16448 19669
rect 24952 19660 25004 19712
rect 25780 19796 25832 19848
rect 26516 19839 26568 19848
rect 26516 19805 26525 19839
rect 26525 19805 26559 19839
rect 26559 19805 26568 19839
rect 26516 19796 26568 19805
rect 25872 19703 25924 19712
rect 25872 19669 25881 19703
rect 25881 19669 25915 19703
rect 25915 19669 25924 19703
rect 25872 19660 25924 19669
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 23388 19456 23440 19508
rect 24032 19456 24084 19508
rect 25872 19456 25924 19508
rect 15752 19388 15804 19440
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 11336 19363 11388 19372
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 9036 19295 9088 19304
rect 2780 19252 2832 19261
rect 9036 19261 9045 19295
rect 9045 19261 9079 19295
rect 9079 19261 9088 19295
rect 9036 19252 9088 19261
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 11704 19320 11756 19372
rect 12624 19320 12676 19372
rect 16488 19320 16540 19372
rect 11060 19252 11112 19304
rect 12532 19252 12584 19304
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 15292 19252 15344 19304
rect 15476 19252 15528 19304
rect 17408 19320 17460 19372
rect 25780 19388 25832 19440
rect 25136 19363 25188 19372
rect 17684 19252 17736 19304
rect 21824 19252 21876 19304
rect 24216 19295 24268 19304
rect 24216 19261 24225 19295
rect 24225 19261 24259 19295
rect 24259 19261 24268 19295
rect 25136 19329 25145 19363
rect 25145 19329 25179 19363
rect 25179 19329 25188 19363
rect 25136 19320 25188 19329
rect 25320 19363 25372 19372
rect 25320 19329 25329 19363
rect 25329 19329 25363 19363
rect 25363 19329 25372 19363
rect 25320 19320 25372 19329
rect 27344 19320 27396 19372
rect 24216 19252 24268 19261
rect 25596 19252 25648 19304
rect 26516 19252 26568 19304
rect 4896 19184 4948 19236
rect 16856 19227 16908 19236
rect 2136 19116 2188 19168
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 3148 19159 3200 19168
rect 3148 19125 3157 19159
rect 3157 19125 3191 19159
rect 3191 19125 3200 19159
rect 3148 19116 3200 19125
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 5080 19116 5132 19168
rect 8116 19159 8168 19168
rect 8116 19125 8125 19159
rect 8125 19125 8159 19159
rect 8159 19125 8168 19159
rect 8116 19116 8168 19125
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11888 19116 11940 19168
rect 16856 19193 16865 19227
rect 16865 19193 16899 19227
rect 16899 19193 16908 19227
rect 16856 19184 16908 19193
rect 19984 19184 20036 19236
rect 13360 19116 13412 19168
rect 15108 19116 15160 19168
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 17868 19159 17920 19168
rect 17868 19125 17877 19159
rect 17877 19125 17911 19159
rect 17911 19125 17920 19159
rect 17868 19116 17920 19125
rect 18328 19159 18380 19168
rect 18328 19125 18337 19159
rect 18337 19125 18371 19159
rect 18371 19125 18380 19159
rect 18328 19116 18380 19125
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 20444 19116 20496 19168
rect 24492 19159 24544 19168
rect 24492 19125 24501 19159
rect 24501 19125 24535 19159
rect 24535 19125 24544 19159
rect 24492 19116 24544 19125
rect 25596 19116 25648 19168
rect 27344 19159 27396 19168
rect 27344 19125 27353 19159
rect 27353 19125 27387 19159
rect 27387 19125 27396 19159
rect 27344 19116 27396 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 3148 18912 3200 18964
rect 4804 18912 4856 18964
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 9036 18912 9088 18964
rect 10232 18955 10284 18964
rect 10232 18921 10241 18955
rect 10241 18921 10275 18955
rect 10275 18921 10284 18955
rect 10232 18912 10284 18921
rect 10876 18912 10928 18964
rect 15752 18912 15804 18964
rect 18328 18912 18380 18964
rect 22560 18955 22612 18964
rect 22560 18921 22569 18955
rect 22569 18921 22603 18955
rect 22603 18921 22612 18955
rect 22560 18912 22612 18921
rect 24492 18912 24544 18964
rect 25320 18955 25372 18964
rect 25320 18921 25329 18955
rect 25329 18921 25363 18955
rect 25363 18921 25372 18955
rect 25320 18912 25372 18921
rect 26332 18912 26384 18964
rect 26976 18955 27028 18964
rect 26976 18921 26985 18955
rect 26985 18921 27019 18955
rect 27019 18921 27028 18955
rect 26976 18912 27028 18921
rect 1952 18887 2004 18896
rect 1952 18853 1961 18887
rect 1961 18853 1995 18887
rect 1995 18853 2004 18887
rect 1952 18844 2004 18853
rect 2688 18844 2740 18896
rect 13084 18844 13136 18896
rect 24216 18887 24268 18896
rect 24216 18853 24250 18887
rect 24250 18853 24268 18887
rect 24216 18844 24268 18853
rect 27068 18844 27120 18896
rect 4712 18776 4764 18828
rect 8116 18776 8168 18828
rect 9588 18776 9640 18828
rect 9680 18776 9732 18828
rect 10784 18776 10836 18828
rect 11336 18776 11388 18828
rect 16304 18776 16356 18828
rect 18144 18819 18196 18828
rect 18144 18785 18178 18819
rect 18178 18785 18196 18819
rect 18144 18776 18196 18785
rect 21640 18776 21692 18828
rect 23388 18776 23440 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 5448 18751 5500 18760
rect 2136 18708 2188 18717
rect 5448 18717 5457 18751
rect 5457 18717 5491 18751
rect 5491 18717 5500 18751
rect 5448 18708 5500 18717
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 1584 18572 1636 18624
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 3700 18615 3752 18624
rect 3700 18581 3709 18615
rect 3709 18581 3743 18615
rect 3743 18581 3752 18615
rect 3700 18572 3752 18581
rect 4896 18615 4948 18624
rect 4896 18581 4905 18615
rect 4905 18581 4939 18615
rect 4939 18581 4948 18615
rect 4896 18572 4948 18581
rect 5264 18572 5316 18624
rect 6920 18572 6972 18624
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 10876 18751 10928 18760
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 16672 18640 16724 18692
rect 17500 18708 17552 18760
rect 17684 18708 17736 18760
rect 20720 18708 20772 18760
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 23940 18751 23992 18760
rect 23940 18717 23949 18751
rect 23949 18717 23983 18751
rect 23983 18717 23992 18751
rect 23940 18708 23992 18717
rect 26332 18708 26384 18760
rect 27344 18708 27396 18760
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 15752 18572 15804 18624
rect 16396 18572 16448 18624
rect 19892 18615 19944 18624
rect 19892 18581 19901 18615
rect 19901 18581 19935 18615
rect 19935 18581 19944 18615
rect 19892 18572 19944 18581
rect 19984 18572 20036 18624
rect 22100 18615 22152 18624
rect 22100 18581 22109 18615
rect 22109 18581 22143 18615
rect 22143 18581 22152 18615
rect 22100 18572 22152 18581
rect 24676 18572 24728 18624
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 2780 18368 2832 18420
rect 4988 18411 5040 18420
rect 4988 18377 4997 18411
rect 4997 18377 5031 18411
rect 5031 18377 5040 18411
rect 4988 18368 5040 18377
rect 5448 18368 5500 18420
rect 5632 18368 5684 18420
rect 6460 18368 6512 18420
rect 6552 18368 6604 18420
rect 10876 18368 10928 18420
rect 11336 18368 11388 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 3700 18300 3752 18352
rect 11520 18300 11572 18352
rect 11796 18343 11848 18352
rect 11796 18309 11805 18343
rect 11805 18309 11839 18343
rect 11839 18309 11848 18343
rect 11796 18300 11848 18309
rect 12440 18411 12492 18420
rect 12440 18377 12449 18411
rect 12449 18377 12483 18411
rect 12483 18377 12492 18411
rect 16580 18411 16632 18420
rect 12440 18368 12492 18377
rect 16580 18377 16589 18411
rect 16589 18377 16623 18411
rect 16623 18377 16632 18411
rect 16580 18368 16632 18377
rect 17500 18411 17552 18420
rect 17500 18377 17509 18411
rect 17509 18377 17543 18411
rect 17543 18377 17552 18411
rect 17500 18368 17552 18377
rect 17776 18368 17828 18420
rect 17868 18368 17920 18420
rect 19892 18368 19944 18420
rect 22560 18368 22612 18420
rect 25872 18368 25924 18420
rect 12900 18300 12952 18352
rect 20168 18343 20220 18352
rect 5632 18275 5684 18284
rect 1584 18096 1636 18148
rect 1676 18028 1728 18080
rect 2964 18164 3016 18216
rect 3148 18164 3200 18216
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 4712 18164 4764 18216
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 2596 18071 2648 18080
rect 2596 18037 2605 18071
rect 2605 18037 2639 18071
rect 2639 18037 2648 18071
rect 2596 18028 2648 18037
rect 2872 18071 2924 18080
rect 2872 18037 2881 18071
rect 2881 18037 2915 18071
rect 2915 18037 2924 18071
rect 2872 18028 2924 18037
rect 4160 18071 4212 18080
rect 4160 18037 4169 18071
rect 4169 18037 4203 18071
rect 4203 18037 4212 18071
rect 4160 18028 4212 18037
rect 4804 18071 4856 18080
rect 4804 18037 4813 18071
rect 4813 18037 4847 18071
rect 4847 18037 4856 18071
rect 4804 18028 4856 18037
rect 7288 18028 7340 18080
rect 8116 18164 8168 18216
rect 12808 18232 12860 18284
rect 20168 18309 20177 18343
rect 20177 18309 20211 18343
rect 20211 18309 20220 18343
rect 20168 18300 20220 18309
rect 21732 18300 21784 18352
rect 26976 18300 27028 18352
rect 18144 18232 18196 18284
rect 19432 18275 19484 18284
rect 19432 18241 19441 18275
rect 19441 18241 19475 18275
rect 19475 18241 19484 18275
rect 19432 18232 19484 18241
rect 19984 18232 20036 18284
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 22652 18275 22704 18284
rect 22652 18241 22661 18275
rect 22661 18241 22695 18275
rect 22695 18241 22704 18275
rect 22652 18232 22704 18241
rect 24676 18275 24728 18284
rect 24676 18241 24685 18275
rect 24685 18241 24719 18275
rect 24719 18241 24728 18275
rect 24676 18232 24728 18241
rect 9312 18164 9364 18216
rect 14924 18164 14976 18216
rect 19892 18164 19944 18216
rect 20720 18207 20772 18216
rect 20720 18173 20729 18207
rect 20729 18173 20763 18207
rect 20763 18173 20772 18207
rect 20720 18164 20772 18173
rect 21640 18164 21692 18216
rect 27068 18164 27120 18216
rect 8576 18096 8628 18148
rect 8116 18028 8168 18080
rect 12348 18096 12400 18148
rect 15752 18096 15804 18148
rect 19340 18096 19392 18148
rect 20168 18096 20220 18148
rect 21364 18096 21416 18148
rect 21916 18096 21968 18148
rect 23940 18096 23992 18148
rect 24216 18096 24268 18148
rect 26240 18096 26292 18148
rect 10140 18028 10192 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 13636 18028 13688 18080
rect 16672 18028 16724 18080
rect 17684 18028 17736 18080
rect 23388 18071 23440 18080
rect 23388 18037 23397 18071
rect 23397 18037 23431 18071
rect 23431 18037 23440 18071
rect 23388 18028 23440 18037
rect 23480 18028 23532 18080
rect 24400 18028 24452 18080
rect 25320 18028 25372 18080
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 4344 17824 4396 17876
rect 4988 17867 5040 17876
rect 4988 17833 4997 17867
rect 4997 17833 5031 17867
rect 5031 17833 5040 17867
rect 4988 17824 5040 17833
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 9680 17824 9732 17876
rect 11704 17824 11756 17876
rect 12900 17867 12952 17876
rect 2596 17756 2648 17808
rect 3516 17756 3568 17808
rect 5632 17756 5684 17808
rect 2044 17688 2096 17740
rect 2964 17688 3016 17740
rect 5172 17688 5224 17740
rect 7932 17688 7984 17740
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 10324 17688 10376 17740
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 12900 17833 12909 17867
rect 12909 17833 12943 17867
rect 12943 17833 12952 17867
rect 12900 17824 12952 17833
rect 15016 17824 15068 17876
rect 15476 17824 15528 17876
rect 17960 17824 18012 17876
rect 18512 17824 18564 17876
rect 18696 17824 18748 17876
rect 20628 17824 20680 17876
rect 21916 17824 21968 17876
rect 22284 17824 22336 17876
rect 22468 17824 22520 17876
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 16580 17756 16632 17808
rect 19432 17756 19484 17808
rect 13452 17688 13504 17740
rect 14924 17688 14976 17740
rect 16672 17731 16724 17740
rect 16672 17697 16681 17731
rect 16681 17697 16715 17731
rect 16715 17697 16724 17731
rect 16672 17688 16724 17697
rect 17684 17688 17736 17740
rect 18972 17688 19024 17740
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4068 17620 4120 17629
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 16488 17620 16540 17672
rect 22652 17756 22704 17808
rect 27252 17756 27304 17808
rect 21364 17688 21416 17740
rect 23020 17688 23072 17740
rect 10876 17552 10928 17604
rect 20444 17620 20496 17672
rect 22192 17663 22244 17672
rect 22192 17629 22201 17663
rect 22201 17629 22235 17663
rect 22235 17629 22244 17663
rect 22192 17620 22244 17629
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 27436 17688 27488 17740
rect 19800 17552 19852 17604
rect 24768 17552 24820 17604
rect 26884 17552 26936 17604
rect 27712 17620 27764 17672
rect 27804 17552 27856 17604
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 9312 17484 9364 17536
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 13268 17484 13320 17536
rect 16304 17527 16356 17536
rect 16304 17493 16313 17527
rect 16313 17493 16347 17527
rect 16347 17493 16356 17527
rect 16304 17484 16356 17493
rect 18972 17527 19024 17536
rect 18972 17493 18981 17527
rect 18981 17493 19015 17527
rect 19015 17493 19024 17527
rect 18972 17484 19024 17493
rect 23572 17527 23624 17536
rect 23572 17493 23581 17527
rect 23581 17493 23615 17527
rect 23615 17493 23624 17527
rect 23572 17484 23624 17493
rect 23756 17484 23808 17536
rect 24400 17484 24452 17536
rect 25228 17484 25280 17536
rect 26516 17527 26568 17536
rect 26516 17493 26525 17527
rect 26525 17493 26559 17527
rect 26559 17493 26568 17527
rect 26516 17484 26568 17493
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 5632 17280 5684 17332
rect 7472 17280 7524 17332
rect 8392 17280 8444 17332
rect 9312 17280 9364 17332
rect 9680 17280 9732 17332
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 11980 17280 12032 17332
rect 12532 17280 12584 17332
rect 16580 17280 16632 17332
rect 21364 17323 21416 17332
rect 21364 17289 21373 17323
rect 21373 17289 21407 17323
rect 21407 17289 21416 17323
rect 21364 17280 21416 17289
rect 21824 17323 21876 17332
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 22192 17280 22244 17332
rect 23388 17280 23440 17332
rect 25780 17280 25832 17332
rect 26424 17323 26476 17332
rect 10324 17212 10376 17264
rect 16672 17212 16724 17264
rect 1492 17076 1544 17128
rect 4344 17119 4396 17128
rect 4344 17085 4378 17119
rect 4378 17085 4396 17119
rect 2228 17008 2280 17060
rect 3148 17008 3200 17060
rect 4344 17076 4396 17085
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 10692 17144 10744 17196
rect 13452 17144 13504 17196
rect 23572 17144 23624 17196
rect 5172 17008 5224 17060
rect 10048 17076 10100 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 12808 17076 12860 17128
rect 14924 17076 14976 17128
rect 17684 17076 17736 17128
rect 21824 17076 21876 17128
rect 26424 17289 26433 17323
rect 26433 17289 26467 17323
rect 26467 17289 26476 17323
rect 26424 17280 26476 17289
rect 26332 17212 26384 17264
rect 26884 17187 26936 17196
rect 26884 17153 26893 17187
rect 26893 17153 26927 17187
rect 26927 17153 26936 17187
rect 26884 17144 26936 17153
rect 27528 17144 27580 17196
rect 26792 17119 26844 17128
rect 8116 17008 8168 17060
rect 8668 17008 8720 17060
rect 10416 17008 10468 17060
rect 12624 17008 12676 17060
rect 15016 17008 15068 17060
rect 18512 17008 18564 17060
rect 21640 17008 21692 17060
rect 23388 17008 23440 17060
rect 26792 17085 26801 17119
rect 26801 17085 26835 17119
rect 26835 17085 26844 17119
rect 26792 17076 26844 17085
rect 24032 17008 24084 17060
rect 6920 16940 6972 16992
rect 11980 16940 12032 16992
rect 13176 16940 13228 16992
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 15752 16940 15804 16992
rect 19892 16940 19944 16992
rect 21548 16940 21600 16992
rect 22192 16940 22244 16992
rect 25504 17008 25556 17060
rect 26424 17008 26476 17060
rect 26332 16983 26384 16992
rect 26332 16949 26341 16983
rect 26341 16949 26375 16983
rect 26375 16949 26384 16983
rect 26332 16940 26384 16949
rect 27252 16940 27304 16992
rect 27436 16983 27488 16992
rect 27436 16949 27445 16983
rect 27445 16949 27479 16983
rect 27479 16949 27488 16983
rect 27436 16940 27488 16949
rect 27712 16940 27764 16992
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 2688 16736 2740 16788
rect 3148 16779 3200 16788
rect 3148 16745 3157 16779
rect 3157 16745 3191 16779
rect 3191 16745 3200 16779
rect 3148 16736 3200 16745
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 4068 16736 4120 16788
rect 4528 16736 4580 16788
rect 5632 16779 5684 16788
rect 5632 16745 5641 16779
rect 5641 16745 5675 16779
rect 5675 16745 5684 16779
rect 5632 16736 5684 16745
rect 6736 16736 6788 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 4620 16668 4672 16720
rect 5908 16711 5960 16720
rect 2596 16600 2648 16652
rect 2964 16600 3016 16652
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 3516 16532 3568 16584
rect 4436 16532 4488 16584
rect 5908 16677 5917 16711
rect 5917 16677 5951 16711
rect 5951 16677 5960 16711
rect 5908 16668 5960 16677
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 8576 16600 8628 16652
rect 7288 16532 7340 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 8668 16575 8720 16584
rect 8668 16541 8677 16575
rect 8677 16541 8711 16575
rect 8711 16541 8720 16575
rect 10232 16736 10284 16788
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 11520 16736 11572 16788
rect 12808 16736 12860 16788
rect 13820 16736 13872 16788
rect 17316 16779 17368 16788
rect 17316 16745 17325 16779
rect 17325 16745 17359 16779
rect 17359 16745 17368 16779
rect 17316 16736 17368 16745
rect 18972 16736 19024 16788
rect 19432 16736 19484 16788
rect 19800 16736 19852 16788
rect 22008 16736 22060 16788
rect 23020 16779 23072 16788
rect 23020 16745 23029 16779
rect 23029 16745 23063 16779
rect 23063 16745 23072 16779
rect 23020 16736 23072 16745
rect 24032 16779 24084 16788
rect 24032 16745 24041 16779
rect 24041 16745 24075 16779
rect 24075 16745 24084 16779
rect 24032 16736 24084 16745
rect 25504 16736 25556 16788
rect 26884 16736 26936 16788
rect 10140 16668 10192 16720
rect 10968 16668 11020 16720
rect 12164 16668 12216 16720
rect 13268 16668 13320 16720
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 13636 16600 13688 16652
rect 16488 16668 16540 16720
rect 17224 16711 17276 16720
rect 17224 16677 17233 16711
rect 17233 16677 17267 16711
rect 17267 16677 17276 16711
rect 17224 16668 17276 16677
rect 18420 16668 18472 16720
rect 21732 16668 21784 16720
rect 22100 16668 22152 16720
rect 24860 16668 24912 16720
rect 25872 16668 25924 16720
rect 10600 16575 10652 16584
rect 8668 16532 8720 16541
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 13820 16532 13872 16584
rect 7564 16507 7616 16516
rect 7564 16473 7573 16507
rect 7573 16473 7607 16507
rect 7607 16473 7616 16507
rect 15384 16600 15436 16652
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16856 16600 16908 16652
rect 18236 16600 18288 16652
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 21272 16600 21324 16652
rect 22652 16600 22704 16652
rect 24768 16643 24820 16652
rect 24768 16609 24777 16643
rect 24777 16609 24811 16643
rect 24811 16609 24820 16643
rect 24768 16600 24820 16609
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 17684 16532 17736 16584
rect 7564 16464 7616 16473
rect 18972 16464 19024 16516
rect 19892 16532 19944 16584
rect 21548 16532 21600 16584
rect 5632 16396 5684 16448
rect 8116 16396 8168 16448
rect 8392 16396 8444 16448
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 12348 16396 12400 16448
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 24952 16600 25004 16652
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 26884 16643 26936 16652
rect 25320 16532 25372 16584
rect 25596 16532 25648 16584
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 26424 16532 26476 16584
rect 27160 16575 27212 16584
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 21916 16396 21968 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 3056 16235 3108 16244
rect 3056 16201 3065 16235
rect 3065 16201 3099 16235
rect 3099 16201 3108 16235
rect 3056 16192 3108 16201
rect 3424 16192 3476 16244
rect 4528 16235 4580 16244
rect 4528 16201 4537 16235
rect 4537 16201 4571 16235
rect 4571 16201 4580 16235
rect 4528 16192 4580 16201
rect 4436 16124 4488 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 3516 16056 3568 16108
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 6460 16192 6512 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 10232 16192 10284 16244
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 15016 16192 15068 16244
rect 15568 16192 15620 16244
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 14740 16124 14792 16133
rect 7564 16099 7616 16108
rect 5816 16056 5868 16065
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 6552 15988 6604 16040
rect 8392 15988 8444 16040
rect 13084 16031 13136 16040
rect 13084 15997 13118 16031
rect 13118 15997 13136 16031
rect 13084 15988 13136 15997
rect 15476 15988 15528 16040
rect 16488 16192 16540 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 18236 16235 18288 16244
rect 18236 16201 18245 16235
rect 18245 16201 18279 16235
rect 18279 16201 18288 16235
rect 18236 16192 18288 16201
rect 21272 16235 21324 16244
rect 21272 16201 21281 16235
rect 21281 16201 21315 16235
rect 21315 16201 21324 16235
rect 21272 16192 21324 16201
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 17316 16124 17368 16176
rect 17684 16056 17736 16108
rect 18236 16056 18288 16108
rect 21364 16056 21416 16108
rect 24032 16192 24084 16244
rect 24676 16192 24728 16244
rect 25780 16192 25832 16244
rect 27160 16192 27212 16244
rect 27528 16167 27580 16176
rect 27528 16133 27537 16167
rect 27537 16133 27571 16167
rect 27571 16133 27580 16167
rect 27528 16124 27580 16133
rect 26148 16099 26200 16108
rect 22100 15988 22152 16040
rect 22376 15988 22428 16040
rect 26148 16065 26157 16099
rect 26157 16065 26191 16099
rect 26191 16065 26200 16099
rect 26148 16056 26200 16065
rect 26424 16031 26476 16040
rect 26424 15997 26458 16031
rect 26458 15997 26476 16031
rect 26424 15988 26476 15997
rect 1952 15963 2004 15972
rect 1952 15929 1961 15963
rect 1961 15929 1995 15963
rect 1995 15929 2004 15963
rect 1952 15920 2004 15929
rect 3056 15920 3108 15972
rect 3424 15920 3476 15972
rect 4988 15920 5040 15972
rect 8300 15920 8352 15972
rect 9036 15920 9088 15972
rect 11612 15920 11664 15972
rect 13636 15920 13688 15972
rect 17040 15920 17092 15972
rect 18328 15920 18380 15972
rect 19064 15920 19116 15972
rect 24492 15920 24544 15972
rect 25412 15920 25464 15972
rect 25872 15920 25924 15972
rect 3240 15852 3292 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 6920 15895 6972 15904
rect 5632 15852 5684 15861
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 7288 15852 7340 15904
rect 8576 15852 8628 15904
rect 10140 15852 10192 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 15660 15852 15712 15904
rect 19340 15852 19392 15904
rect 21916 15852 21968 15904
rect 22192 15852 22244 15904
rect 25596 15895 25648 15904
rect 25596 15861 25605 15895
rect 25605 15861 25639 15895
rect 25639 15861 25648 15895
rect 25596 15852 25648 15861
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 1952 15648 2004 15700
rect 4620 15691 4672 15700
rect 4620 15657 4629 15691
rect 4629 15657 4663 15691
rect 4663 15657 4672 15691
rect 4620 15648 4672 15657
rect 5356 15648 5408 15700
rect 7564 15648 7616 15700
rect 8484 15648 8536 15700
rect 10784 15648 10836 15700
rect 12348 15648 12400 15700
rect 13728 15691 13780 15700
rect 13728 15657 13737 15691
rect 13737 15657 13771 15691
rect 13771 15657 13780 15691
rect 13728 15648 13780 15657
rect 13820 15648 13872 15700
rect 2596 15580 2648 15632
rect 7288 15580 7340 15632
rect 8576 15580 8628 15632
rect 10692 15580 10744 15632
rect 1952 15512 2004 15564
rect 4068 15512 4120 15564
rect 4988 15512 5040 15564
rect 5448 15512 5500 15564
rect 7656 15512 7708 15564
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 2872 15444 2924 15496
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 2044 15376 2096 15428
rect 8300 15376 8352 15428
rect 10600 15444 10652 15496
rect 12348 15512 12400 15564
rect 11244 15444 11296 15496
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 9588 15376 9640 15428
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 8392 15308 8444 15360
rect 9496 15308 9548 15360
rect 13452 15376 13504 15428
rect 15844 15648 15896 15700
rect 16304 15648 16356 15700
rect 17408 15648 17460 15700
rect 18420 15691 18472 15700
rect 18420 15657 18429 15691
rect 18429 15657 18463 15691
rect 18463 15657 18472 15691
rect 18420 15648 18472 15657
rect 21364 15648 21416 15700
rect 22376 15648 22428 15700
rect 22652 15648 22704 15700
rect 23388 15648 23440 15700
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 26148 15691 26200 15700
rect 26148 15657 26157 15691
rect 26157 15657 26191 15691
rect 26191 15657 26200 15691
rect 26148 15648 26200 15657
rect 26516 15648 26568 15700
rect 27620 15648 27672 15700
rect 15568 15623 15620 15632
rect 15568 15589 15602 15623
rect 15602 15589 15620 15623
rect 15568 15580 15620 15589
rect 17960 15580 18012 15632
rect 25320 15580 25372 15632
rect 25596 15580 25648 15632
rect 18788 15555 18840 15564
rect 18788 15521 18797 15555
rect 18797 15521 18831 15555
rect 18831 15521 18840 15555
rect 18788 15512 18840 15521
rect 22192 15555 22244 15564
rect 22192 15521 22226 15555
rect 22226 15521 22244 15555
rect 22192 15512 22244 15521
rect 25136 15512 25188 15564
rect 18972 15487 19024 15496
rect 11520 15308 11572 15360
rect 14648 15308 14700 15360
rect 18972 15453 18981 15487
rect 18981 15453 19015 15487
rect 19015 15453 19024 15487
rect 18972 15444 19024 15453
rect 21916 15487 21968 15496
rect 21916 15453 21925 15487
rect 21925 15453 21959 15487
rect 21959 15453 21968 15487
rect 21916 15444 21968 15453
rect 25044 15444 25096 15496
rect 25688 15512 25740 15564
rect 26424 15512 26476 15564
rect 26332 15444 26384 15496
rect 27528 15444 27580 15496
rect 24032 15376 24084 15428
rect 25780 15376 25832 15428
rect 26424 15376 26476 15428
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 24124 15308 24176 15360
rect 26516 15351 26568 15360
rect 26516 15317 26525 15351
rect 26525 15317 26559 15351
rect 26559 15317 26568 15351
rect 26516 15308 26568 15317
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 3516 15104 3568 15156
rect 6828 15104 6880 15156
rect 8300 15104 8352 15156
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 9956 15104 10008 15156
rect 15752 15104 15804 15156
rect 10600 15036 10652 15088
rect 1860 14900 1912 14952
rect 2320 14900 2372 14952
rect 1952 14764 2004 14816
rect 4068 14900 4120 14952
rect 6920 14900 6972 14952
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 4712 14832 4764 14884
rect 7932 14832 7984 14884
rect 11520 14968 11572 15020
rect 12716 14968 12768 15020
rect 15660 15036 15712 15088
rect 16304 15036 16356 15088
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 11796 14900 11848 14952
rect 12624 14900 12676 14952
rect 11244 14875 11296 14884
rect 11244 14841 11253 14875
rect 11253 14841 11287 14875
rect 11287 14841 11296 14875
rect 11244 14832 11296 14841
rect 4988 14764 5040 14816
rect 5448 14764 5500 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7748 14764 7800 14816
rect 8392 14764 8444 14816
rect 10784 14764 10836 14816
rect 11888 14764 11940 14816
rect 12992 14832 13044 14884
rect 16580 15104 16632 15156
rect 17868 15104 17920 15156
rect 18972 15104 19024 15156
rect 21640 15104 21692 15156
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 25688 15147 25740 15156
rect 23388 15104 23440 15113
rect 18236 15036 18288 15088
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 21548 15036 21600 15088
rect 21916 15036 21968 15088
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 25688 15113 25697 15147
rect 25697 15113 25731 15147
rect 25731 15113 25740 15147
rect 25688 15104 25740 15113
rect 27528 15104 27580 15156
rect 25596 15036 25648 15088
rect 21456 14900 21508 14952
rect 21824 14900 21876 14952
rect 26424 14943 26476 14952
rect 26424 14909 26458 14943
rect 26458 14909 26476 14943
rect 26424 14900 26476 14909
rect 19340 14875 19392 14884
rect 19340 14841 19374 14875
rect 19374 14841 19392 14875
rect 19340 14832 19392 14841
rect 20352 14832 20404 14884
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 13268 14764 13320 14816
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 15016 14764 15068 14816
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 15752 14764 15804 14816
rect 16764 14807 16816 14816
rect 16764 14773 16773 14807
rect 16773 14773 16807 14807
rect 16807 14773 16816 14807
rect 16764 14764 16816 14773
rect 18236 14764 18288 14816
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 21916 14832 21968 14884
rect 24032 14875 24084 14884
rect 24032 14841 24041 14875
rect 24041 14841 24075 14875
rect 24075 14841 24084 14875
rect 24032 14832 24084 14841
rect 22192 14764 22244 14816
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 25044 14764 25096 14816
rect 25136 14764 25188 14816
rect 27344 14764 27396 14816
rect 27712 14764 27764 14816
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 2872 14603 2924 14612
rect 2872 14569 2881 14603
rect 2881 14569 2915 14603
rect 2915 14569 2924 14603
rect 2872 14560 2924 14569
rect 4712 14603 4764 14612
rect 4712 14569 4721 14603
rect 4721 14569 4755 14603
rect 4755 14569 4764 14603
rect 4712 14560 4764 14569
rect 5816 14560 5868 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 9496 14560 9548 14612
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 12348 14560 12400 14612
rect 15200 14560 15252 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 16948 14560 17000 14612
rect 18788 14560 18840 14612
rect 19708 14603 19760 14612
rect 19708 14569 19717 14603
rect 19717 14569 19751 14603
rect 19751 14569 19760 14603
rect 19708 14560 19760 14569
rect 20352 14603 20404 14612
rect 20352 14569 20361 14603
rect 20361 14569 20395 14603
rect 20395 14569 20404 14603
rect 20352 14560 20404 14569
rect 21272 14560 21324 14612
rect 23480 14560 23532 14612
rect 24952 14560 25004 14612
rect 25228 14560 25280 14612
rect 26424 14560 26476 14612
rect 26516 14560 26568 14612
rect 28264 14560 28316 14612
rect 1860 14492 1912 14544
rect 5356 14492 5408 14544
rect 7288 14492 7340 14544
rect 10600 14492 10652 14544
rect 16672 14535 16724 14544
rect 16672 14501 16706 14535
rect 16706 14501 16724 14535
rect 16672 14492 16724 14501
rect 24032 14492 24084 14544
rect 25504 14492 25556 14544
rect 27620 14535 27672 14544
rect 27620 14501 27629 14535
rect 27629 14501 27663 14535
rect 27663 14501 27672 14535
rect 27620 14492 27672 14501
rect 2780 14424 2832 14476
rect 4252 14424 4304 14476
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 10416 14467 10468 14476
rect 10416 14433 10450 14467
rect 10450 14433 10468 14467
rect 10416 14424 10468 14433
rect 12716 14424 12768 14476
rect 13268 14424 13320 14476
rect 18972 14424 19024 14476
rect 19432 14424 19484 14476
rect 19524 14424 19576 14476
rect 22100 14424 22152 14476
rect 26516 14424 26568 14476
rect 4988 14356 5040 14408
rect 8668 14399 8720 14408
rect 2872 14220 2924 14272
rect 4068 14220 4120 14272
rect 4988 14220 5040 14272
rect 8668 14365 8677 14399
rect 8677 14365 8711 14399
rect 8711 14365 8720 14399
rect 8668 14356 8720 14365
rect 10140 14399 10192 14408
rect 8300 14288 8352 14340
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 14648 14356 14700 14408
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 21272 14356 21324 14408
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 27160 14399 27212 14408
rect 14004 14331 14056 14340
rect 14004 14297 14013 14331
rect 14013 14297 14047 14331
rect 14047 14297 14056 14331
rect 14004 14288 14056 14297
rect 19340 14288 19392 14340
rect 23204 14288 23256 14340
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 6368 14220 6420 14272
rect 6736 14220 6788 14272
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 19708 14220 19760 14272
rect 22192 14220 22244 14272
rect 26332 14288 26384 14340
rect 26608 14288 26660 14340
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 4252 14016 4304 14068
rect 5356 14016 5408 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7288 14016 7340 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 4344 13948 4396 14000
rect 5540 13948 5592 14000
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 7380 13923 7432 13932
rect 5816 13880 5868 13889
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9312 13880 9364 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 4988 13812 5040 13864
rect 6828 13812 6880 13864
rect 8668 13812 8720 13864
rect 10416 13880 10468 13932
rect 12072 14016 12124 14068
rect 12624 14016 12676 14068
rect 14648 14016 14700 14068
rect 15200 14016 15252 14068
rect 16672 14016 16724 14068
rect 18512 14016 18564 14068
rect 19064 14016 19116 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 21824 14059 21876 14068
rect 21824 14025 21833 14059
rect 21833 14025 21867 14059
rect 21867 14025 21876 14059
rect 21824 14016 21876 14025
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 24216 14016 24268 14068
rect 24400 14016 24452 14068
rect 26700 14059 26752 14068
rect 26700 14025 26709 14059
rect 26709 14025 26743 14059
rect 26743 14025 26752 14059
rect 26700 14016 26752 14025
rect 27160 14016 27212 14068
rect 28264 14059 28316 14068
rect 28264 14025 28273 14059
rect 28273 14025 28307 14059
rect 28307 14025 28316 14059
rect 28264 14016 28316 14025
rect 12716 13880 12768 13932
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 26056 13948 26108 14000
rect 26148 13948 26200 14000
rect 19156 13880 19208 13932
rect 20352 13880 20404 13932
rect 22652 13880 22704 13932
rect 27344 13880 27396 13932
rect 27620 13880 27672 13932
rect 10048 13812 10100 13864
rect 2872 13744 2924 13796
rect 5540 13787 5592 13796
rect 5540 13753 5549 13787
rect 5549 13753 5583 13787
rect 5583 13753 5592 13787
rect 5540 13744 5592 13753
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 7288 13744 7340 13753
rect 12072 13812 12124 13864
rect 14832 13855 14884 13864
rect 11428 13744 11480 13796
rect 14832 13821 14841 13855
rect 14841 13821 14875 13855
rect 14875 13821 14884 13855
rect 14832 13812 14884 13821
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 18972 13812 19024 13864
rect 12808 13787 12860 13796
rect 12808 13753 12817 13787
rect 12817 13753 12851 13787
rect 12851 13753 12860 13787
rect 12808 13744 12860 13753
rect 15568 13744 15620 13796
rect 19064 13787 19116 13796
rect 19064 13753 19073 13787
rect 19073 13753 19107 13787
rect 19107 13753 19116 13787
rect 19064 13744 19116 13753
rect 19524 13812 19576 13864
rect 20076 13812 20128 13864
rect 22100 13812 22152 13864
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 25504 13812 25556 13864
rect 26700 13812 26752 13864
rect 20168 13744 20220 13796
rect 2780 13676 2832 13728
rect 5356 13676 5408 13728
rect 6368 13676 6420 13728
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 10140 13676 10192 13728
rect 10508 13676 10560 13728
rect 11336 13676 11388 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 14004 13719 14056 13728
rect 12900 13676 12952 13685
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 14924 13676 14976 13728
rect 16396 13676 16448 13728
rect 17132 13676 17184 13728
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 23204 13744 23256 13796
rect 23664 13744 23716 13796
rect 24768 13744 24820 13796
rect 27160 13744 27212 13796
rect 22468 13676 22520 13728
rect 26884 13719 26936 13728
rect 26884 13685 26893 13719
rect 26893 13685 26927 13719
rect 26927 13685 26936 13719
rect 26884 13676 26936 13685
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 5172 13472 5224 13524
rect 5816 13472 5868 13524
rect 9312 13515 9364 13524
rect 9312 13481 9321 13515
rect 9321 13481 9355 13515
rect 9355 13481 9364 13515
rect 9312 13472 9364 13481
rect 10416 13472 10468 13524
rect 11336 13472 11388 13524
rect 12256 13472 12308 13524
rect 13176 13472 13228 13524
rect 15200 13472 15252 13524
rect 19892 13472 19944 13524
rect 19984 13472 20036 13524
rect 20168 13472 20220 13524
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 23664 13472 23716 13524
rect 25320 13515 25372 13524
rect 25320 13481 25329 13515
rect 25329 13481 25363 13515
rect 25363 13481 25372 13515
rect 25320 13472 25372 13481
rect 26148 13472 26200 13524
rect 26884 13515 26936 13524
rect 26884 13481 26893 13515
rect 26893 13481 26927 13515
rect 26927 13481 26936 13515
rect 26884 13472 26936 13481
rect 27620 13515 27672 13524
rect 27620 13481 27629 13515
rect 27629 13481 27663 13515
rect 27663 13481 27672 13515
rect 27620 13472 27672 13481
rect 5356 13404 5408 13456
rect 15292 13404 15344 13456
rect 16856 13404 16908 13456
rect 17776 13404 17828 13456
rect 19616 13447 19668 13456
rect 19616 13413 19625 13447
rect 19625 13413 19659 13447
rect 19659 13413 19668 13447
rect 19616 13404 19668 13413
rect 2412 13336 2464 13388
rect 6736 13379 6788 13388
rect 6736 13345 6770 13379
rect 6770 13345 6788 13379
rect 6736 13336 6788 13345
rect 11336 13336 11388 13388
rect 12164 13336 12216 13388
rect 15016 13336 15068 13388
rect 20812 13336 20864 13388
rect 23020 13336 23072 13388
rect 24400 13404 24452 13456
rect 24676 13336 24728 13388
rect 26056 13336 26108 13388
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 2964 13268 3016 13320
rect 5264 13268 5316 13320
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 6368 13268 6420 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 13176 13311 13228 13320
rect 4896 13243 4948 13252
rect 4896 13209 4905 13243
rect 4905 13209 4939 13243
rect 4939 13209 4948 13243
rect 4896 13200 4948 13209
rect 8208 13200 8260 13252
rect 11520 13200 11572 13252
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 20444 13268 20496 13320
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 26976 13311 27028 13320
rect 26976 13277 26985 13311
rect 26985 13277 27019 13311
rect 27019 13277 27028 13311
rect 26976 13268 27028 13277
rect 27528 13268 27580 13320
rect 12900 13200 12952 13252
rect 15384 13200 15436 13252
rect 26516 13243 26568 13252
rect 26516 13209 26525 13243
rect 26525 13209 26559 13243
rect 26559 13209 26568 13243
rect 26516 13200 26568 13209
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 2780 13132 2832 13184
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 7196 13132 7248 13184
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 12808 13132 12860 13184
rect 14556 13132 14608 13184
rect 14924 13132 14976 13184
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 18512 13132 18564 13141
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 20996 13132 21048 13184
rect 22100 13132 22152 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 2596 12928 2648 12980
rect 5080 12928 5132 12980
rect 5264 12928 5316 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 11060 12928 11112 12980
rect 11428 12928 11480 12980
rect 13176 12928 13228 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 14464 12928 14516 12980
rect 15016 12971 15068 12980
rect 2872 12860 2924 12912
rect 5448 12860 5500 12912
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 11520 12792 11572 12844
rect 13360 12792 13412 12844
rect 1768 12724 1820 12776
rect 6828 12724 6880 12776
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8392 12724 8444 12776
rect 2780 12656 2832 12708
rect 2964 12656 3016 12708
rect 3700 12656 3752 12708
rect 6736 12656 6788 12708
rect 8116 12656 8168 12708
rect 9956 12724 10008 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 10508 12656 10560 12708
rect 12256 12699 12308 12708
rect 12256 12665 12265 12699
rect 12265 12665 12299 12699
rect 12299 12665 12308 12699
rect 14280 12724 14332 12776
rect 15016 12937 15025 12971
rect 15025 12937 15059 12971
rect 15059 12937 15068 12971
rect 15016 12928 15068 12937
rect 15844 12928 15896 12980
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 18788 12928 18840 12980
rect 20536 12928 20588 12980
rect 20904 12928 20956 12980
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 23572 12928 23624 12980
rect 24400 12928 24452 12980
rect 21364 12903 21416 12912
rect 21364 12869 21373 12903
rect 21373 12869 21407 12903
rect 21407 12869 21416 12903
rect 21364 12860 21416 12869
rect 24952 12860 25004 12912
rect 15292 12792 15344 12844
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20720 12792 20772 12844
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 16396 12724 16448 12776
rect 22192 12792 22244 12844
rect 26976 12928 27028 12980
rect 27344 12971 27396 12980
rect 27344 12937 27353 12971
rect 27353 12937 27387 12971
rect 27387 12937 27396 12971
rect 27344 12928 27396 12937
rect 27528 12860 27580 12912
rect 22008 12724 22060 12776
rect 23940 12767 23992 12776
rect 23940 12733 23949 12767
rect 23949 12733 23983 12767
rect 23983 12733 23992 12767
rect 23940 12724 23992 12733
rect 24860 12724 24912 12776
rect 25320 12767 25372 12776
rect 25320 12733 25354 12767
rect 25354 12733 25372 12767
rect 25320 12724 25372 12733
rect 27528 12767 27580 12776
rect 27528 12733 27537 12767
rect 27537 12733 27571 12767
rect 27571 12733 27580 12767
rect 27528 12724 27580 12733
rect 12256 12656 12308 12665
rect 13360 12656 13412 12708
rect 13544 12656 13596 12708
rect 2504 12588 2556 12640
rect 4344 12588 4396 12640
rect 5356 12588 5408 12640
rect 6368 12588 6420 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 7748 12631 7800 12640
rect 7748 12597 7757 12631
rect 7757 12597 7791 12631
rect 7791 12597 7800 12631
rect 7748 12588 7800 12597
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 11612 12588 11664 12640
rect 16764 12656 16816 12708
rect 17868 12699 17920 12708
rect 17868 12665 17877 12699
rect 17877 12665 17911 12699
rect 17911 12665 17920 12699
rect 17868 12656 17920 12665
rect 19800 12656 19852 12708
rect 16488 12631 16540 12640
rect 16488 12597 16497 12631
rect 16497 12597 16531 12631
rect 16531 12597 16540 12631
rect 16488 12588 16540 12597
rect 17132 12588 17184 12640
rect 17776 12588 17828 12640
rect 19248 12588 19300 12640
rect 20628 12588 20680 12640
rect 22376 12631 22428 12640
rect 22376 12597 22385 12631
rect 22385 12597 22419 12631
rect 22419 12597 22428 12631
rect 22376 12588 22428 12597
rect 26424 12631 26476 12640
rect 26424 12597 26433 12631
rect 26433 12597 26467 12631
rect 26467 12597 26476 12631
rect 26424 12588 26476 12597
rect 27804 12588 27856 12640
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 2504 12384 2556 12436
rect 6828 12384 6880 12436
rect 7104 12384 7156 12436
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 8208 12384 8260 12436
rect 10048 12384 10100 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 13084 12384 13136 12436
rect 15108 12384 15160 12436
rect 15660 12384 15712 12436
rect 1860 12316 1912 12368
rect 6368 12316 6420 12368
rect 11336 12316 11388 12368
rect 11520 12316 11572 12368
rect 15384 12316 15436 12368
rect 16672 12384 16724 12436
rect 20812 12384 20864 12436
rect 22008 12384 22060 12436
rect 24216 12384 24268 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 25320 12384 25372 12436
rect 27344 12384 27396 12436
rect 16764 12359 16816 12368
rect 16764 12325 16773 12359
rect 16773 12325 16807 12359
rect 16807 12325 16816 12359
rect 16764 12316 16816 12325
rect 17868 12316 17920 12368
rect 18512 12316 18564 12368
rect 1584 12248 1636 12300
rect 5816 12248 5868 12300
rect 7288 12248 7340 12300
rect 8208 12248 8260 12300
rect 10876 12248 10928 12300
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 21272 12316 21324 12368
rect 22192 12316 22244 12368
rect 23940 12316 23992 12368
rect 24584 12316 24636 12368
rect 21180 12291 21232 12300
rect 21180 12257 21214 12291
rect 21214 12257 21232 12291
rect 21180 12248 21232 12257
rect 23480 12248 23532 12300
rect 25412 12316 25464 12368
rect 25136 12248 25188 12300
rect 26516 12248 26568 12300
rect 3056 12223 3108 12232
rect 2228 12112 2280 12164
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 7932 12180 7984 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10508 12180 10560 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17776 12180 17828 12232
rect 20628 12180 20680 12232
rect 25044 12180 25096 12232
rect 25412 12223 25464 12232
rect 25412 12189 25421 12223
rect 25421 12189 25455 12223
rect 25455 12189 25464 12223
rect 25412 12180 25464 12189
rect 25688 12180 25740 12232
rect 27620 12180 27672 12232
rect 28080 12180 28132 12232
rect 2044 12044 2096 12096
rect 3424 12112 3476 12164
rect 3700 12112 3752 12164
rect 2504 12044 2556 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4160 12044 4212 12096
rect 7380 12112 7432 12164
rect 16856 12112 16908 12164
rect 24584 12112 24636 12164
rect 26424 12112 26476 12164
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 15384 12044 15436 12096
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 19156 12044 19208 12096
rect 24676 12044 24728 12096
rect 26976 12044 27028 12096
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 2596 11840 2648 11892
rect 4436 11840 4488 11892
rect 4620 11840 4672 11892
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 7564 11840 7616 11892
rect 7840 11840 7892 11892
rect 9956 11883 10008 11892
rect 9956 11849 9965 11883
rect 9965 11849 9999 11883
rect 9999 11849 10008 11883
rect 9956 11840 10008 11849
rect 10048 11840 10100 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 11520 11840 11572 11892
rect 12532 11840 12584 11892
rect 3240 11772 3292 11824
rect 3700 11772 3752 11824
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 4988 11772 5040 11824
rect 6368 11772 6420 11824
rect 11336 11772 11388 11824
rect 12624 11772 12676 11824
rect 6644 11704 6696 11756
rect 7104 11704 7156 11756
rect 7932 11704 7984 11756
rect 8484 11704 8536 11756
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 16672 11840 16724 11892
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 20720 11840 20772 11892
rect 23480 11883 23532 11892
rect 23480 11849 23489 11883
rect 23489 11849 23523 11883
rect 23523 11849 23532 11883
rect 23480 11840 23532 11849
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 25688 11883 25740 11892
rect 25688 11849 25697 11883
rect 25697 11849 25731 11883
rect 25731 11849 25740 11883
rect 25688 11840 25740 11849
rect 16764 11772 16816 11824
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17408 11704 17460 11756
rect 17776 11704 17828 11756
rect 17960 11772 18012 11824
rect 18328 11772 18380 11824
rect 18420 11704 18472 11756
rect 21272 11772 21324 11824
rect 24860 11772 24912 11824
rect 26516 11840 26568 11892
rect 28080 11883 28132 11892
rect 28080 11849 28089 11883
rect 28089 11849 28123 11883
rect 28123 11849 28132 11883
rect 28080 11840 28132 11849
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 23756 11704 23808 11756
rect 20536 11636 20588 11688
rect 24216 11704 24268 11756
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 24584 11704 24636 11713
rect 26148 11679 26200 11688
rect 26148 11645 26157 11679
rect 26157 11645 26191 11679
rect 26191 11645 26200 11679
rect 26148 11636 26200 11645
rect 4252 11568 4304 11620
rect 6276 11568 6328 11620
rect 8944 11568 8996 11620
rect 14556 11568 14608 11620
rect 16856 11611 16908 11620
rect 16856 11577 16865 11611
rect 16865 11577 16899 11611
rect 16899 11577 16908 11611
rect 16856 11568 16908 11577
rect 17776 11568 17828 11620
rect 19156 11568 19208 11620
rect 20812 11568 20864 11620
rect 22192 11568 22244 11620
rect 25412 11568 25464 11620
rect 1492 11500 1544 11552
rect 4528 11500 4580 11552
rect 4804 11500 4856 11552
rect 5816 11500 5868 11552
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 16488 11500 16540 11552
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 20168 11500 20220 11552
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 24032 11543 24084 11552
rect 24032 11509 24041 11543
rect 24041 11509 24075 11543
rect 24075 11509 24084 11543
rect 24032 11500 24084 11509
rect 27068 11500 27120 11552
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 1400 11296 1452 11348
rect 2412 11339 2464 11348
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 2964 11296 3016 11348
rect 3516 11296 3568 11348
rect 4344 11296 4396 11348
rect 5816 11296 5868 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 10416 11296 10468 11348
rect 14556 11296 14608 11348
rect 15568 11296 15620 11348
rect 16396 11296 16448 11348
rect 4252 11228 4304 11280
rect 6644 11271 6696 11280
rect 6644 11237 6653 11271
rect 6653 11237 6687 11271
rect 6687 11237 6696 11271
rect 6644 11228 6696 11237
rect 7196 11228 7248 11280
rect 8024 11228 8076 11280
rect 8116 11228 8168 11280
rect 9588 11228 9640 11280
rect 10232 11228 10284 11280
rect 15384 11228 15436 11280
rect 16488 11228 16540 11280
rect 16948 11271 17000 11280
rect 16948 11237 16957 11271
rect 16957 11237 16991 11271
rect 16991 11237 17000 11271
rect 16948 11228 17000 11237
rect 17592 11296 17644 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 21456 11339 21508 11348
rect 21456 11305 21465 11339
rect 21465 11305 21499 11339
rect 21499 11305 21508 11339
rect 21456 11296 21508 11305
rect 22008 11296 22060 11348
rect 22192 11339 22244 11348
rect 22192 11305 22201 11339
rect 22201 11305 22235 11339
rect 22235 11305 22244 11339
rect 22192 11296 22244 11305
rect 23020 11296 23072 11348
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 25136 11296 25188 11348
rect 25412 11339 25464 11348
rect 25412 11305 25421 11339
rect 25421 11305 25455 11339
rect 25455 11305 25464 11339
rect 25412 11296 25464 11305
rect 26700 11296 26752 11348
rect 26976 11339 27028 11348
rect 26976 11305 26985 11339
rect 26985 11305 27019 11339
rect 27019 11305 27028 11339
rect 26976 11296 27028 11305
rect 27620 11296 27672 11348
rect 17960 11271 18012 11280
rect 17960 11237 17969 11271
rect 17969 11237 18003 11271
rect 18003 11237 18012 11271
rect 17960 11228 18012 11237
rect 3516 11160 3568 11212
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 3056 11135 3108 11144
rect 2320 11092 2372 11101
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 4804 11160 4856 11212
rect 6368 11092 6420 11144
rect 6736 11092 6788 11144
rect 9772 11092 9824 11144
rect 18512 11203 18564 11212
rect 9680 11067 9732 11076
rect 9680 11033 9689 11067
rect 9689 11033 9723 11067
rect 9723 11033 9732 11067
rect 9680 11024 9732 11033
rect 18512 11169 18521 11203
rect 18521 11169 18555 11203
rect 18555 11169 18564 11203
rect 18512 11160 18564 11169
rect 19248 11160 19300 11212
rect 19800 11228 19852 11280
rect 21364 11160 21416 11212
rect 22652 11228 22704 11280
rect 24032 11228 24084 11280
rect 26148 11271 26200 11280
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 18052 11135 18104 11144
rect 16488 11092 16540 11101
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 20168 11092 20220 11144
rect 22928 11135 22980 11144
rect 22928 11101 22937 11135
rect 22937 11101 22971 11135
rect 22971 11101 22980 11135
rect 22928 11092 22980 11101
rect 23572 11160 23624 11212
rect 26148 11237 26157 11271
rect 26157 11237 26191 11271
rect 26191 11237 26200 11271
rect 26148 11228 26200 11237
rect 16948 11024 17000 11076
rect 19156 11024 19208 11076
rect 23388 11024 23440 11076
rect 24768 11160 24820 11212
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 27068 11135 27120 11144
rect 27068 11101 27077 11135
rect 27077 11101 27111 11135
rect 27111 11101 27120 11135
rect 27068 11092 27120 11101
rect 16856 10956 16908 11008
rect 21180 10999 21232 11008
rect 21180 10965 21189 10999
rect 21189 10965 21223 10999
rect 21223 10965 21232 10999
rect 21180 10956 21232 10965
rect 23112 10956 23164 11008
rect 26332 11024 26384 11076
rect 26608 10956 26660 11008
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 2964 10752 3016 10804
rect 3792 10752 3844 10804
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 4620 10684 4672 10736
rect 4712 10684 4764 10736
rect 2780 10616 2832 10668
rect 3792 10616 3844 10668
rect 3884 10616 3936 10668
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 5448 10616 5500 10668
rect 6644 10752 6696 10804
rect 7380 10752 7432 10804
rect 8760 10752 8812 10804
rect 8300 10684 8352 10736
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 3516 10548 3568 10557
rect 4620 10548 4672 10600
rect 6368 10548 6420 10600
rect 7932 10591 7984 10600
rect 2228 10412 2280 10464
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 4068 10480 4120 10532
rect 4344 10480 4396 10532
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 15568 10752 15620 10804
rect 16488 10752 16540 10804
rect 17868 10752 17920 10804
rect 17960 10752 18012 10804
rect 19248 10752 19300 10804
rect 19340 10752 19392 10804
rect 17408 10684 17460 10736
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 18512 10659 18564 10668
rect 18512 10625 18521 10659
rect 18521 10625 18555 10659
rect 18555 10625 18564 10659
rect 18512 10616 18564 10625
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 20720 10752 20772 10804
rect 22928 10752 22980 10804
rect 23112 10795 23164 10804
rect 23112 10761 23121 10795
rect 23121 10761 23155 10795
rect 23155 10761 23164 10795
rect 23112 10752 23164 10761
rect 24400 10752 24452 10804
rect 26700 10752 26752 10804
rect 27620 10752 27672 10804
rect 21364 10684 21416 10736
rect 25320 10684 25372 10736
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 20720 10616 20772 10668
rect 21180 10616 21232 10668
rect 21456 10616 21508 10668
rect 22008 10616 22060 10668
rect 23572 10616 23624 10668
rect 20260 10548 20312 10600
rect 2504 10412 2556 10421
rect 4436 10412 4488 10464
rect 9312 10480 9364 10532
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6736 10412 6788 10464
rect 8576 10455 8628 10464
rect 8576 10421 8585 10455
rect 8585 10421 8619 10455
rect 8619 10421 8628 10455
rect 8576 10412 8628 10421
rect 9772 10412 9824 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 16856 10412 16908 10464
rect 20536 10480 20588 10532
rect 23480 10480 23532 10532
rect 24584 10480 24636 10532
rect 27068 10616 27120 10668
rect 26608 10591 26660 10600
rect 26608 10557 26617 10591
rect 26617 10557 26651 10591
rect 26651 10557 26660 10591
rect 26608 10548 26660 10557
rect 25964 10523 26016 10532
rect 25964 10489 25973 10523
rect 25973 10489 26007 10523
rect 26007 10489 26016 10523
rect 25964 10480 26016 10489
rect 26424 10480 26476 10532
rect 20720 10455 20772 10464
rect 20720 10421 20729 10455
rect 20729 10421 20763 10455
rect 20763 10421 20772 10455
rect 20720 10412 20772 10421
rect 21548 10455 21600 10464
rect 21548 10421 21557 10455
rect 21557 10421 21591 10455
rect 21591 10421 21600 10455
rect 21548 10412 21600 10421
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 3424 10208 3476 10260
rect 4252 10208 4304 10260
rect 4344 10183 4396 10192
rect 4344 10149 4378 10183
rect 4378 10149 4396 10183
rect 8208 10208 8260 10260
rect 8576 10208 8628 10260
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 18052 10208 18104 10260
rect 18236 10251 18288 10260
rect 18236 10217 18245 10251
rect 18245 10217 18279 10251
rect 18279 10217 18288 10251
rect 18236 10208 18288 10217
rect 18420 10208 18472 10260
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 21548 10251 21600 10260
rect 21548 10217 21557 10251
rect 21557 10217 21591 10251
rect 21591 10217 21600 10251
rect 21548 10208 21600 10217
rect 21732 10208 21784 10260
rect 22652 10251 22704 10260
rect 22652 10217 22661 10251
rect 22661 10217 22695 10251
rect 22695 10217 22704 10251
rect 22652 10208 22704 10217
rect 23020 10251 23072 10260
rect 23020 10217 23029 10251
rect 23029 10217 23063 10251
rect 23063 10217 23072 10251
rect 23020 10208 23072 10217
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 26608 10208 26660 10260
rect 27068 10251 27120 10260
rect 27068 10217 27077 10251
rect 27077 10217 27111 10251
rect 27111 10217 27120 10251
rect 27068 10208 27120 10217
rect 27160 10208 27212 10260
rect 4344 10140 4396 10149
rect 9036 10140 9088 10192
rect 9312 10140 9364 10192
rect 17408 10140 17460 10192
rect 18328 10183 18380 10192
rect 18328 10149 18337 10183
rect 18337 10149 18371 10183
rect 18371 10149 18380 10183
rect 18328 10140 18380 10149
rect 19800 10140 19852 10192
rect 20444 10140 20496 10192
rect 21916 10183 21968 10192
rect 21916 10149 21925 10183
rect 21925 10149 21959 10183
rect 21959 10149 21968 10183
rect 21916 10140 21968 10149
rect 22928 10140 22980 10192
rect 24676 10140 24728 10192
rect 25044 10140 25096 10192
rect 3332 10072 3384 10124
rect 6368 10072 6420 10124
rect 20720 10072 20772 10124
rect 22008 10072 22060 10124
rect 23572 10115 23624 10124
rect 23572 10081 23581 10115
rect 23581 10081 23615 10115
rect 23615 10081 23624 10115
rect 23572 10072 23624 10081
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 1768 10004 1820 10056
rect 4068 10047 4120 10056
rect 2780 9936 2832 9988
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 3056 9936 3108 9988
rect 2688 9868 2740 9920
rect 6276 9868 6328 9920
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 16488 10004 16540 10056
rect 18696 10004 18748 10056
rect 22192 10047 22244 10056
rect 22192 10013 22201 10047
rect 22201 10013 22235 10047
rect 22235 10013 22244 10047
rect 22192 10004 22244 10013
rect 16764 9936 16816 9988
rect 6368 9868 6420 9877
rect 6736 9868 6788 9920
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 26884 9868 26936 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 3884 9664 3936 9716
rect 4068 9664 4120 9716
rect 2412 9596 2464 9648
rect 3424 9596 3476 9648
rect 2136 9528 2188 9580
rect 2964 9528 3016 9580
rect 5264 9596 5316 9648
rect 6460 9664 6512 9716
rect 7656 9596 7708 9648
rect 4344 9528 4396 9580
rect 4896 9528 4948 9580
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 6368 9528 6420 9580
rect 9588 9596 9640 9648
rect 18236 9664 18288 9716
rect 21456 9664 21508 9716
rect 22928 9664 22980 9716
rect 24768 9664 24820 9716
rect 17960 9596 18012 9648
rect 18144 9596 18196 9648
rect 19616 9639 19668 9648
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 17408 9571 17460 9580
rect 8024 9528 8076 9537
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 19616 9605 19625 9639
rect 19625 9605 19659 9639
rect 19659 9605 19668 9639
rect 19616 9596 19668 9605
rect 21824 9596 21876 9648
rect 23848 9639 23900 9648
rect 23848 9605 23857 9639
rect 23857 9605 23891 9639
rect 23891 9605 23900 9639
rect 23848 9596 23900 9605
rect 18696 9571 18748 9580
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 19708 9528 19760 9580
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 22192 9571 22244 9580
rect 20720 9528 20772 9537
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 24768 9528 24820 9580
rect 4804 9460 4856 9512
rect 5356 9460 5408 9512
rect 5448 9460 5500 9512
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 21364 9503 21416 9512
rect 21364 9469 21373 9503
rect 21373 9469 21407 9503
rect 21407 9469 21416 9503
rect 21364 9460 21416 9469
rect 21824 9460 21876 9512
rect 26700 9664 26752 9716
rect 26976 9596 27028 9648
rect 26516 9460 26568 9512
rect 27528 9503 27580 9512
rect 27528 9469 27537 9503
rect 27537 9469 27571 9503
rect 27571 9469 27580 9503
rect 27528 9460 27580 9469
rect 2044 9392 2096 9444
rect 2596 9392 2648 9444
rect 4252 9392 4304 9444
rect 4436 9392 4488 9444
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 5080 9324 5132 9376
rect 23480 9392 23532 9444
rect 5908 9324 5960 9376
rect 6000 9324 6052 9376
rect 6736 9324 6788 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 10784 9324 10836 9376
rect 14740 9324 14792 9376
rect 19984 9367 20036 9376
rect 19984 9333 19993 9367
rect 19993 9333 20027 9367
rect 20027 9333 20036 9367
rect 19984 9324 20036 9333
rect 24400 9324 24452 9376
rect 27712 9367 27764 9376
rect 27712 9333 27721 9367
rect 27721 9333 27755 9367
rect 27755 9333 27764 9367
rect 27712 9324 27764 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 2964 9120 3016 9172
rect 4160 9120 4212 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 8024 9120 8076 9172
rect 18144 9163 18196 9172
rect 18144 9129 18153 9163
rect 18153 9129 18187 9163
rect 18187 9129 18196 9163
rect 18144 9120 18196 9129
rect 18696 9120 18748 9172
rect 19984 9120 20036 9172
rect 21732 9120 21784 9172
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 23572 9163 23624 9172
rect 23572 9129 23581 9163
rect 23581 9129 23615 9163
rect 23615 9129 23624 9163
rect 23572 9120 23624 9129
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 25320 9120 25372 9172
rect 3148 8984 3200 9036
rect 6368 9052 6420 9104
rect 24860 9095 24912 9104
rect 24860 9061 24869 9095
rect 24869 9061 24903 9095
rect 24903 9061 24912 9095
rect 24860 9052 24912 9061
rect 26148 9052 26200 9104
rect 4344 8984 4396 9036
rect 4988 8984 5040 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 2964 8848 3016 8900
rect 4712 8848 4764 8900
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5448 8916 5500 8968
rect 6000 8984 6052 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 24676 8916 24728 8968
rect 2320 8780 2372 8832
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 7380 8780 7432 8832
rect 8300 8780 8352 8832
rect 26700 8823 26752 8832
rect 26700 8789 26709 8823
rect 26709 8789 26743 8823
rect 26743 8789 26752 8823
rect 26700 8780 26752 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1584 8576 1636 8628
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 3148 8508 3200 8560
rect 6276 8576 6328 8628
rect 24676 8576 24728 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25320 8576 25372 8628
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 26516 8576 26568 8628
rect 27712 8619 27764 8628
rect 27712 8585 27721 8619
rect 27721 8585 27755 8619
rect 27755 8585 27764 8619
rect 27712 8576 27764 8585
rect 2044 8440 2096 8492
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 4712 8508 4764 8560
rect 5448 8508 5500 8560
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 3608 8372 3660 8424
rect 4344 8372 4396 8424
rect 5908 8372 5960 8424
rect 6828 8372 6880 8424
rect 26608 8551 26660 8560
rect 26608 8517 26617 8551
rect 26617 8517 26651 8551
rect 26651 8517 26660 8551
rect 26608 8508 26660 8517
rect 26792 8508 26844 8560
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 8760 8440 8812 8492
rect 8392 8372 8444 8424
rect 25228 8372 25280 8424
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 2412 8347 2464 8356
rect 2412 8313 2421 8347
rect 2421 8313 2455 8347
rect 2455 8313 2464 8347
rect 2412 8304 2464 8313
rect 5724 8304 5776 8356
rect 6920 8304 6972 8356
rect 6368 8236 6420 8288
rect 8392 8236 8444 8288
rect 9036 8236 9088 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 2504 8032 2556 8084
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 2964 8032 3016 8084
rect 3608 8075 3660 8084
rect 3608 8041 3617 8075
rect 3617 8041 3651 8075
rect 3651 8041 3660 8075
rect 3608 8032 3660 8041
rect 4252 8032 4304 8084
rect 5264 8032 5316 8084
rect 6276 8032 6328 8084
rect 25872 8032 25924 8084
rect 4896 7964 4948 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2964 7896 3016 7948
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 6828 7896 6880 7948
rect 7380 7896 7432 7948
rect 25412 7896 25464 7948
rect 27252 7896 27304 7948
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 3976 7760 4028 7812
rect 6368 7760 6420 7812
rect 8300 7828 8352 7880
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 6920 7692 6972 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 26332 7692 26384 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 1400 7488 1452 7540
rect 2596 7488 2648 7540
rect 3240 7488 3292 7540
rect 4068 7488 4120 7540
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 6276 7488 6328 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 27252 7488 27304 7540
rect 1584 7463 1636 7472
rect 1584 7429 1593 7463
rect 1593 7429 1627 7463
rect 1627 7429 1636 7463
rect 1584 7420 1636 7429
rect 3976 7420 4028 7472
rect 27712 7463 27764 7472
rect 27712 7429 27721 7463
rect 27721 7429 27755 7463
rect 27755 7429 27764 7463
rect 27712 7420 27764 7429
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 6460 7352 6512 7404
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 4528 7284 4580 7336
rect 27068 7284 27120 7336
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 2964 7216 3016 7268
rect 4804 7216 4856 7268
rect 7196 7216 7248 7268
rect 9680 7216 9732 7268
rect 6368 7148 6420 7200
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 26792 7148 26844 7200
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 2872 6944 2924 6996
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 6552 6944 6604 6996
rect 6276 6876 6328 6928
rect 6736 6876 6788 6928
rect 1860 6808 1912 6860
rect 2136 6808 2188 6860
rect 2228 6808 2280 6860
rect 3516 6808 3568 6860
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5632 6808 5684 6860
rect 27436 6808 27488 6860
rect 3424 6740 3476 6792
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 1952 6672 2004 6724
rect 4160 6604 4212 6656
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1860 6400 1912 6452
rect 1584 6375 1636 6384
rect 1584 6341 1593 6375
rect 1593 6341 1627 6375
rect 1627 6341 1636 6375
rect 1584 6332 1636 6341
rect 2596 6332 2648 6384
rect 4068 6400 4120 6452
rect 5632 6400 5684 6452
rect 6276 6400 6328 6452
rect 26424 6400 26476 6452
rect 26608 6443 26660 6452
rect 26608 6409 26617 6443
rect 26617 6409 26651 6443
rect 26651 6409 26660 6443
rect 26608 6400 26660 6409
rect 27436 6400 27488 6452
rect 3332 6332 3384 6384
rect 3424 6332 3476 6384
rect 4436 6332 4488 6384
rect 3240 6264 3292 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 3792 6196 3844 6248
rect 26424 6239 26476 6248
rect 26424 6205 26433 6239
rect 26433 6205 26467 6239
rect 26467 6205 26476 6239
rect 26424 6196 26476 6205
rect 1400 6060 1452 6112
rect 1860 6060 1912 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 6368 6060 6420 6112
rect 8300 6060 8352 6112
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 2412 5788 2464 5840
rect 1768 5720 1820 5772
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 8392 5720 8444 5772
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 26700 5627 26752 5636
rect 26700 5593 26709 5627
rect 26709 5593 26743 5627
rect 26743 5593 26752 5627
rect 26700 5584 26752 5593
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2044 5355 2096 5364
rect 2044 5321 2053 5355
rect 2053 5321 2087 5355
rect 2087 5321 2096 5355
rect 2044 5312 2096 5321
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 26516 5312 26568 5364
rect 2044 5108 2096 5160
rect 26332 5108 26384 5160
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 1768 4768 1820 4820
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2044 2932 2096 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 5540 2592 5592 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 7196 2499 7248 2508
rect 7196 2465 7230 2499
rect 7230 2465 7248 2499
rect 7196 2456 7248 2465
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 938 23520 994 24000
rect 2778 23520 2834 24000
rect 3514 23624 3570 23633
rect 3514 23559 3570 23568
rect 952 20602 980 23520
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 1952 20256 2004 20262
rect 2792 20233 2820 23520
rect 3528 23458 3556 23559
rect 4618 23520 4674 24000
rect 6550 23520 6606 24000
rect 8390 23520 8446 24000
rect 10230 23520 10286 24000
rect 12162 23520 12218 24000
rect 14002 23520 14058 24000
rect 15934 23520 15990 24000
rect 17774 23520 17830 24000
rect 19614 23520 19670 24000
rect 21546 23520 21602 24000
rect 23386 23520 23442 24000
rect 24950 23624 25006 23633
rect 24950 23559 25006 23568
rect 3516 23452 3568 23458
rect 3516 23394 3568 23400
rect 3514 23080 3570 23089
rect 3514 23015 3570 23024
rect 3528 22574 3556 23015
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3238 22400 3294 22409
rect 3238 22335 3294 22344
rect 3054 20632 3110 20641
rect 3054 20567 3110 20576
rect 1952 20198 2004 20204
rect 2502 20224 2558 20233
rect 1964 19961 1992 20198
rect 2502 20159 2558 20168
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 1950 19952 2006 19961
rect 1950 19887 2006 19896
rect 1398 19816 1454 19825
rect 1398 19751 1454 19760
rect 1412 11914 1440 19751
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 18902 1992 19654
rect 2410 19544 2466 19553
rect 2410 19479 2466 19488
rect 2424 19174 2452 19479
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 1952 18896 2004 18902
rect 1952 18838 2004 18844
rect 2148 18766 2176 19110
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1596 18154 1624 18566
rect 2044 18284 2096 18290
rect 2148 18272 2176 18702
rect 2096 18244 2176 18272
rect 2044 18226 2096 18232
rect 1584 18148 1636 18154
rect 1584 18090 1636 18096
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1504 17134 1532 17614
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1596 16250 1624 18090
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 16794 1716 18022
rect 2056 17746 2084 18226
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 2042 16688 2098 16697
rect 2042 16623 2098 16632
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 2056 16114 2084 16623
rect 2240 16590 2268 17002
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 16114 2268 16526
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 1950 16008 2006 16017
rect 1950 15943 1952 15952
rect 2004 15943 2006 15952
rect 1952 15914 2004 15920
rect 1964 15706 1992 15914
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1872 14550 1900 14894
rect 1964 14822 1992 15506
rect 2056 15434 2084 16050
rect 2516 15994 2544 20159
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2688 18896 2740 18902
rect 2688 18838 2740 18844
rect 2700 18306 2728 18838
rect 2792 18426 2820 19246
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2700 18278 2820 18306
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2608 17814 2636 18022
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2240 15966 2544 15994
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 2042 15328 2098 15337
rect 2042 15263 2098 15272
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1860 14544 1912 14550
rect 1860 14486 1912 14492
rect 1872 13870 1900 14486
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13190 1900 13806
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1768 12776 1820 12782
rect 1872 12764 1900 13126
rect 1964 13025 1992 14758
rect 1950 13016 2006 13025
rect 1950 12951 2006 12960
rect 1820 12736 1900 12764
rect 1768 12718 1820 12724
rect 1872 12374 1900 12736
rect 1964 12481 1992 12951
rect 1950 12472 2006 12481
rect 1950 12407 2006 12416
rect 1860 12368 1912 12374
rect 1582 12336 1638 12345
rect 1860 12310 1912 12316
rect 1582 12271 1584 12280
rect 1636 12271 1638 12280
rect 1584 12242 1636 12248
rect 1320 11886 1440 11914
rect 1320 11234 1348 11886
rect 1398 11792 1454 11801
rect 1398 11727 1454 11736
rect 1412 11694 1440 11727
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11354 1440 11630
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1320 11206 1440 11234
rect 1412 7954 1440 11206
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7546 1440 7890
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 377 1440 6054
rect 1504 3913 1532 11494
rect 1596 8634 1624 12242
rect 2056 12102 2084 15263
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11898 2084 12038
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9722 1808 9998
rect 1950 9888 2006 9897
rect 1950 9823 2006 9832
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1582 8120 1638 8129
rect 1582 8055 1584 8064
rect 1636 8055 1638 8064
rect 1584 8026 1636 8032
rect 1766 7848 1822 7857
rect 1766 7783 1822 7792
rect 1584 7472 1636 7478
rect 1582 7440 1584 7449
rect 1636 7440 1638 7449
rect 1582 7375 1638 7384
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6730 1624 6831
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1584 6384 1636 6390
rect 1582 6352 1584 6361
rect 1636 6352 1638 6361
rect 1582 6287 1638 6296
rect 1780 5778 1808 7783
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 6458 1900 6802
rect 1964 6730 1992 9823
rect 2148 9586 2176 13126
rect 2240 12170 2268 15966
rect 2608 15638 2636 16594
rect 2700 16561 2728 16730
rect 2792 16640 2820 18278
rect 2976 18222 3004 18566
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17882 2912 18022
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 17338 3004 17682
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2964 16652 3016 16658
rect 2792 16612 2964 16640
rect 2964 16594 3016 16600
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 2700 16250 2728 16487
rect 3068 16250 3096 20567
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3160 18970 3188 19110
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3160 18222 3188 18906
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16794 3188 17002
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 2700 15881 2728 16186
rect 3068 15978 3096 16186
rect 3146 16008 3202 16017
rect 3056 15972 3108 15978
rect 3252 15994 3280 22335
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 4080 20806 4108 21791
rect 4434 21312 4490 21321
rect 4434 21247 4490 21256
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3790 19952 3846 19961
rect 3790 19887 3846 19896
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3436 16250 3464 18566
rect 3712 18358 3740 18566
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3528 16794 3556 17750
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3528 16590 3556 16730
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3528 16114 3556 16526
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3252 15966 3372 15994
rect 3146 15943 3202 15952
rect 3056 15914 3108 15920
rect 2686 15872 2742 15881
rect 2686 15807 2742 15816
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2332 14958 2360 15438
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2884 14618 2912 15438
rect 3160 15314 3188 15943
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15366 3280 15846
rect 3068 15286 3188 15314
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 13734 2820 14418
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13802 2912 14214
rect 3068 13954 3096 15286
rect 3252 15201 3280 15302
rect 3238 15192 3294 15201
rect 2976 13926 3096 13954
rect 3160 15150 3238 15178
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2424 11354 2452 13330
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12986 2636 13262
rect 2792 13190 2820 13670
rect 2780 13184 2832 13190
rect 2700 13132 2780 13138
rect 2700 13126 2832 13132
rect 2700 13110 2820 13126
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 12442 2544 12582
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 2056 8498 2084 9386
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2042 7440 2098 7449
rect 2042 7375 2044 7384
rect 2096 7375 2098 7384
rect 2044 7346 2096 7352
rect 2148 6866 2176 9522
rect 2240 9382 2268 10406
rect 2332 10266 2360 11086
rect 2516 10470 2544 12038
rect 2608 11898 2636 12922
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 6866 2268 9318
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8430 2360 8774
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1872 6118 1900 6394
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 2332 5914 2360 8366
rect 2424 8362 2452 9590
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2424 5846 2452 8298
rect 2516 8090 2544 10406
rect 2700 10010 2728 13110
rect 2884 12918 2912 13738
rect 2976 13433 3004 13926
rect 3054 13832 3110 13841
rect 3054 13767 3110 13776
rect 2962 13424 3018 13433
rect 2962 13359 3018 13368
rect 2964 13320 3016 13326
rect 3068 13297 3096 13767
rect 2964 13262 3016 13268
rect 3054 13288 3110 13297
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 10674 2820 12650
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2608 9982 2728 10010
rect 2792 9994 2820 10610
rect 2884 10146 2912 12854
rect 2976 12714 3004 13262
rect 3054 13223 3110 13232
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 3068 12322 3096 13223
rect 2976 12294 3096 12322
rect 2976 11354 3004 12294
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3068 11762 3096 12174
rect 3160 11801 3188 15150
rect 3238 15127 3294 15136
rect 3238 12880 3294 12889
rect 3238 12815 3294 12824
rect 3252 11830 3280 12815
rect 3344 11914 3372 15966
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3436 15042 3464 15914
rect 3528 15162 3556 16050
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3436 15014 3556 15042
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3436 12073 3464 12106
rect 3422 12064 3478 12073
rect 3422 11999 3478 12008
rect 3344 11886 3464 11914
rect 3240 11824 3292 11830
rect 3146 11792 3202 11801
rect 3056 11756 3108 11762
rect 3240 11766 3292 11772
rect 3146 11727 3202 11736
rect 3056 11698 3108 11704
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2976 10810 3004 11290
rect 3068 11150 3096 11698
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2884 10118 3004 10146
rect 2780 9988 2832 9994
rect 2608 9450 2636 9982
rect 2780 9930 2832 9936
rect 2688 9920 2740 9926
rect 2740 9868 2912 9874
rect 2688 9862 2912 9868
rect 2700 9846 2912 9862
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2594 9344 2650 9353
rect 2594 9279 2650 9288
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2608 7546 2636 9279
rect 2884 8974 2912 9846
rect 2976 9586 3004 10118
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9178 3004 9522
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2686 8664 2742 8673
rect 2686 8599 2742 8608
rect 2700 8090 2728 8599
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 7970 2820 8327
rect 2700 7942 2820 7970
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2596 6384 2648 6390
rect 2700 6372 2728 7942
rect 2884 7002 2912 8910
rect 2976 8906 3004 9114
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2976 8090 3004 8842
rect 3068 8634 3096 9930
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3160 8566 3188 8978
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7274 3004 7890
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2648 6344 2728 6372
rect 2596 6326 2648 6332
rect 3160 5914 3188 8502
rect 3252 7546 3280 11591
rect 3436 10266 3464 11886
rect 3528 11354 3556 15014
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3606 12472 3662 12481
rect 3606 12407 3662 12416
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3528 10606 3556 11154
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3330 10160 3386 10169
rect 3330 10095 3332 10104
rect 3384 10095 3386 10104
rect 3332 10066 3384 10072
rect 3344 9722 3372 10066
rect 3436 10033 3464 10202
rect 3422 10024 3478 10033
rect 3422 9959 3478 9968
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3344 6390 3372 9658
rect 3436 9654 3464 9959
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3528 6866 3556 10542
rect 3620 8430 3648 12407
rect 3712 12170 3740 12650
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3620 8090 3648 8366
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3606 7984 3662 7993
rect 3606 7919 3662 7928
rect 3620 7342 3648 7919
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 7002 3648 7278
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3436 6390 3464 6734
rect 3332 6384 3384 6390
rect 3238 6352 3294 6361
rect 3332 6326 3384 6332
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3238 6287 3240 6296
rect 3292 6287 3294 6296
rect 3240 6258 3292 6264
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5914 3648 6190
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 1582 5672 1638 5681
rect 1582 5607 1584 5616
rect 1636 5607 1638 5616
rect 1584 5578 1636 5584
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 5030 1624 5063
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1780 4826 1808 5714
rect 2042 5400 2098 5409
rect 2516 5370 2544 5714
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2042 5335 2044 5344
rect 2096 5335 2098 5344
rect 2504 5364 2556 5370
rect 2044 5306 2096 5312
rect 2504 5306 2556 5312
rect 2056 5166 2084 5306
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1490 3904 1546 3913
rect 1490 3839 1546 3848
rect 2042 3496 2098 3505
rect 2042 3431 2098 3440
rect 2056 3194 2084 3431
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2689 1624 2790
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 2700 1465 2728 5510
rect 3712 4457 3740 11766
rect 3804 10810 3832 19887
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4080 16794 4108 17614
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4080 14958 4108 15506
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3974 14648 4030 14657
rect 3974 14583 4030 14592
rect 3988 13705 4016 14583
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3974 13696 4030 13705
rect 3974 13631 4030 13640
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3896 10674 3924 12038
rect 4080 11121 4108 14214
rect 4172 12209 4200 18022
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4250 17640 4306 17649
rect 4250 17575 4306 17584
rect 4264 14482 4292 17575
rect 4356 17134 4384 17818
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4448 16674 4476 21247
rect 4632 19553 4660 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 4618 19544 4674 19553
rect 4618 19479 4674 19488
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4816 18970 4844 19110
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4724 18222 4752 18770
rect 4908 18630 4936 19178
rect 5092 19174 5120 19654
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4356 16646 4476 16674
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 14074 4292 14418
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4356 14006 4384 16646
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 16182 4476 16526
rect 4540 16250 4568 16730
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12345 4292 13126
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4356 12356 4384 12582
rect 4448 12424 4476 16118
rect 4632 15706 4660 16662
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4724 15586 4752 18158
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4632 15558 4752 15586
rect 4632 13297 4660 15558
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4724 14618 4752 14826
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4618 13288 4674 13297
rect 4618 13223 4674 13232
rect 4816 12889 4844 18022
rect 4908 13258 4936 18566
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5000 17882 5028 18362
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 4986 16416 5042 16425
rect 4986 16351 5042 16360
rect 5000 15978 5028 16351
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 5000 14822 5028 15506
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14414 5028 14758
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5000 13870 5028 14214
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4896 13252 4948 13258
rect 4896 13194 4948 13200
rect 4802 12880 4858 12889
rect 4802 12815 4858 12824
rect 4448 12396 4752 12424
rect 4356 12345 4476 12356
rect 4250 12336 4306 12345
rect 4356 12336 4490 12345
rect 4356 12328 4434 12336
rect 4250 12271 4306 12280
rect 4434 12271 4490 12280
rect 4158 12200 4214 12209
rect 4214 12158 4292 12186
rect 4158 12135 4214 12144
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3804 6254 3832 10610
rect 3896 9722 3924 10610
rect 4172 10554 4200 12038
rect 4264 11626 4292 12158
rect 4448 11898 4476 12271
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4264 11506 4292 11562
rect 4540 11558 4568 12174
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11552 4580 11558
rect 4264 11478 4476 11506
rect 4528 11494 4580 11500
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4264 10674 4292 11222
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4080 10538 4200 10554
rect 4068 10532 4200 10538
rect 4120 10526 4200 10532
rect 4068 10474 4120 10480
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 7818 4016 10367
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9722 4108 9998
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4068 9376 4120 9382
rect 4066 9344 4068 9353
rect 4120 9344 4122 9353
rect 4066 9279 4122 9288
rect 4172 9178 4200 10526
rect 4264 10266 4292 10610
rect 4356 10538 4384 11290
rect 4448 10826 4476 11478
rect 4448 10798 4568 10826
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4436 10464 4488 10470
rect 4434 10432 4436 10441
rect 4488 10432 4490 10441
rect 4434 10367 4490 10376
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4356 9586 4384 10134
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4080 8498 4108 9007
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4080 7954 4108 8434
rect 4264 8090 4292 9386
rect 4356 9042 4384 9522
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4344 8424 4396 8430
rect 4342 8392 4344 8401
rect 4396 8392 4398 8401
rect 4342 8327 4398 8336
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 4080 7546 4108 7890
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3698 4448 3754 4457
rect 3698 4383 3754 4392
rect 3804 3369 3832 6054
rect 3790 3360 3846 3369
rect 3790 3295 3846 3304
rect 2686 1456 2742 1465
rect 2686 1391 2742 1400
rect 3988 921 4016 7414
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4080 6458 4108 6802
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 4706 4200 6598
rect 4448 6390 4476 9386
rect 4540 7546 4568 10798
rect 4632 10742 4660 11834
rect 4724 10742 4752 12396
rect 5000 11830 5028 13806
rect 5092 12986 5120 19110
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 17066 5212 17682
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 13530 5212 15846
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5276 13326 5304 18566
rect 5368 15706 5396 19314
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5460 18426 5488 18702
rect 5644 18426 5672 18702
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 17814 5672 18226
rect 5736 18170 5764 20742
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 6564 18426 6592 23520
rect 8404 23474 8432 23520
rect 8312 23446 8432 23474
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 5814 18184 5870 18193
rect 5736 18142 5814 18170
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5644 17338 5672 17750
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5644 16794 5672 17274
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5644 15910 5672 16390
rect 5540 15904 5592 15910
rect 5632 15904 5684 15910
rect 5540 15846 5592 15852
rect 5630 15872 5632 15881
rect 5684 15872 5686 15881
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5368 14550 5396 15642
rect 5552 15609 5580 15846
rect 5630 15807 5686 15816
rect 5538 15600 5594 15609
rect 5448 15564 5500 15570
rect 5538 15535 5594 15544
rect 5448 15506 5500 15512
rect 5460 14822 5488 15506
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5368 14074 5396 14486
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5368 13462 5396 13670
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12986 5304 13262
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5368 12646 5396 13398
rect 5460 13326 5488 14758
rect 5540 14000 5592 14006
rect 5538 13968 5540 13977
rect 5592 13968 5594 13977
rect 5538 13903 5594 13912
rect 5552 13802 5580 13903
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12918 5488 13262
rect 5644 13138 5672 15807
rect 5552 13110 5672 13138
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5356 12640 5408 12646
rect 5170 12608 5226 12617
rect 5356 12582 5408 12588
rect 5170 12543 5226 12552
rect 5184 11898 5212 12543
rect 5172 11892 5224 11898
rect 5552 11880 5580 13110
rect 5630 13016 5686 13025
rect 5630 12951 5686 12960
rect 5644 12753 5672 12951
rect 5630 12744 5686 12753
rect 5630 12679 5686 12688
rect 5172 11834 5224 11840
rect 5460 11852 5580 11880
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5000 11665 5028 11766
rect 4986 11656 5042 11665
rect 4986 11591 5042 11600
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 5170 11520 5226 11529
rect 4816 11218 4844 11494
rect 5170 11455 5226 11464
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4540 7342 4568 7482
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4632 5409 4660 10542
rect 4724 9024 4752 10678
rect 4816 9518 4844 11154
rect 5184 10810 5212 11455
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5460 10674 5488 11852
rect 5538 11792 5594 11801
rect 5538 11727 5594 11736
rect 5552 11694 5580 11727
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5264 9648 5316 9654
rect 5552 9625 5580 10406
rect 5264 9590 5316 9596
rect 5538 9616 5594 9625
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4724 8996 4844 9024
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4724 8566 4752 8842
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4724 6866 4752 8502
rect 4816 7274 4844 8996
rect 4908 8974 4936 9522
rect 5080 9376 5132 9382
rect 5000 9324 5080 9330
rect 5000 9318 5132 9324
rect 5000 9302 5120 9318
rect 5000 9042 5028 9302
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 8022 4936 8910
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 5000 6866 5028 8978
rect 5276 8090 5304 9590
rect 5538 9551 5594 9560
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5368 9058 5396 9454
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5368 9030 5488 9058
rect 5460 8974 5488 9030
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8566 5488 8910
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5276 7546 5304 8026
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4618 5400 4674 5409
rect 4618 5335 4674 5344
rect 4080 4678 4200 4706
rect 4080 2145 4108 4678
rect 5460 2666 5488 8502
rect 5644 6866 5672 12679
rect 5736 8362 5764 18142
rect 5814 18119 5870 18128
rect 6472 17882 6500 18362
rect 6550 18320 6606 18329
rect 6550 18255 6606 18264
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5908 16720 5960 16726
rect 5906 16688 5908 16697
rect 5960 16688 5962 16697
rect 5906 16623 5962 16632
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 6472 16250 6500 17818
rect 6564 16425 6592 18255
rect 6840 18222 6868 18906
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6932 18068 6960 18566
rect 6748 18040 6960 18068
rect 6642 17096 6698 17105
rect 6642 17031 6698 17040
rect 6550 16416 6606 16425
rect 6550 16351 6606 16360
rect 6564 16250 6592 16351
rect 6656 16289 6684 17031
rect 6748 16794 6776 18040
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 16794 6960 16934
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6642 16280 6698 16289
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6552 16244 6604 16250
rect 6642 16215 6698 16224
rect 6552 16186 6604 16192
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5828 14618 5856 16050
rect 6564 16046 6592 16186
rect 6552 16040 6604 16046
rect 6472 16000 6552 16028
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5828 13938 5856 14554
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5828 13530 5856 13874
rect 6380 13734 6408 14214
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6380 13326 6408 13670
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6380 12646 6408 13262
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12374 6408 12582
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 11558 5856 12242
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6380 11830 6408 12310
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11354 5856 11494
rect 6288 11393 6316 11562
rect 6274 11384 6330 11393
rect 5816 11348 5868 11354
rect 6274 11319 6276 11328
rect 5816 11290 5868 11296
rect 6328 11319 6330 11328
rect 6276 11290 6328 11296
rect 6380 11150 6408 11766
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6366 10840 6422 10849
rect 6366 10775 6422 10784
rect 6380 10606 6408 10775
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9926 6408 10066
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 8838 5856 9522
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6000 9376 6052 9382
rect 6288 9353 6316 9862
rect 6380 9586 6408 9862
rect 6472 9722 6500 16000
rect 6552 15982 6604 15988
rect 6840 15892 6868 16594
rect 6920 15904 6972 15910
rect 6840 15864 6920 15892
rect 6840 15162 6868 15864
rect 6920 15846 6972 15852
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6656 11880 6684 14010
rect 6748 13394 6776 14214
rect 6840 13870 6868 14758
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6748 12714 6776 13330
rect 6840 12782 6868 13670
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6840 12442 6868 12718
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6932 12322 6960 14894
rect 7010 13696 7066 13705
rect 7010 13631 7066 13640
rect 6564 11852 6684 11880
rect 6840 12294 6960 12322
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6000 9318 6052 9324
rect 6274 9344 6330 9353
rect 5920 8945 5948 9318
rect 6012 9042 6040 9318
rect 6274 9279 6330 9288
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5906 8936 5962 8945
rect 5906 8871 5962 8880
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8498 5856 8774
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 6288 8634 6316 9279
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 5906 8528 5962 8537
rect 5816 8492 5868 8498
rect 5906 8463 5962 8472
rect 5816 8434 5868 8440
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5724 7880 5776 7886
rect 5828 7868 5856 8434
rect 5920 8430 5948 8463
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6380 8294 6408 9046
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 5776 7840 5856 7868
rect 5724 7822 5776 7828
rect 5736 7546 5764 7822
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 6288 7546 6316 8026
rect 6380 7818 6408 8230
rect 6564 7834 6592 11852
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6656 11558 6684 11698
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 11286 6684 11494
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6656 10810 6684 11222
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6748 10470 6776 11086
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 9926 6776 10406
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9382 6776 9862
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6840 8514 6868 12294
rect 7024 9058 7052 13631
rect 7116 12442 7144 20334
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 16590 7328 18022
rect 7944 17746 7972 22510
rect 8312 20618 8340 23446
rect 8220 20602 8340 20618
rect 10244 20602 10272 23520
rect 11980 23452 12032 23458
rect 11980 23394 12032 23400
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 8208 20596 8340 20602
rect 8260 20590 8340 20596
rect 10232 20596 10284 20602
rect 8208 20538 8260 20544
rect 10232 20538 10284 20544
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9218 19544 9274 19553
rect 9218 19479 9274 19488
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8128 18834 8156 19110
rect 9048 18970 9076 19246
rect 9232 19174 9260 19479
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 18086 8156 18158
rect 8588 18154 8616 18702
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15638 7328 15846
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7300 14074 7328 14486
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7300 13802 7328 14010
rect 7392 13938 7420 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11762 7144 12038
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7208 11286 7236 13126
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12306 7328 12582
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7392 11694 7420 12106
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7484 11642 7512 17274
rect 7944 17134 7972 17682
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7932 17128 7984 17134
rect 7930 17096 7932 17105
rect 7984 17096 7986 17105
rect 7930 17031 7986 17040
rect 8036 16833 8064 17478
rect 8128 17066 8156 18022
rect 8298 17776 8354 17785
rect 8298 17711 8354 17720
rect 8482 17776 8538 17785
rect 8482 17711 8538 17720
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8022 16824 8078 16833
rect 8022 16759 8078 16768
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7576 16114 7604 16458
rect 8128 16454 8156 17002
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8312 16153 8340 17711
rect 8496 17678 8524 17711
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8392 17332 8444 17338
rect 8496 17320 8524 17614
rect 8444 17292 8524 17320
rect 8392 17274 8444 17280
rect 8680 17066 8708 17614
rect 9324 17542 9352 18158
rect 9600 17762 9628 18770
rect 9692 17882 9720 18770
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9600 17734 9720 17762
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17338 9352 17478
rect 9692 17338 9720 17734
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8298 16144 8354 16153
rect 7564 16108 7616 16114
rect 8298 16079 8354 16088
rect 7564 16050 7616 16056
rect 7576 15706 7604 16050
rect 8404 16046 8432 16390
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 14958 7696 15506
rect 8312 15434 8340 15914
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8312 15162 8340 15370
rect 8404 15366 8432 15982
rect 8496 15706 8524 16526
rect 8588 16017 8616 16594
rect 8680 16590 8708 17002
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8574 16008 8630 16017
rect 9048 15978 9076 16390
rect 8574 15943 8630 15952
rect 9036 15972 9088 15978
rect 8588 15910 8616 15943
rect 9036 15914 9088 15920
rect 8576 15904 8628 15910
rect 8628 15864 8800 15892
rect 8576 15846 8628 15852
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8022 15056 8078 15065
rect 8022 14991 8078 15000
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7668 14249 7696 14894
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7654 14240 7710 14249
rect 7654 14175 7710 14184
rect 7656 12776 7708 12782
rect 7760 12753 7788 14758
rect 7944 14618 7972 14826
rect 8036 14618 8064 14991
rect 8300 14952 8352 14958
rect 8404 14940 8432 15302
rect 8496 15201 8524 15438
rect 8482 15192 8538 15201
rect 8482 15127 8538 15136
rect 8352 14912 8432 14940
rect 8300 14894 8352 14900
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8312 14346 8340 14894
rect 8392 14816 8444 14822
rect 8496 14804 8524 15127
rect 8444 14776 8524 14804
rect 8392 14758 8444 14764
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7656 12718 7708 12724
rect 7746 12744 7802 12753
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7576 11898 7604 12378
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7392 10810 7420 11630
rect 7484 11614 7604 11642
rect 7472 11552 7524 11558
rect 7470 11520 7472 11529
rect 7524 11520 7526 11529
rect 7470 11455 7526 11464
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7024 9030 7236 9058
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6472 7806 6592 7834
rect 6748 8486 6868 8514
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6380 7206 6408 7754
rect 6472 7410 6500 7806
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6458 5672 6802
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6458 6316 6870
rect 6380 6798 6408 7142
rect 6564 7002 6592 7686
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6748 6934 6776 8486
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7954 6868 8366
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6932 7750 6960 8298
rect 7208 7886 7236 9030
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8498 7420 8774
rect 7576 8537 7604 11614
rect 7668 9654 7696 12718
rect 7746 12679 7802 12688
rect 7748 12640 7800 12646
rect 7746 12608 7748 12617
rect 7800 12608 7802 12617
rect 7746 12543 7802 12552
rect 7944 12238 7972 12786
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7852 11898 7880 12174
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7944 11762 7972 12174
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8128 11286 8156 12650
rect 8220 12442 8248 13194
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12782 8432 13126
rect 8588 13025 8616 15574
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 13870 8708 14350
rect 8668 13864 8720 13870
rect 8772 13841 8800 15864
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9218 14920 9274 14929
rect 9218 14855 9274 14864
rect 9232 14074 9260 14855
rect 9508 14634 9536 15302
rect 9600 15178 9628 15370
rect 9600 15162 9720 15178
rect 9968 15162 9996 20198
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10230 19952 10286 19961
rect 10230 19887 10286 19896
rect 11888 19916 11940 19922
rect 10244 18970 10272 19887
rect 11888 19858 11940 19864
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10980 19292 11008 19654
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11060 19304 11112 19310
rect 10980 19264 11060 19292
rect 11060 19246 11112 19252
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10796 18834 10824 19110
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10888 18766 10916 18906
rect 11348 18834 11376 19314
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 10692 18760 10744 18766
rect 10690 18728 10692 18737
rect 10876 18760 10928 18766
rect 10744 18728 10746 18737
rect 10876 18702 10928 18708
rect 10690 18663 10746 18672
rect 10888 18426 10916 18702
rect 11348 18426 11376 18770
rect 11716 18630 11744 19314
rect 11900 19174 11928 19858
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18873 11928 19110
rect 11886 18864 11942 18873
rect 11886 18799 11942 18808
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10060 17134 10088 17682
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10152 16726 10180 18022
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10232 17672 10284 17678
rect 10336 17649 10364 17682
rect 10232 17614 10284 17620
rect 10322 17640 10378 17649
rect 10244 16794 10272 17614
rect 10888 17610 10916 18022
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 11532 17746 11560 18294
rect 11716 17882 11744 18566
rect 11808 18358 11836 18702
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 10322 17575 10378 17584
rect 10876 17604 10928 17610
rect 10336 17270 10364 17575
rect 10876 17546 10928 17552
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10704 17202 10732 17478
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10888 17134 10916 17546
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16833 10456 17002
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10414 16824 10470 16833
rect 10232 16788 10284 16794
rect 10956 16816 11252 16836
rect 11532 16794 11560 17274
rect 10414 16759 10416 16768
rect 10232 16730 10284 16736
rect 10468 16759 10470 16768
rect 11520 16788 11572 16794
rect 10416 16730 10468 16736
rect 11520 16730 11572 16736
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10244 16250 10272 16730
rect 10968 16720 11020 16726
rect 11020 16668 11100 16674
rect 10968 16662 11100 16668
rect 10980 16646 11100 16662
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10612 15910 10640 16526
rect 11072 16250 11100 16646
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 9600 15156 9732 15162
rect 9600 15150 9680 15156
rect 9680 15098 9732 15104
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9416 14618 9536 14634
rect 9416 14612 9548 14618
rect 9416 14606 9496 14612
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 8668 13806 8720 13812
rect 8758 13832 8814 13841
rect 8758 13767 8814 13776
rect 8574 13016 8630 13025
rect 8574 12951 8630 12960
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8036 10674 8064 11222
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7932 10600 7984 10606
rect 7930 10568 7932 10577
rect 7984 10568 7986 10577
rect 7930 10503 7986 10512
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 8036 9586 8064 10610
rect 8220 10266 8248 12242
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11801 8340 12038
rect 8298 11792 8354 11801
rect 8298 11727 8354 11736
rect 8484 11756 8536 11762
rect 8312 10742 8340 11727
rect 8484 11698 8536 11704
rect 8496 11354 8524 11698
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8772 10810 8800 13767
rect 9324 13530 9352 13874
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9310 13016 9366 13025
rect 9416 12986 9444 14606
rect 9496 14554 9548 14560
rect 9494 14512 9550 14521
rect 9494 14447 9496 14456
rect 9548 14447 9550 14456
rect 9496 14418 9548 14424
rect 10152 14414 10180 15846
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10600 15496 10652 15502
rect 10598 15464 10600 15473
rect 10652 15464 10654 15473
rect 10598 15399 10654 15408
rect 10612 15094 10640 15399
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10612 14550 10640 15030
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10140 14408 10192 14414
rect 10428 14385 10456 14418
rect 10140 14350 10192 14356
rect 10414 14376 10470 14385
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13870 10088 14214
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10152 13734 10180 14350
rect 10414 14311 10470 14320
rect 10428 13938 10456 14311
rect 10704 14074 10732 15574
rect 10796 14822 10824 15642
rect 11348 15586 11376 15846
rect 11164 15558 11376 15586
rect 11164 15065 11192 15558
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11150 15056 11206 15065
rect 11150 14991 11206 15000
rect 11164 14958 11192 14991
rect 11152 14952 11204 14958
rect 11256 14929 11284 15438
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11532 15026 11560 15302
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11152 14894 11204 14900
rect 11242 14920 11298 14929
rect 11242 14855 11244 14864
rect 11296 14855 11298 14864
rect 11244 14826 11296 14832
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9600 13433 9628 13670
rect 10428 13530 10456 13874
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9310 12951 9366 12960
rect 9404 12980 9456 12986
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 12481 8892 12582
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8956 11626 8984 12038
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8588 10266 8616 10406
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7840 9376 7892 9382
rect 7838 9344 7840 9353
rect 7892 9344 7894 9353
rect 7838 9279 7894 9288
rect 8036 9178 8064 9522
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7562 8528 7618 8537
rect 7380 8492 7432 8498
rect 7562 8463 7618 8472
rect 7380 8434 7432 8440
rect 8312 8412 8340 8774
rect 8772 8498 8800 10746
rect 9324 10538 9352 12951
rect 9404 12922 9456 12928
rect 9968 12782 9996 13126
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10046 12744 10102 12753
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11393 9720 12038
rect 9968 11898 9996 12718
rect 10520 12714 10548 13670
rect 10796 13297 10824 14758
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 11532 14618 11560 14962
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 10874 14240 10930 14249
rect 10874 14175 10930 14184
rect 10888 13977 10916 14175
rect 10874 13968 10930 13977
rect 10874 13903 10930 13912
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10046 12679 10102 12688
rect 10508 12708 10560 12714
rect 10060 12442 10088 12679
rect 10508 12650 10560 12656
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10060 11898 10088 12378
rect 10520 12238 10548 12650
rect 10888 12306 10916 13903
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11348 13530 11376 13670
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12986 11100 13126
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 11348 12374 11376 13330
rect 11440 12986 11468 13738
rect 11624 13326 11652 15914
rect 11900 15586 11928 18799
rect 11992 17338 12020 23394
rect 12176 19553 12204 23520
rect 14016 20602 14044 23520
rect 15948 23474 15976 23520
rect 15856 23446 15976 23474
rect 15856 20602 15884 23446
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 17788 20602 17816 23520
rect 19628 20602 19656 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19996 20466 20024 20742
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12162 19544 12218 19553
rect 12162 19479 12218 19488
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11992 16998 12020 17274
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12070 16144 12126 16153
rect 12070 16079 12126 16088
rect 11716 15558 11928 15586
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11532 12850 11560 13194
rect 11624 12889 11652 13262
rect 11610 12880 11666 12889
rect 11520 12844 11572 12850
rect 11610 12815 11666 12824
rect 11520 12786 11572 12792
rect 11532 12374 11560 12786
rect 11624 12646 11652 12815
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11336 12368 11388 12374
rect 11256 12328 11336 12356
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9678 11384 9734 11393
rect 9678 11319 9734 11328
rect 10244 11286 10272 12174
rect 10888 11898 10916 12242
rect 11256 12209 11284 12328
rect 11336 12310 11388 12316
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11336 12232 11388 12238
rect 11242 12200 11298 12209
rect 11336 12174 11388 12180
rect 11242 12135 11298 12144
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11348 11830 11376 12174
rect 11532 11898 11560 12310
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 10232 11280 10284 11286
rect 10428 11257 10456 11290
rect 10232 11222 10284 11228
rect 10414 11248 10470 11257
rect 9600 10674 9628 11222
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10198 9352 10474
rect 9586 10432 9642 10441
rect 9586 10367 9642 10376
rect 9036 10192 9088 10198
rect 9036 10134 9088 10140
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8392 8424 8444 8430
rect 8312 8384 8392 8412
rect 7378 8256 7434 8265
rect 7378 8191 7434 8200
rect 7392 7954 7420 8191
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7208 7274 7236 7822
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7392 7206 7420 7890
rect 8312 7886 8340 8384
rect 8392 8366 8444 8372
rect 9048 8294 9076 10134
rect 9600 10033 9628 10367
rect 9586 10024 9642 10033
rect 9586 9959 9642 9968
rect 9588 9648 9640 9654
rect 9692 9636 9720 11018
rect 9784 10470 9812 11086
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9640 9608 9720 9636
rect 9588 9590 9640 9596
rect 9784 9466 9812 10406
rect 10244 10266 10272 11222
rect 10414 11183 10470 11192
rect 10428 10470 10456 11183
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 9692 9438 9812 9466
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8404 7750 8432 8230
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6288 6361 6316 6394
rect 6274 6352 6330 6361
rect 6274 6287 6330 6296
rect 6380 6118 6408 6734
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 7392 3505 7420 7142
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7378 3496 7434 3505
rect 7378 3431 7434 3440
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 5000 2650 5580 2666
rect 8312 2650 8340 6054
rect 8404 5778 8432 7686
rect 9692 7274 9720 9438
rect 10428 8265 10456 10406
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 11716 10169 11744 15558
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11808 14958 11836 15438
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14113 11928 14758
rect 11886 14104 11942 14113
rect 12084 14074 12112 16079
rect 12176 15910 12204 16662
rect 12268 16017 12296 19994
rect 12452 19961 12480 20334
rect 12438 19952 12494 19961
rect 12438 19887 12494 19896
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12360 18154 12388 19654
rect 12636 19378 12664 19790
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12820 19310 12848 19654
rect 14844 19514 14872 20334
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17512 20058 17540 20198
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14462 19408 14518 19417
rect 14462 19343 14518 19352
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12438 18728 12494 18737
rect 12438 18663 12494 18672
rect 12452 18426 12480 18663
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12544 17338 12572 19246
rect 12820 18290 12848 19246
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12912 17882 12940 18294
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16658 12664 17002
rect 12820 16794 12848 17070
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12254 16008 12310 16017
rect 12254 15943 12310 15952
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11886 14039 11942 14048
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13870 12112 14010
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12176 13394 12204 15846
rect 12268 13530 12296 15943
rect 12360 15706 12388 16390
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12360 15570 12388 15642
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12360 14618 12388 15506
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 14521 12480 14758
rect 12438 14512 12494 14521
rect 12438 14447 12494 14456
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12452 13433 12480 13670
rect 12438 13424 12494 13433
rect 12164 13388 12216 13394
rect 12438 13359 12494 13368
rect 12164 13330 12216 13336
rect 12254 13152 12310 13161
rect 12254 13087 12310 13096
rect 12268 12714 12296 13087
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12544 11898 12572 16487
rect 12636 15745 12664 16594
rect 12820 16114 12848 16730
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13096 16046 13124 18838
rect 13372 18737 13400 19110
rect 13358 18728 13414 18737
rect 13358 18663 13414 18672
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13176 16992 13228 16998
rect 13174 16960 13176 16969
rect 13228 16960 13230 16969
rect 13174 16895 13230 16904
rect 13280 16726 13308 17478
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 13174 16552 13230 16561
rect 13174 16487 13230 16496
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12622 15736 12678 15745
rect 12622 15671 12678 15680
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12636 14414 12664 14894
rect 12728 14482 12756 14962
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 14074 12664 14350
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12636 11830 12664 14010
rect 12728 13938 12756 14418
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 12442 12756 13874
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12820 13705 12848 13738
rect 12900 13728 12952 13734
rect 12806 13696 12862 13705
rect 12900 13670 12952 13676
rect 12806 13631 12862 13640
rect 12912 13258 12940 13670
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12782 12848 13126
rect 12808 12776 12860 12782
rect 12806 12744 12808 12753
rect 12860 12744 12862 12753
rect 12806 12679 12862 12688
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 11702 10160 11758 10169
rect 11702 10095 11758 10104
rect 13004 9489 13032 14826
rect 13188 13530 13216 16487
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14482 13308 14758
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 13569 13308 14418
rect 13372 13954 13400 18663
rect 13544 18080 13596 18086
rect 13542 18048 13544 18057
rect 13636 18080 13688 18086
rect 13596 18048 13598 18057
rect 13636 18022 13688 18028
rect 13542 17983 13598 17992
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13464 17202 13492 17682
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13464 16998 13492 17138
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 15434 13492 16934
rect 13648 16658 13676 18022
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 15978 13676 16594
rect 13832 16590 13860 16730
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13634 15736 13690 15745
rect 13740 15706 13768 16526
rect 13832 15706 13860 16526
rect 14370 16416 14426 16425
rect 14370 16351 14426 16360
rect 14384 16017 14412 16351
rect 14370 16008 14426 16017
rect 14370 15943 14426 15952
rect 13634 15671 13690 15680
rect 13728 15700 13780 15706
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13372 13926 13584 13954
rect 13266 13560 13322 13569
rect 13176 13524 13228 13530
rect 13096 13484 13176 13512
rect 13096 12442 13124 13484
rect 13266 13495 13322 13504
rect 13176 13466 13228 13472
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13188 12986 13216 13262
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13096 12345 13124 12378
rect 13082 12336 13138 12345
rect 13082 12271 13138 12280
rect 12990 9480 13046 9489
rect 12990 9415 13046 9424
rect 10784 9376 10836 9382
rect 10782 9344 10784 9353
rect 10836 9344 10838 9353
rect 10782 9279 10838 9288
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 10414 8256 10470 8265
rect 10414 8191 10470 8200
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 13280 7857 13308 13495
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12850 13400 13262
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13372 7993 13400 12650
rect 13464 11121 13492 12922
rect 13556 12714 13584 13926
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13450 11112 13506 11121
rect 13450 11047 13506 11056
rect 13464 9217 13492 11047
rect 13648 10305 13676 15671
rect 13728 15642 13780 15648
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 14002 14376 14058 14385
rect 14002 14311 14004 14320
rect 14056 14311 14058 14320
rect 14004 14282 14056 14288
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 13297 14044 13670
rect 14002 13288 14058 13297
rect 14002 13223 14058 13232
rect 14278 13288 14334 13297
rect 14278 13223 14334 13232
rect 14292 12782 14320 13223
rect 14476 12986 14504 19343
rect 15120 19174 15148 19654
rect 15304 19310 15332 19654
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18329 15056 18566
rect 15014 18320 15070 18329
rect 15014 18255 15070 18264
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14936 17746 14964 18158
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14936 17134 14964 17682
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 15028 17066 15056 17818
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15120 16538 15148 19110
rect 15382 18048 15438 18057
rect 15382 17983 15438 17992
rect 15396 16658 15424 17983
rect 15488 17882 15516 19246
rect 15672 18329 15700 19858
rect 15764 19446 15792 19858
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15764 18970 15792 19382
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15752 18624 15804 18630
rect 15856 18612 15884 19790
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 16408 19281 16436 19654
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 16394 19272 16450 19281
rect 16394 19207 16450 19216
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 15804 18584 15884 18612
rect 15752 18566 15804 18572
rect 15658 18320 15714 18329
rect 15658 18255 15714 18264
rect 15764 18154 15792 18566
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15764 16998 15792 18090
rect 16316 17542 16344 18770
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15120 16510 15424 16538
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14738 16280 14794 16289
rect 15028 16250 15056 16390
rect 14738 16215 14794 16224
rect 15016 16244 15068 16250
rect 14752 16182 14780 16215
rect 15016 16186 15068 16192
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 14822 14688 15302
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14660 14414 14688 14758
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 14074 14688 14350
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 13025 14596 13126
rect 14554 13016 14610 13025
rect 14464 12980 14516 12986
rect 14554 12951 14610 12960
rect 14464 12922 14516 12928
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14568 11626 14596 12951
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 11354 14596 11562
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 13634 10296 13690 10305
rect 13634 10231 13690 10240
rect 14752 9382 14780 16118
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15016 14816 15068 14822
rect 15200 14816 15252 14822
rect 15068 14776 15148 14804
rect 15016 14758 15068 14764
rect 14832 13864 14884 13870
rect 14830 13832 14832 13841
rect 14884 13832 14886 13841
rect 14830 13767 14886 13776
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13190 14964 13670
rect 15120 13512 15148 14776
rect 15200 14758 15252 14764
rect 15212 14618 15240 14758
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15212 14074 15240 14554
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15200 13524 15252 13530
rect 15120 13484 15200 13512
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 15028 12986 15056 13330
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15120 12442 15148 13484
rect 15200 13466 15252 13472
rect 15304 13462 15332 15846
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15304 12850 15332 13398
rect 15396 13258 15424 16510
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15396 12102 15424 12310
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11762 15424 12038
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 10713 14872 11494
rect 15396 11286 15424 11698
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15488 10849 15516 15982
rect 15580 15638 15608 16186
rect 15672 15910 15700 16594
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 14618 15608 15574
rect 15764 15450 15792 16934
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 15706 15884 16526
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 15764 15422 15884 15450
rect 15750 15192 15806 15201
rect 15750 15127 15752 15136
rect 15804 15127 15806 15136
rect 15752 15098 15804 15104
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15580 13938 15608 14554
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15566 13832 15622 13841
rect 15566 13767 15568 13776
rect 15620 13767 15622 13776
rect 15568 13738 15620 13744
rect 15580 11354 15608 13738
rect 15672 12850 15700 15030
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 13977 15792 14758
rect 15750 13968 15806 13977
rect 15750 13903 15806 13912
rect 15856 13326 15884 15422
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16316 15094 16344 15642
rect 16408 15314 16436 18566
rect 16500 18442 16528 19314
rect 16854 19272 16910 19281
rect 16854 19207 16856 19216
rect 16908 19207 16910 19216
rect 16856 19178 16908 19184
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16500 18426 16620 18442
rect 16500 18420 16632 18426
rect 16500 18414 16580 18420
rect 16580 18362 16632 18368
rect 16592 17814 16620 18362
rect 16684 18086 16712 18634
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16580 17808 16632 17814
rect 16580 17750 16632 17756
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 16726 16528 17614
rect 16592 17338 16620 17750
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 17270 16712 17682
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16776 17105 16804 19110
rect 16854 18320 16910 18329
rect 16854 18255 16910 18264
rect 16762 17096 16818 17105
rect 16762 17031 16818 17040
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16868 16658 16896 18255
rect 17314 17640 17370 17649
rect 17314 17575 17370 17584
rect 17328 16794 17356 17575
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17224 16720 17276 16726
rect 17328 16697 17356 16730
rect 17224 16662 17276 16668
rect 17314 16688 17370 16697
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16486 16416 16542 16425
rect 16486 16351 16542 16360
rect 16500 16250 16528 16351
rect 17236 16250 17264 16662
rect 17314 16623 17370 16632
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 16182 17356 16623
rect 17420 16590 17448 19314
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18426 17540 18702
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 16408 15286 16620 15314
rect 16592 15162 16620 15286
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16670 14648 16726 14657
rect 16670 14583 16726 14592
rect 16684 14550 16712 14583
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16408 13734 16436 14350
rect 16684 14074 16712 14486
rect 16776 14385 16804 14758
rect 16762 14376 16818 14385
rect 16762 14311 16818 14320
rect 16868 14113 16896 14894
rect 16960 14618 16988 14962
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16854 14104 16910 14113
rect 16672 14068 16724 14074
rect 16854 14039 16910 14048
rect 16672 14010 16724 14016
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12986 15884 13262
rect 16394 13152 16450 13161
rect 15956 13084 16252 13104
rect 16394 13087 16450 13096
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 12442 15700 12786
rect 16408 12782 16436 13087
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 15842 12472 15898 12481
rect 15660 12436 15712 12442
rect 15842 12407 15898 12416
rect 15660 12378 15712 12384
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15474 10840 15530 10849
rect 15580 10810 15608 11290
rect 15474 10775 15530 10784
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 14830 10704 14886 10713
rect 14830 10639 14886 10648
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 13450 9208 13506 9217
rect 13450 9143 13506 9152
rect 13358 7984 13414 7993
rect 13358 7919 13414 7928
rect 13266 7848 13322 7857
rect 13266 7783 13322 7792
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 9692 5273 9720 7210
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 14752 6225 14780 9318
rect 15856 7449 15884 12407
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 16316 11393 16344 12038
rect 16500 11558 16528 12582
rect 16684 12442 16712 14010
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16868 12986 16896 13398
rect 17052 13297 17080 15914
rect 17420 15706 17448 16526
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13326 17172 13670
rect 17132 13320 17184 13326
rect 17038 13288 17094 13297
rect 17132 13262 17184 13268
rect 17038 13223 17094 13232
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 12374 16804 12650
rect 16764 12368 16816 12374
rect 16762 12336 16764 12345
rect 16816 12336 16818 12345
rect 16672 12300 16724 12306
rect 16868 12322 16896 12922
rect 17144 12646 17172 13262
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 16868 12294 17080 12322
rect 16762 12271 16818 12280
rect 16672 12242 16724 12248
rect 16684 12209 16712 12242
rect 16670 12200 16726 12209
rect 16670 12135 16726 12144
rect 16684 11898 16712 12135
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16776 11830 16804 12271
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16868 11626 16896 12106
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16302 11384 16358 11393
rect 16408 11354 16436 11494
rect 16302 11319 16358 11328
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16500 11150 16528 11222
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16500 10810 16528 11086
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16500 10062 16528 10746
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16776 9994 16804 11494
rect 16960 11286 16988 12174
rect 17052 11762 17080 12294
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17420 11558 17448 11698
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16960 11082 16988 11222
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10470 16896 10950
rect 17420 10742 17448 11494
rect 17604 11354 17632 20334
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 18050 19952 18106 19961
rect 17960 19916 18012 19922
rect 18050 19887 18106 19896
rect 17960 19858 18012 19864
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17696 18766 17724 19246
rect 17868 19168 17920 19174
rect 17972 19156 18000 19858
rect 17920 19128 18000 19156
rect 17868 19110 17920 19116
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17696 18086 17724 18702
rect 17880 18426 17908 19110
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17696 17746 17724 18022
rect 17788 17864 17816 18362
rect 17960 17876 18012 17882
rect 17788 17836 17960 17864
rect 17960 17818 18012 17824
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17696 17134 17724 17682
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17696 16590 17724 17070
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 16114 17724 16526
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17960 15632 18012 15638
rect 17880 15580 17960 15586
rect 17880 15574 18012 15580
rect 17880 15558 18000 15574
rect 17880 15162 17908 15558
rect 18064 15314 18092 19887
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18234 19408 18290 19417
rect 18234 19343 18290 19352
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18156 18290 18184 18770
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18248 17513 18276 19343
rect 18340 19174 18368 19722
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18970 18368 19110
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18234 17504 18290 17513
rect 18234 17439 18290 17448
rect 18248 16658 18276 17439
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18248 16250 18276 16594
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 17972 15286 18092 15314
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13462 17816 14214
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17866 12744 17922 12753
rect 17866 12679 17868 12688
rect 17920 12679 17922 12688
rect 17868 12650 17920 12656
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12238 17816 12582
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17788 11762 17816 12174
rect 17880 11898 17908 12310
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17880 11608 17908 11834
rect 17972 11830 18000 15286
rect 18248 15094 18276 16050
rect 18340 15978 18368 18906
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18524 17066 18552 17818
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18432 15706 18460 16662
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18050 13968 18106 13977
rect 18050 13903 18106 13912
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18064 11778 18092 13903
rect 18064 11750 18184 11778
rect 17880 11580 18092 11608
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17788 10690 17816 11562
rect 17880 10810 17908 11580
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17972 10826 18000 11222
rect 18064 11150 18092 11580
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17972 10810 18092 10826
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17960 10804 18092 10810
rect 18012 10798 18092 10804
rect 17960 10746 18012 10752
rect 17788 10662 18000 10690
rect 17406 10568 17462 10577
rect 17406 10503 17462 10512
rect 16856 10464 16908 10470
rect 16854 10432 16856 10441
rect 16908 10432 16910 10441
rect 16854 10367 16910 10376
rect 17420 10198 17448 10503
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 17420 9586 17448 10134
rect 17972 9654 18000 10662
rect 18064 10266 18092 10798
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18156 9654 18184 11750
rect 18248 10266 18276 14758
rect 18524 14074 18552 17002
rect 18616 16969 18644 20198
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18708 19174 18736 19858
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18708 17882 18736 19110
rect 19352 18154 19380 20198
rect 19444 19854 19472 20266
rect 19432 19848 19484 19854
rect 19430 19816 19432 19825
rect 19484 19816 19486 19825
rect 19430 19751 19486 19760
rect 19996 19242 20024 20402
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20732 19258 20760 20334
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 20548 19230 20760 19258
rect 19996 18630 20024 19178
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20166 18728 20222 18737
rect 20166 18663 20222 18672
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19904 18426 19932 18566
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 19444 17814 19472 18226
rect 19904 18222 19932 18362
rect 19996 18290 20024 18566
rect 20180 18358 20208 18663
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 18984 17542 19012 17682
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18602 16960 18658 16969
rect 18602 16895 18658 16904
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 13705 18552 13806
rect 18510 13696 18566 13705
rect 18510 13631 18566 13640
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18418 12744 18474 12753
rect 18418 12679 18474 12688
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18248 9722 18276 10202
rect 18340 10198 18368 11766
rect 18432 11762 18460 12679
rect 18524 12374 18552 13126
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18616 11801 18644 16895
rect 18984 16794 19012 17478
rect 19444 16794 19472 17750
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19812 16794 19840 17546
rect 19892 16992 19944 16998
rect 19996 16980 20024 18226
rect 20180 18154 20208 18294
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 20456 17678 20484 19110
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 19944 16952 20024 16980
rect 19892 16934 19944 16940
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18878 15600 18934 15609
rect 18788 15564 18840 15570
rect 18878 15535 18934 15544
rect 18788 15506 18840 15512
rect 18800 14618 18828 15506
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18800 12986 18828 14554
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18892 11937 18920 15535
rect 18984 15502 19012 16458
rect 19076 15978 19104 16594
rect 19904 16590 19932 16934
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19430 16280 19486 16289
rect 19430 16215 19486 16224
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 15162 19012 15438
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18984 13954 19012 14418
rect 19076 14074 19104 15914
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19352 14890 19380 15846
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19352 14346 19380 14826
rect 19444 14482 19472 16215
rect 20166 15056 20222 15065
rect 20166 14991 20222 15000
rect 19706 14920 19762 14929
rect 19706 14855 19762 14864
rect 19720 14618 19748 14855
rect 19708 14612 19760 14618
rect 19628 14572 19708 14600
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19246 14240 19248 14249
rect 19300 14240 19302 14249
rect 19246 14175 19302 14184
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18984 13926 19104 13954
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18878 11928 18934 11937
rect 18878 11863 18934 11872
rect 18602 11792 18658 11801
rect 18420 11756 18472 11762
rect 18602 11727 18658 11736
rect 18420 11698 18472 11704
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18418 10704 18474 10713
rect 18524 10674 18552 11154
rect 18418 10639 18474 10648
rect 18512 10668 18564 10674
rect 18432 10606 18460 10639
rect 18512 10610 18564 10616
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 10266 18460 10542
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 17960 9648 18012 9654
rect 17774 9616 17830 9625
rect 17408 9580 17460 9586
rect 17960 9590 18012 9596
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 17774 9551 17776 9560
rect 17408 9522 17460 9528
rect 17828 9551 17830 9560
rect 17776 9522 17828 9528
rect 18156 9178 18184 9590
rect 18708 9586 18736 9998
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 18432 8537 18460 9454
rect 18708 9178 18736 9522
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18418 8528 18474 8537
rect 18418 8463 18474 8472
rect 18984 7857 19012 13806
rect 19076 13802 19104 13926
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 19076 13569 19104 13738
rect 19062 13560 19118 13569
rect 19062 13495 19118 13504
rect 19168 12850 19196 13874
rect 19536 13870 19564 14418
rect 19524 13864 19576 13870
rect 19522 13832 19524 13841
rect 19576 13832 19578 13841
rect 19522 13767 19578 13776
rect 19628 13462 19656 14572
rect 19708 14554 19760 14560
rect 19892 14408 19944 14414
rect 20180 14385 20208 14991
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20364 14618 20392 14826
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14657 20484 14758
rect 20442 14648 20498 14657
rect 20352 14612 20404 14618
rect 20442 14583 20498 14592
rect 20352 14554 20404 14560
rect 20258 14512 20314 14521
rect 20258 14447 20314 14456
rect 19892 14350 19944 14356
rect 20166 14376 20222 14385
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19338 13288 19394 13297
rect 19338 13223 19394 13232
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19352 12764 19380 13223
rect 19260 12736 19380 12764
rect 19260 12646 19288 12736
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11626 19196 12038
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19168 11082 19196 11562
rect 19246 11520 19302 11529
rect 19246 11455 19302 11464
rect 19260 11354 19288 11455
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19260 10810 19288 11154
rect 19352 10810 19380 12736
rect 19614 11928 19670 11937
rect 19614 11863 19670 11872
rect 19628 11354 19656 11863
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19614 10432 19670 10441
rect 19614 10367 19670 10376
rect 19628 9654 19656 10367
rect 19720 10266 19748 14214
rect 19904 13841 19932 14350
rect 20166 14311 20222 14320
rect 20074 14104 20130 14113
rect 20074 14039 20076 14048
rect 20128 14039 20130 14048
rect 20076 14010 20128 14016
rect 20088 13870 20116 14010
rect 20076 13864 20128 13870
rect 19890 13832 19946 13841
rect 20076 13806 20128 13812
rect 19890 13767 19946 13776
rect 19904 13530 19932 13767
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19812 11286 19840 12650
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19720 9586 19748 10202
rect 19812 10198 19840 11222
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19996 9382 20024 13466
rect 20088 9897 20116 13806
rect 20180 13802 20208 14311
rect 20272 14074 20300 14447
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20364 13938 20392 14554
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 20180 13530 20208 13738
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20180 11150 20208 11494
rect 20258 11384 20314 11393
rect 20258 11319 20260 11328
rect 20312 11319 20314 11328
rect 20260 11290 20312 11296
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20180 10674 20208 11086
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20272 10606 20300 11290
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20456 10198 20484 13262
rect 20548 12986 20576 19230
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 18222 20760 18702
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20628 17876 20680 17882
rect 20732 17864 20760 18158
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 18057 21404 18090
rect 21362 18048 21418 18057
rect 20956 17980 21252 18000
rect 21362 17983 21418 17992
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 20680 17836 20760 17864
rect 20628 17818 20680 17824
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21376 17338 21404 17682
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21284 16250 21312 16594
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 21284 14618 21312 16186
rect 21376 16114 21404 17274
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21376 15706 21404 16050
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21362 15464 21418 15473
rect 21468 15450 21496 20742
rect 21560 20602 21588 23520
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 23400 19514 23428 23520
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 20262 23888 20946
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 22558 19272 22614 19281
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21652 18222 21680 18770
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21640 18216 21692 18222
rect 21638 18184 21640 18193
rect 21692 18184 21694 18193
rect 21638 18119 21694 18128
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16590 21588 16934
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21418 15422 21496 15450
rect 21362 15399 21418 15408
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21284 13734 21312 14350
rect 21376 13818 21404 15399
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21468 14958 21496 15302
rect 21652 15162 21680 17002
rect 21744 16726 21772 18294
rect 21836 17338 21864 19246
rect 22558 19207 22614 19216
rect 22466 19136 22522 19145
rect 22466 19071 22522 19080
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21928 17882 21956 18090
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21836 16250 21864 17070
rect 22112 16810 22140 18566
rect 22480 18290 22508 19071
rect 22572 18970 22600 19207
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22572 18426 22600 18906
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22664 18290 22692 18702
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22480 17882 22508 18226
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 17338 22232 17614
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22204 16998 22232 17274
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22020 16794 22232 16810
rect 22008 16788 22232 16794
rect 22060 16782 22232 16788
rect 22008 16730 22060 16736
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21928 15910 21956 16390
rect 22112 16046 22140 16662
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22204 15910 22232 16782
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 21730 15736 21786 15745
rect 21730 15671 21786 15680
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21560 14414 21588 15030
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21744 13954 21772 15671
rect 21928 15502 21956 15846
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21928 15094 21956 15438
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21836 14074 21864 14894
rect 21928 14890 21956 15030
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 22204 14822 22232 15506
rect 22192 14816 22244 14822
rect 21914 14784 21970 14793
rect 22192 14758 22244 14764
rect 21914 14719 21970 14728
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21744 13926 21864 13954
rect 21376 13790 21772 13818
rect 21272 13728 21324 13734
rect 20810 13696 20866 13705
rect 21272 13670 21324 13676
rect 20810 13631 20866 13640
rect 20824 13512 20852 13631
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20824 13484 20944 13512
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20732 12850 20760 13126
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 12238 20668 12582
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20640 11778 20668 12174
rect 20732 11898 20760 12786
rect 20824 12442 20852 13330
rect 20916 12986 20944 13484
rect 21180 13320 21232 13326
rect 21284 13274 21312 13670
rect 21232 13268 21312 13274
rect 21180 13262 21312 13268
rect 21192 13246 21312 13262
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21008 12850 21036 13126
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 21284 12374 21312 13246
rect 21364 12912 21416 12918
rect 21362 12880 21364 12889
rect 21416 12880 21418 12889
rect 21362 12815 21418 12824
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20640 11750 20760 11778
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20548 10538 20576 11630
rect 20732 10810 20760 11750
rect 21192 11642 21220 12242
rect 21284 11830 21312 12310
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21362 11792 21418 11801
rect 21362 11727 21418 11736
rect 20812 11620 20864 11626
rect 21192 11614 21312 11642
rect 20812 11562 20864 11568
rect 20824 11529 20852 11562
rect 21284 11558 21312 11614
rect 21272 11552 21324 11558
rect 20810 11520 20866 11529
rect 21272 11494 21324 11500
rect 20810 11455 20866 11464
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 21376 11218 21404 11727
rect 21454 11656 21510 11665
rect 21454 11591 21510 11600
rect 21468 11354 21496 11591
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21180 11008 21232 11014
rect 21180 10950 21232 10956
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 21192 10674 21220 10950
rect 21376 10742 21404 11154
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20732 10470 20760 10610
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20732 10130 20760 10406
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20074 9888 20130 9897
rect 20074 9823 20130 9832
rect 20088 9518 20116 9823
rect 20732 9586 20760 10066
rect 21468 9722 21496 10610
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 10266 21588 10406
rect 21744 10266 21772 13790
rect 21836 12073 21864 13926
rect 21928 12986 21956 14719
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22112 13870 22140 14418
rect 22204 14278 22232 14758
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22006 13424 22062 13433
rect 22006 13359 22062 13368
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22020 12782 22048 13359
rect 22112 13190 22140 13806
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22098 13016 22154 13025
rect 22098 12951 22154 12960
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21822 12064 21878 12073
rect 21822 11999 21878 12008
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20076 9512 20128 9518
rect 21364 9512 21416 9518
rect 20076 9454 20128 9460
rect 21362 9480 21364 9489
rect 21416 9480 21418 9489
rect 21362 9415 21418 9424
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9178 20024 9318
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 21744 9178 21772 10202
rect 21836 9654 21864 11999
rect 22020 11762 22048 12378
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11354 22048 11698
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22020 10674 22048 11290
rect 22112 11257 22140 12951
rect 22204 12850 22232 14214
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12374 22232 12786
rect 22192 12368 22244 12374
rect 22192 12310 22244 12316
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22204 11354 22232 11562
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22098 11248 22154 11257
rect 22098 11183 22154 11192
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21836 9518 21864 9590
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21928 9178 21956 10134
rect 22020 10130 22048 10610
rect 22296 10146 22324 17818
rect 22664 17814 22692 18226
rect 23400 18204 23428 18770
rect 23400 18176 23704 18204
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22664 16658 22692 17750
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23032 16794 23060 17682
rect 23400 17338 23428 18022
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23400 17066 23428 17274
rect 23388 17060 23440 17066
rect 23388 17002 23440 17008
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22388 15706 22416 15982
rect 22664 15706 22692 16594
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 22388 15026 22416 15642
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22664 13938 22692 15642
rect 23400 15162 23428 15642
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23492 14929 23520 18022
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23584 17202 23612 17478
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23478 14920 23534 14929
rect 23478 14855 23534 14864
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 23216 13802 23244 14282
rect 23492 14074 23520 14554
rect 23676 14385 23704 18176
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23768 15065 23796 17478
rect 23754 15056 23810 15065
rect 23754 14991 23810 15000
rect 23662 14376 23718 14385
rect 23662 14311 23718 14320
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23492 13977 23520 14010
rect 23478 13968 23534 13977
rect 23478 13903 23534 13912
rect 23662 13832 23718 13841
rect 23204 13796 23256 13802
rect 23662 13767 23664 13776
rect 23204 13738 23256 13744
rect 23716 13767 23718 13776
rect 23664 13738 23716 13744
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22480 13161 22508 13670
rect 23216 13530 23244 13738
rect 23676 13530 23704 13738
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 22466 13152 22522 13161
rect 22466 13087 22522 13096
rect 22376 12640 22428 12646
rect 22374 12608 22376 12617
rect 22428 12608 22430 12617
rect 22374 12543 22430 12552
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22112 10118 22324 10146
rect 22112 9602 22140 10118
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22020 9574 22140 9602
rect 22204 9586 22232 9998
rect 22192 9580 22244 9586
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22020 8809 22048 9574
rect 22192 9522 22244 9528
rect 22006 8800 22062 8809
rect 22006 8735 22062 8744
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 18970 7848 19026 7857
rect 18970 7783 19026 7792
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 22480 7449 22508 13087
rect 23032 12986 23060 13330
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23492 11937 23520 12242
rect 23478 11928 23534 11937
rect 23478 11863 23480 11872
rect 23532 11863 23534 11872
rect 23480 11834 23532 11840
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22652 11280 22704 11286
rect 22652 11222 22704 11228
rect 22664 10266 22692 11222
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22940 10810 22968 11086
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22940 10198 22968 10746
rect 23032 10266 23060 11290
rect 23584 11218 23612 12922
rect 23768 12481 23796 14991
rect 23754 12472 23810 12481
rect 23754 12407 23810 12416
rect 23754 11792 23810 11801
rect 23754 11727 23756 11736
rect 23808 11727 23810 11736
rect 23756 11698 23808 11704
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 23124 10810 23152 10950
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 22940 9722 22968 10134
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 23400 9466 23428 11018
rect 23584 10674 23612 11154
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23492 10266 23520 10474
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23584 10130 23612 10610
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23400 9450 23520 9466
rect 23400 9444 23532 9450
rect 23400 9438 23480 9444
rect 23480 9386 23532 9392
rect 23584 9178 23612 10066
rect 23860 9654 23888 20198
rect 24044 19514 24072 20198
rect 24964 19802 24992 23559
rect 25226 23520 25282 24000
rect 27158 23520 27214 24000
rect 28998 23520 29054 24000
rect 25134 21312 25190 21321
rect 25134 21247 25190 21256
rect 25148 20806 25176 21247
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25240 20602 25268 23520
rect 25318 23080 25374 23089
rect 25318 23015 25374 23024
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25332 20346 25360 23015
rect 25410 22400 25466 22409
rect 25410 22335 25466 22344
rect 24872 19774 24992 19802
rect 25056 20318 25360 20346
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 24216 19304 24268 19310
rect 24216 19246 24268 19252
rect 24228 18902 24256 19246
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24504 18970 24532 19110
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24216 18896 24268 18902
rect 24216 18838 24268 18844
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23952 18154 23980 18702
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 24216 18148 24268 18154
rect 24216 18090 24268 18096
rect 23938 17096 23994 17105
rect 23938 17031 23994 17040
rect 24032 17060 24084 17066
rect 23952 12782 23980 17031
rect 24032 17002 24084 17008
rect 24044 16794 24072 17002
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 24044 16250 24072 16730
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24032 15428 24084 15434
rect 24032 15370 24084 15376
rect 24044 14890 24072 15370
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 24044 14793 24072 14826
rect 24136 14822 24164 15302
rect 24124 14816 24176 14822
rect 24030 14784 24086 14793
rect 24124 14758 24176 14764
rect 24030 14719 24086 14728
rect 24032 14544 24084 14550
rect 24136 14521 24164 14758
rect 24032 14486 24084 14492
rect 24122 14512 24178 14521
rect 24044 13870 24072 14486
rect 24122 14447 24178 14456
rect 24228 14362 24256 18090
rect 24400 18080 24452 18086
rect 24306 18048 24362 18057
rect 24400 18022 24452 18028
rect 24306 17983 24362 17992
rect 24136 14334 24256 14362
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 12776 23992 12782
rect 24044 12753 24072 13806
rect 23940 12718 23992 12724
rect 24030 12744 24086 12753
rect 24030 12679 24086 12688
rect 23940 12368 23992 12374
rect 23940 12310 23992 12316
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23952 8945 23980 12310
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 24044 11286 24072 11494
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 24136 10146 24164 14334
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24228 12442 24256 14010
rect 24320 12866 24348 17983
rect 24412 17542 24440 18022
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24504 15978 24532 18906
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24688 18290 24716 18566
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24688 16250 24716 18226
rect 24872 18057 24900 19774
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24858 18048 24914 18057
rect 24858 17983 24914 17992
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24780 16658 24808 17546
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24674 16144 24730 16153
rect 24674 16079 24730 16088
rect 24492 15972 24544 15978
rect 24492 15914 24544 15920
rect 24688 15609 24716 16079
rect 24398 15600 24454 15609
rect 24398 15535 24454 15544
rect 24674 15600 24730 15609
rect 24780 15586 24808 16594
rect 24872 15706 24900 16662
rect 24964 16658 24992 19654
rect 25056 16697 25084 20318
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25240 19922 25268 20198
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25148 19378 25176 19722
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25240 19009 25268 19858
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25226 19000 25282 19009
rect 25332 18970 25360 19314
rect 25424 19122 25452 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25502 21584 25558 21593
rect 25502 21519 25558 21528
rect 25516 19281 25544 21519
rect 27172 21146 27200 23520
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 29012 21078 29040 23520
rect 29000 21072 29052 21078
rect 29000 21014 29052 21020
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 25700 20330 25728 20742
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25688 20324 25740 20330
rect 25688 20266 25740 20272
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25608 19990 25636 20198
rect 25596 19984 25648 19990
rect 25596 19926 25648 19932
rect 25608 19310 25636 19926
rect 25792 19854 25820 20402
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25792 19446 25820 19790
rect 25884 19718 25912 20198
rect 26160 19802 26188 20198
rect 26516 19848 26568 19854
rect 26160 19774 26372 19802
rect 26516 19790 26568 19796
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25884 19514 25912 19654
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 25780 19440 25832 19446
rect 25832 19388 25912 19394
rect 25780 19382 25912 19388
rect 25792 19366 25912 19382
rect 25792 19317 25820 19366
rect 25596 19304 25648 19310
rect 25502 19272 25558 19281
rect 25596 19246 25648 19252
rect 25502 19207 25558 19216
rect 25596 19168 25648 19174
rect 25424 19116 25596 19122
rect 25424 19110 25648 19116
rect 25424 19094 25636 19110
rect 25226 18935 25282 18944
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25410 18864 25466 18873
rect 25410 18799 25466 18808
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25134 17776 25190 17785
rect 25134 17711 25190 17720
rect 25042 16688 25098 16697
rect 24952 16652 25004 16658
rect 25042 16623 25098 16632
rect 24952 16594 25004 16600
rect 24950 15872 25006 15881
rect 24950 15807 25006 15816
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24780 15558 24900 15586
rect 24674 15535 24730 15544
rect 24412 14074 24440 15535
rect 24582 15192 24638 15201
rect 24582 15127 24638 15136
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24412 13462 24440 13806
rect 24400 13456 24452 13462
rect 24400 13398 24452 13404
rect 24412 12986 24440 13398
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24320 12838 24440 12866
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24228 11762 24256 12378
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24412 11354 24440 12838
rect 24596 12374 24624 15127
rect 24766 13832 24822 13841
rect 24766 13767 24768 13776
rect 24820 13767 24822 13776
rect 24768 13738 24820 13744
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24688 13297 24716 13330
rect 24674 13288 24730 13297
rect 24674 13223 24730 13232
rect 24688 12442 24716 13223
rect 24872 13161 24900 15558
rect 24964 14618 24992 15807
rect 25148 15722 25176 17711
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25240 16658 25268 17478
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25056 15694 25176 15722
rect 25056 15609 25084 15694
rect 25042 15600 25098 15609
rect 25042 15535 25098 15544
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25056 14822 25084 15438
rect 25148 14822 25176 15506
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24858 13152 24914 13161
rect 24858 13087 24914 13096
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24596 11762 24624 12106
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24412 10810 24440 11290
rect 24596 11150 24624 11698
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24596 10538 24624 11086
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 24688 10418 24716 12038
rect 24872 11830 24900 12718
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24596 10390 24716 10418
rect 24214 10160 24270 10169
rect 24136 10118 24214 10146
rect 24136 9897 24164 10118
rect 24214 10095 24270 10104
rect 24122 9888 24178 9897
rect 24122 9823 24178 9832
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24412 9178 24440 9318
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 23938 8936 23994 8945
rect 23938 8871 23994 8880
rect 24596 8242 24624 10390
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24688 8974 24716 10134
rect 24780 9722 24808 11154
rect 24964 11121 24992 12854
rect 25056 12345 25084 14758
rect 25148 12889 25176 14758
rect 25240 14618 25268 16594
rect 25332 16590 25360 18022
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25332 15638 25360 16526
rect 25424 16153 25452 18799
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25516 17066 25544 17614
rect 25504 17060 25556 17066
rect 25504 17002 25556 17008
rect 25516 16794 25544 17002
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25608 16674 25636 19094
rect 25884 18426 25912 19366
rect 26344 18970 26372 19774
rect 26528 19310 26556 19790
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26422 19000 26478 19009
rect 26332 18964 26384 18970
rect 26422 18935 26478 18944
rect 26332 18906 26384 18912
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26252 17882 26280 18090
rect 26240 17876 26292 17882
rect 26344 17864 26372 18702
rect 26292 17836 26372 17864
rect 26240 17818 26292 17824
rect 25686 17640 25742 17649
rect 25686 17575 25742 17584
rect 25516 16646 25636 16674
rect 25410 16144 25466 16153
rect 25410 16079 25466 16088
rect 25412 15972 25464 15978
rect 25412 15914 25464 15920
rect 25320 15632 25372 15638
rect 25320 15574 25372 15580
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25226 14376 25282 14385
rect 25226 14311 25282 14320
rect 25134 12880 25190 12889
rect 25134 12815 25190 12824
rect 25042 12336 25098 12345
rect 25148 12306 25176 12815
rect 25042 12271 25098 12280
rect 25136 12300 25188 12306
rect 25056 12238 25084 12271
rect 25136 12242 25188 12248
rect 25044 12232 25096 12238
rect 25148 12209 25176 12242
rect 25044 12174 25096 12180
rect 25134 12200 25190 12209
rect 25056 11898 25084 12174
rect 25134 12135 25190 12144
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25056 11257 25084 11834
rect 25148 11354 25176 12135
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25042 11248 25098 11257
rect 25042 11183 25098 11192
rect 24950 11112 25006 11121
rect 24950 11047 25006 11056
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 25056 10198 25084 10406
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24964 9602 24992 9862
rect 24780 9586 24992 9602
rect 24768 9580 24992 9586
rect 24820 9574 24992 9580
rect 24768 9522 24820 9528
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24688 8634 24716 8910
rect 24872 8634 24900 9046
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24596 8214 24900 8242
rect 15842 7440 15898 7449
rect 15842 7375 15898 7384
rect 22466 7440 22522 7449
rect 22466 7375 22522 7384
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 14738 6216 14794 6225
rect 14738 6151 14794 6160
rect 24766 6216 24822 6225
rect 24766 6151 24822 6160
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 9678 5264 9734 5273
rect 9678 5199 9734 5208
rect 24780 5137 24808 6151
rect 24766 5128 24822 5137
rect 24766 5063 24822 5072
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 24872 4593 24900 8214
rect 24858 4584 24914 4593
rect 24858 4519 24914 4528
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 5000 2644 5592 2650
rect 5000 2638 5540 2644
rect 4066 2136 4122 2145
rect 4066 2071 4122 2080
rect 3974 912 4030 921
rect 3974 847 4030 856
rect 5000 480 5028 2638
rect 5540 2586 5592 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7208 2417 7236 2450
rect 7194 2408 7250 2417
rect 7194 2343 7250 2352
rect 14922 2408 14978 2417
rect 14922 2343 14978 2352
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 14936 480 14964 2343
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 24964 480 24992 9574
rect 25240 8430 25268 14311
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25332 12782 25360 13466
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 25332 12442 25360 12718
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25424 12374 25452 15914
rect 25516 15201 25544 16646
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25608 15910 25636 16526
rect 25700 16289 25728 17575
rect 25778 17504 25834 17513
rect 25778 17439 25834 17448
rect 25792 17338 25820 17439
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 26344 17270 26372 17836
rect 26436 17338 26464 18935
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 26332 17264 26384 17270
rect 26332 17206 26384 17212
rect 25778 17096 25834 17105
rect 25778 17031 25834 17040
rect 26424 17060 26476 17066
rect 25792 16425 25820 17031
rect 26424 17002 26476 17008
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 25872 16720 25924 16726
rect 25872 16662 25924 16668
rect 25778 16416 25834 16425
rect 25778 16351 25834 16360
rect 25686 16280 25742 16289
rect 25686 16215 25742 16224
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25608 15745 25636 15846
rect 25594 15736 25650 15745
rect 25594 15671 25650 15680
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25502 15192 25558 15201
rect 25502 15127 25558 15136
rect 25608 15094 25636 15574
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25700 15162 25728 15506
rect 25792 15434 25820 16186
rect 25884 15978 25912 16662
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 26160 15706 26188 16050
rect 26238 16008 26294 16017
rect 26344 15994 26372 16934
rect 26436 16590 26464 17002
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26436 16046 26464 16526
rect 26294 15966 26372 15994
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 26238 15943 26294 15952
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26436 15570 26464 15982
rect 26528 15706 26556 17478
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 25780 15428 25832 15434
rect 25780 15370 25832 15376
rect 25778 15328 25834 15337
rect 25778 15263 25834 15272
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25596 15088 25648 15094
rect 25516 15048 25596 15076
rect 25516 14550 25544 15048
rect 25792 15042 25820 15263
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25596 15030 25648 15036
rect 25700 15014 25820 15042
rect 25594 14648 25650 14657
rect 25594 14583 25650 14592
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25516 13870 25544 14486
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25608 13025 25636 14583
rect 25594 13016 25650 13025
rect 25594 12951 25650 12960
rect 25412 12368 25464 12374
rect 25412 12310 25464 12316
rect 25700 12238 25728 15014
rect 26344 14346 26372 15438
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26436 14958 26464 15370
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14618 26464 14894
rect 26528 14618 26556 15302
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 25780 14272 25832 14278
rect 25778 14240 25780 14249
rect 25832 14240 25834 14249
rect 25778 14175 25834 14184
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 26056 14000 26108 14006
rect 26056 13942 26108 13948
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26068 13394 26096 13942
rect 26160 13530 26188 13942
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26068 13297 26096 13330
rect 26054 13288 26110 13297
rect 26528 13258 26556 14418
rect 26620 14346 26648 20742
rect 26974 20088 27030 20097
rect 26974 20023 27030 20032
rect 26988 19825 27016 20023
rect 26974 19816 27030 19825
rect 26974 19751 27030 19760
rect 26988 18970 27016 19751
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27356 19174 27384 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 26988 18358 27016 18906
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 26976 18352 27028 18358
rect 26976 18294 27028 18300
rect 27080 18222 27108 18838
rect 27356 18766 27384 19110
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 26896 17202 26924 17546
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 26698 16688 26754 16697
rect 26698 16623 26754 16632
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 26606 14104 26662 14113
rect 26712 14074 26740 16623
rect 26606 14039 26662 14048
rect 26700 14068 26752 14074
rect 26054 13223 26110 13232
rect 26516 13252 26568 13258
rect 26516 13194 26568 13200
rect 25778 13152 25834 13161
rect 25778 13087 25834 13096
rect 25792 12481 25820 13087
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 25778 12472 25834 12481
rect 25778 12407 25834 12416
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25424 11626 25452 12174
rect 25700 11898 25728 12174
rect 26436 12170 26464 12582
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26528 11898 26556 12242
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25424 11354 25452 11562
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 26160 11286 26188 11630
rect 26148 11280 26200 11286
rect 26148 11222 26200 11228
rect 26514 11248 26570 11257
rect 26514 11183 26570 11192
rect 26332 11076 26384 11082
rect 26332 11018 26384 11024
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25332 9178 25360 10678
rect 25962 10568 26018 10577
rect 25962 10503 25964 10512
rect 26016 10503 26018 10512
rect 25964 10474 26016 10480
rect 25870 10432 25926 10441
rect 25870 10367 25926 10376
rect 25410 10296 25466 10305
rect 25410 10231 25466 10240
rect 25424 9761 25452 10231
rect 25502 10024 25558 10033
rect 25502 9959 25558 9968
rect 25410 9752 25466 9761
rect 25410 9687 25466 9696
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25332 8634 25360 9114
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25424 7954 25452 9687
rect 25516 8634 25544 9959
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25778 8256 25834 8265
rect 25778 8191 25834 8200
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 25424 7546 25452 7890
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25792 3505 25820 8191
rect 25884 8090 25912 10367
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26344 9194 26372 11018
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26160 9166 26372 9194
rect 26160 9110 26188 9166
rect 26148 9104 26200 9110
rect 26148 9046 26200 9052
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 26344 5250 26372 7686
rect 26436 6458 26464 10474
rect 26528 10130 26556 11183
rect 26620 11014 26648 14039
rect 26700 14010 26752 14016
rect 26712 13870 26740 14010
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26698 12472 26754 12481
rect 26698 12407 26754 12416
rect 26712 11354 26740 12407
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26620 10606 26648 10950
rect 26712 10810 26740 11290
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26620 10266 26648 10542
rect 26608 10260 26660 10266
rect 26608 10202 26660 10208
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26528 9518 26556 10066
rect 26712 9722 26740 10746
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26516 9512 26568 9518
rect 26516 9454 26568 9460
rect 26514 9072 26570 9081
rect 26514 9007 26516 9016
rect 26568 9007 26570 9016
rect 26516 8978 26568 8984
rect 26528 8634 26556 8978
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26620 8401 26648 8502
rect 26606 8392 26662 8401
rect 26606 8327 26662 8336
rect 26712 8265 26740 8774
rect 26804 8566 26832 17070
rect 26896 16794 26924 17138
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26896 16425 26924 16594
rect 26974 16552 27030 16561
rect 26974 16487 27030 16496
rect 26882 16416 26938 16425
rect 26882 16351 26938 16360
rect 26988 15337 27016 16487
rect 26974 15328 27030 15337
rect 26974 15263 27030 15272
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26896 13530 26924 13670
rect 26884 13524 26936 13530
rect 26884 13466 26936 13472
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26988 12986 27016 13262
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 27080 12186 27108 18158
rect 27252 17808 27304 17814
rect 27252 17750 27304 17756
rect 27264 16998 27292 17750
rect 27436 17740 27488 17746
rect 27436 17682 27488 17688
rect 27448 16998 27476 17682
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 27436 16992 27488 16998
rect 27436 16934 27488 16940
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27172 16250 27200 16526
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27172 14074 27200 14350
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27160 13796 27212 13802
rect 27160 13738 27212 13744
rect 26896 12158 27108 12186
rect 26896 10305 26924 12158
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26988 11354 27016 12038
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 26976 11348 27028 11354
rect 26976 11290 27028 11296
rect 27080 11150 27108 11494
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27080 10674 27108 11086
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26882 10296 26938 10305
rect 27080 10266 27108 10610
rect 27172 10266 27200 13738
rect 27264 13274 27292 16934
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27356 13938 27384 14758
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27448 13433 27476 16934
rect 27540 16182 27568 17138
rect 27724 16998 27752 17614
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27528 16176 27580 16182
rect 27528 16118 27580 16124
rect 27620 15700 27672 15706
rect 27620 15642 27672 15648
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27540 15162 27568 15438
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27434 13424 27490 13433
rect 27434 13359 27490 13368
rect 27540 13326 27568 15098
rect 27632 14550 27660 15642
rect 27724 14822 27752 16934
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27620 14544 27672 14550
rect 27620 14486 27672 14492
rect 27816 14113 27844 17546
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 27802 14104 27858 14113
rect 28276 14074 28304 14554
rect 27802 14039 27858 14048
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 27632 13841 27660 13874
rect 27618 13832 27674 13841
rect 27618 13767 27674 13776
rect 27632 13530 27660 13767
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27528 13320 27580 13326
rect 27264 13246 27476 13274
rect 27528 13262 27580 13268
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27250 12608 27306 12617
rect 27250 12543 27306 12552
rect 26882 10231 26938 10240
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 27066 10160 27122 10169
rect 27066 10095 27122 10104
rect 26884 9920 26936 9926
rect 26884 9862 26936 9868
rect 26792 8560 26844 8566
rect 26792 8502 26844 8508
rect 26698 8256 26754 8265
rect 26698 8191 26754 8200
rect 26514 7848 26570 7857
rect 26514 7783 26570 7792
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26436 6254 26464 6394
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 26528 5778 26556 7783
rect 26792 7200 26844 7206
rect 26792 7142 26844 7148
rect 26606 6896 26662 6905
rect 26606 6831 26662 6840
rect 26620 6458 26648 6831
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26712 6361 26740 6598
rect 26698 6352 26754 6361
rect 26698 6287 26754 6296
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26528 5370 26556 5714
rect 26698 5672 26754 5681
rect 26698 5607 26700 5616
rect 26752 5607 26754 5616
rect 26700 5578 26752 5584
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 25884 5222 26372 5250
rect 26422 5264 26478 5273
rect 25778 3496 25834 3505
rect 25778 3431 25834 3440
rect 25884 1465 25912 5222
rect 26422 5199 26478 5208
rect 26332 5160 26384 5166
rect 26330 5128 26332 5137
rect 26384 5128 26386 5137
rect 26330 5063 26386 5072
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26436 2990 26464 5199
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26608 2848 26660 2854
rect 26606 2816 26608 2825
rect 26660 2816 26662 2825
rect 26606 2751 26662 2760
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 1456 25926 1465
rect 25870 1391 25926 1400
rect 1398 368 1454 377
rect 1398 303 1454 312
rect 4986 0 5042 480
rect 14922 0 14978 480
rect 24950 0 25006 480
rect 26804 377 26832 7142
rect 26896 921 26924 9862
rect 26976 9648 27028 9654
rect 26976 9590 27028 9596
rect 26988 2145 27016 9590
rect 27080 7342 27108 10095
rect 27264 7954 27292 12543
rect 27356 12442 27384 12922
rect 27344 12436 27396 12442
rect 27344 12378 27396 12384
rect 27252 7948 27304 7954
rect 27252 7890 27304 7896
rect 27264 7546 27292 7890
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27448 6866 27476 13246
rect 27540 12918 27568 13262
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27528 12776 27580 12782
rect 27526 12744 27528 12753
rect 27580 12744 27582 12753
rect 27526 12679 27582 12688
rect 27632 12238 27660 13466
rect 27804 12640 27856 12646
rect 27804 12582 27856 12588
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27632 10810 27660 11290
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27528 9512 27580 9518
rect 27526 9480 27528 9489
rect 27580 9480 27582 9489
rect 27526 9415 27582 9424
rect 27712 9376 27764 9382
rect 27710 9344 27712 9353
rect 27764 9344 27766 9353
rect 27710 9279 27766 9288
rect 27710 8664 27766 8673
rect 27710 8599 27712 8608
rect 27764 8599 27766 8608
rect 27712 8570 27764 8576
rect 27526 8528 27582 8537
rect 27526 8463 27582 8472
rect 27540 8430 27568 8463
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27712 7472 27764 7478
rect 27526 7440 27582 7449
rect 27526 7375 27582 7384
rect 27710 7440 27712 7449
rect 27764 7440 27766 7449
rect 27710 7375 27766 7384
rect 27540 7342 27568 7375
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 27448 6458 27476 6802
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27816 3913 27844 12582
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 28092 11898 28120 12174
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 27802 3904 27858 3913
rect 27802 3839 27858 3848
rect 26974 2136 27030 2145
rect 26974 2071 27030 2080
rect 26882 912 26938 921
rect 26882 847 26938 856
rect 26790 368 26846 377
rect 26790 303 26846 312
<< via2 >>
rect 3514 23568 3570 23624
rect 24950 23568 25006 23624
rect 3514 23024 3570 23080
rect 3238 22344 3294 22400
rect 3054 20576 3110 20632
rect 2502 20168 2558 20224
rect 2778 20168 2834 20224
rect 1950 19896 2006 19952
rect 1398 19760 1454 19816
rect 2410 19488 2466 19544
rect 2042 16632 2098 16688
rect 1950 15972 2006 16008
rect 1950 15952 1952 15972
rect 1952 15952 2004 15972
rect 2004 15952 2006 15972
rect 2042 15272 2098 15328
rect 1950 12960 2006 13016
rect 1950 12416 2006 12472
rect 1582 12300 1638 12336
rect 1582 12280 1584 12300
rect 1584 12280 1636 12300
rect 1636 12280 1638 12300
rect 1398 11736 1454 11792
rect 1950 9832 2006 9888
rect 1582 8084 1638 8120
rect 1582 8064 1584 8084
rect 1584 8064 1636 8084
rect 1636 8064 1638 8084
rect 1766 7792 1822 7848
rect 1582 7420 1584 7440
rect 1584 7420 1636 7440
rect 1636 7420 1638 7440
rect 1582 7384 1638 7420
rect 1582 6840 1638 6896
rect 1582 6332 1584 6352
rect 1584 6332 1636 6352
rect 1636 6332 1638 6352
rect 1582 6296 1638 6332
rect 2686 16496 2742 16552
rect 3146 15952 3202 16008
rect 4066 21800 4122 21856
rect 4434 21256 4490 21312
rect 3790 19896 3846 19952
rect 2686 15816 2742 15872
rect 2042 7404 2098 7440
rect 2042 7384 2044 7404
rect 2044 7384 2096 7404
rect 2096 7384 2098 7404
rect 3054 13776 3110 13832
rect 2962 13368 3018 13424
rect 3054 13232 3110 13288
rect 3238 15136 3294 15192
rect 3238 12824 3294 12880
rect 3422 12008 3478 12064
rect 3146 11736 3202 11792
rect 3238 11600 3294 11656
rect 2594 9288 2650 9344
rect 2686 8608 2742 8664
rect 2778 8336 2834 8392
rect 3606 12416 3662 12472
rect 3330 10124 3386 10160
rect 3330 10104 3332 10124
rect 3332 10104 3384 10124
rect 3384 10104 3386 10124
rect 3422 9968 3478 10024
rect 3606 7928 3662 7984
rect 3238 6316 3294 6352
rect 3238 6296 3240 6316
rect 3240 6296 3292 6316
rect 3292 6296 3294 6316
rect 1582 5636 1638 5672
rect 1582 5616 1584 5636
rect 1584 5616 1636 5636
rect 1636 5616 1638 5636
rect 1582 5072 1638 5128
rect 2042 5364 2098 5400
rect 2042 5344 2044 5364
rect 2044 5344 2096 5364
rect 2096 5344 2098 5364
rect 1490 3848 1546 3904
rect 2042 3440 2098 3496
rect 1582 2624 1638 2680
rect 3974 14592 4030 14648
rect 3974 13640 4030 13696
rect 4250 17584 4306 17640
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 4618 19488 4674 19544
rect 4618 13232 4674 13288
rect 4986 16360 5042 16416
rect 4802 12824 4858 12880
rect 4250 12280 4306 12336
rect 4434 12280 4490 12336
rect 4158 12144 4214 12200
rect 4066 11056 4122 11112
rect 3974 10376 4030 10432
rect 4066 9324 4068 9344
rect 4068 9324 4120 9344
rect 4120 9324 4122 9344
rect 4066 9288 4122 9324
rect 4434 10412 4436 10432
rect 4436 10412 4488 10432
rect 4488 10412 4490 10432
rect 4434 10376 4490 10412
rect 4066 9016 4122 9072
rect 4342 8372 4344 8392
rect 4344 8372 4396 8392
rect 4396 8372 4398 8392
rect 4342 8336 4398 8372
rect 3698 4392 3754 4448
rect 3790 3304 3846 3360
rect 2686 1400 2742 1456
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5630 15852 5632 15872
rect 5632 15852 5684 15872
rect 5684 15852 5686 15872
rect 5630 15816 5686 15852
rect 5538 15544 5594 15600
rect 5538 13948 5540 13968
rect 5540 13948 5592 13968
rect 5592 13948 5594 13968
rect 5538 13912 5594 13948
rect 5170 12552 5226 12608
rect 5630 12960 5686 13016
rect 5630 12688 5686 12744
rect 4986 11600 5042 11656
rect 5170 11464 5226 11520
rect 5538 11736 5594 11792
rect 5538 9560 5594 9616
rect 4618 5344 4674 5400
rect 5814 18128 5870 18184
rect 6550 18264 6606 18320
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5906 16668 5908 16688
rect 5908 16668 5960 16688
rect 5960 16668 5962 16688
rect 5906 16632 5962 16668
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 6642 17040 6698 17096
rect 6550 16360 6606 16416
rect 6642 16224 6698 16280
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 6274 11348 6330 11384
rect 6274 11328 6276 11348
rect 6276 11328 6328 11348
rect 6328 11328 6330 11348
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 6366 10784 6422 10840
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 7010 13640 7066 13696
rect 6274 9288 6330 9344
rect 5906 8880 5962 8936
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 5906 8472 5962 8528
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 9218 19488 9274 19544
rect 7930 17076 7932 17096
rect 7932 17076 7984 17096
rect 7984 17076 7986 17096
rect 7930 17040 7986 17076
rect 8298 17720 8354 17776
rect 8482 17720 8538 17776
rect 8022 16768 8078 16824
rect 8298 16088 8354 16144
rect 8574 15952 8630 16008
rect 8022 15000 8078 15056
rect 7654 14184 7710 14240
rect 8482 15136 8538 15192
rect 7470 11500 7472 11520
rect 7472 11500 7524 11520
rect 7524 11500 7526 11520
rect 7470 11464 7526 11500
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 7746 12688 7802 12744
rect 7746 12588 7748 12608
rect 7748 12588 7800 12608
rect 7800 12588 7802 12608
rect 7746 12552 7802 12588
rect 9218 14864 9274 14920
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10230 19896 10286 19952
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 10690 18708 10692 18728
rect 10692 18708 10744 18728
rect 10744 18708 10746 18728
rect 10690 18672 10746 18708
rect 11886 18808 11942 18864
rect 10322 17584 10378 17640
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10414 16788 10470 16824
rect 10414 16768 10416 16788
rect 10416 16768 10468 16788
rect 10468 16768 10470 16788
rect 8758 13776 8814 13832
rect 8574 12960 8630 13016
rect 7930 10548 7932 10568
rect 7932 10548 7984 10568
rect 7984 10548 7986 10568
rect 7930 10512 7986 10548
rect 8298 11736 8354 11792
rect 9310 12960 9366 13016
rect 9494 14476 9550 14512
rect 9494 14456 9496 14476
rect 9496 14456 9548 14476
rect 9548 14456 9550 14476
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10598 15444 10600 15464
rect 10600 15444 10652 15464
rect 10652 15444 10654 15464
rect 10598 15408 10654 15444
rect 10414 14320 10470 14376
rect 11150 15000 11206 15056
rect 11242 14884 11298 14920
rect 11242 14864 11244 14884
rect 11244 14864 11296 14884
rect 11296 14864 11298 14884
rect 9586 13368 9642 13424
rect 8850 12416 8906 12472
rect 7838 9324 7840 9344
rect 7840 9324 7892 9344
rect 7892 9324 7894 9344
rect 7838 9288 7894 9324
rect 7562 8472 7618 8528
rect 10046 12688 10102 12744
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10874 14184 10930 14240
rect 10874 13912 10930 13968
rect 10782 13232 10838 13288
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 12162 19488 12218 19544
rect 12070 16088 12126 16144
rect 11610 12824 11666 12880
rect 9678 11328 9734 11384
rect 11242 12144 11298 12200
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 9586 10376 9642 10432
rect 7378 8200 7434 8256
rect 9586 9968 9642 10024
rect 10414 11192 10470 11248
rect 6274 6296 6330 6352
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 7378 3440 7434 3496
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 11886 14048 11942 14104
rect 12438 19896 12494 19952
rect 14462 19352 14518 19408
rect 12438 18672 12494 18728
rect 12530 16496 12586 16552
rect 12254 15952 12310 16008
rect 12438 14456 12494 14512
rect 12438 13368 12494 13424
rect 12254 13096 12310 13152
rect 13358 18672 13414 18728
rect 13174 16940 13176 16960
rect 13176 16940 13228 16960
rect 13228 16940 13230 16960
rect 13174 16904 13230 16940
rect 13174 16496 13230 16552
rect 12622 15680 12678 15736
rect 12806 13640 12862 13696
rect 12806 12724 12808 12744
rect 12808 12724 12860 12744
rect 12860 12724 12862 12744
rect 12806 12688 12862 12724
rect 11702 10104 11758 10160
rect 13542 18028 13544 18048
rect 13544 18028 13596 18048
rect 13596 18028 13598 18048
rect 13542 17992 13598 18028
rect 13634 15680 13690 15736
rect 14370 16360 14426 16416
rect 14370 15952 14426 16008
rect 13266 13504 13322 13560
rect 13082 12280 13138 12336
rect 12990 9424 13046 9480
rect 10782 9324 10784 9344
rect 10784 9324 10836 9344
rect 10836 9324 10838 9344
rect 10782 9288 10838 9324
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10414 8200 10470 8256
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 13450 11056 13506 11112
rect 14002 14340 14058 14376
rect 14002 14320 14004 14340
rect 14004 14320 14056 14340
rect 14056 14320 14058 14340
rect 14002 13232 14058 13288
rect 14278 13232 14334 13288
rect 15014 18264 15070 18320
rect 15382 17992 15438 18048
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 16394 19216 16450 19272
rect 15658 18264 15714 18320
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 14738 16224 14794 16280
rect 14554 12960 14610 13016
rect 13634 10240 13690 10296
rect 14830 13812 14832 13832
rect 14832 13812 14884 13832
rect 14884 13812 14886 13832
rect 14830 13776 14886 13812
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15750 15156 15806 15192
rect 15750 15136 15752 15156
rect 15752 15136 15804 15156
rect 15804 15136 15806 15156
rect 15566 13796 15622 13832
rect 15566 13776 15568 13796
rect 15568 13776 15620 13796
rect 15620 13776 15622 13796
rect 15750 13912 15806 13968
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 16854 19236 16910 19272
rect 16854 19216 16856 19236
rect 16856 19216 16908 19236
rect 16908 19216 16910 19236
rect 16854 18264 16910 18320
rect 16762 17040 16818 17096
rect 17314 17584 17370 17640
rect 16486 16360 16542 16416
rect 17314 16632 17370 16688
rect 16670 14592 16726 14648
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 16762 14320 16818 14376
rect 16854 14048 16910 14104
rect 16394 13096 16450 13152
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15842 12416 15898 12472
rect 15474 10784 15530 10840
rect 14830 10648 14886 10704
rect 13450 9152 13506 9208
rect 13358 7928 13414 7984
rect 13266 7792 13322 7848
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 17038 13232 17094 13288
rect 16762 12316 16764 12336
rect 16764 12316 16816 12336
rect 16816 12316 16818 12336
rect 16762 12280 16818 12316
rect 16670 12144 16726 12200
rect 16302 11328 16358 11384
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 18050 19896 18106 19952
rect 18234 19352 18290 19408
rect 18234 17448 18290 17504
rect 17866 12708 17922 12744
rect 17866 12688 17868 12708
rect 17868 12688 17920 12708
rect 17920 12688 17922 12708
rect 18050 13912 18106 13968
rect 17406 10512 17462 10568
rect 16854 10412 16856 10432
rect 16856 10412 16908 10432
rect 16908 10412 16910 10432
rect 16854 10376 16910 10412
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 19430 19796 19432 19816
rect 19432 19796 19484 19816
rect 19484 19796 19486 19816
rect 19430 19760 19486 19796
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 20166 18672 20222 18728
rect 18602 16904 18658 16960
rect 18510 13640 18566 13696
rect 18418 12688 18474 12744
rect 18878 15544 18934 15600
rect 19430 16224 19486 16280
rect 20166 15000 20222 15056
rect 19706 14864 19762 14920
rect 19246 14220 19248 14240
rect 19248 14220 19300 14240
rect 19300 14220 19302 14240
rect 19246 14184 19302 14220
rect 18878 11872 18934 11928
rect 18602 11736 18658 11792
rect 18418 10648 18474 10704
rect 17774 9580 17830 9616
rect 17774 9560 17776 9580
rect 17776 9560 17828 9580
rect 17828 9560 17830 9580
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 18418 8472 18474 8528
rect 19062 13504 19118 13560
rect 19522 13812 19524 13832
rect 19524 13812 19576 13832
rect 19576 13812 19578 13832
rect 19522 13776 19578 13812
rect 20442 14592 20498 14648
rect 20258 14456 20314 14512
rect 19338 13232 19394 13288
rect 19246 11464 19302 11520
rect 19614 11872 19670 11928
rect 19614 10376 19670 10432
rect 20166 14320 20222 14376
rect 20074 14068 20130 14104
rect 20074 14048 20076 14068
rect 20076 14048 20128 14068
rect 20128 14048 20130 14068
rect 19890 13776 19946 13832
rect 20258 11348 20314 11384
rect 20258 11328 20260 11348
rect 20260 11328 20312 11348
rect 20312 11328 20314 11348
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 21362 17992 21418 18048
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 21362 15408 21418 15464
rect 21638 18164 21640 18184
rect 21640 18164 21692 18184
rect 21692 18164 21694 18184
rect 21638 18128 21694 18164
rect 22558 19216 22614 19272
rect 22466 19080 22522 19136
rect 21730 15680 21786 15736
rect 21914 14728 21970 14784
rect 20810 13640 20866 13696
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 21362 12860 21364 12880
rect 21364 12860 21416 12880
rect 21416 12860 21418 12880
rect 21362 12824 21418 12860
rect 21362 11736 21418 11792
rect 20810 11464 20866 11520
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 21454 11600 21510 11656
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20074 9832 20130 9888
rect 22006 13368 22062 13424
rect 22098 12960 22154 13016
rect 21822 12008 21878 12064
rect 21362 9460 21364 9480
rect 21364 9460 21416 9480
rect 21416 9460 21418 9480
rect 21362 9424 21418 9460
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 22098 11192 22154 11248
rect 23478 14864 23534 14920
rect 23754 15000 23810 15056
rect 23662 14320 23718 14376
rect 23478 13912 23534 13968
rect 23662 13796 23718 13832
rect 23662 13776 23664 13796
rect 23664 13776 23716 13796
rect 23716 13776 23718 13796
rect 22466 13096 22522 13152
rect 22374 12588 22376 12608
rect 22376 12588 22428 12608
rect 22428 12588 22430 12608
rect 22374 12552 22430 12588
rect 22006 8744 22062 8800
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 18970 7792 19026 7848
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 23478 11892 23534 11928
rect 23478 11872 23480 11892
rect 23480 11872 23532 11892
rect 23532 11872 23534 11892
rect 23754 12416 23810 12472
rect 23754 11756 23810 11792
rect 23754 11736 23756 11756
rect 23756 11736 23808 11756
rect 23808 11736 23810 11756
rect 25134 21256 25190 21312
rect 25318 23024 25374 23080
rect 25410 22344 25466 22400
rect 23938 17040 23994 17096
rect 24030 14728 24086 14784
rect 24122 14456 24178 14512
rect 24306 17992 24362 18048
rect 24030 12688 24086 12744
rect 24858 17992 24914 18048
rect 24674 16088 24730 16144
rect 24398 15544 24454 15600
rect 24674 15544 24730 15600
rect 25226 18944 25282 19000
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25502 21528 25558 21584
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25502 19216 25558 19272
rect 25410 18808 25466 18864
rect 25134 17720 25190 17776
rect 25042 16632 25098 16688
rect 24950 15816 25006 15872
rect 24582 15136 24638 15192
rect 24766 13796 24822 13832
rect 24766 13776 24768 13796
rect 24768 13776 24820 13796
rect 24820 13776 24822 13796
rect 24674 13232 24730 13288
rect 25042 15544 25098 15600
rect 24858 13096 24914 13152
rect 24214 10104 24270 10160
rect 24122 9832 24178 9888
rect 23938 8880 23994 8936
rect 26422 18944 26478 19000
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25686 17584 25742 17640
rect 25410 16088 25466 16144
rect 25226 14320 25282 14376
rect 25134 12824 25190 12880
rect 25042 12280 25098 12336
rect 25134 12144 25190 12200
rect 25042 11192 25098 11248
rect 24950 11056 25006 11112
rect 15842 7384 15898 7440
rect 22466 7384 22522 7440
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 14738 6160 14794 6216
rect 24766 6160 24822 6216
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 9678 5208 9734 5264
rect 24766 5072 24822 5128
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 24858 4528 24914 4584
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 4066 2080 4122 2136
rect 3974 856 4030 912
rect 7194 2352 7250 2408
rect 14922 2352 14978 2408
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 25778 17448 25834 17504
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25778 17040 25834 17096
rect 25778 16360 25834 16416
rect 25686 16224 25742 16280
rect 25594 15680 25650 15736
rect 25502 15136 25558 15192
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 26238 15952 26294 16008
rect 25778 15272 25834 15328
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25594 14592 25650 14648
rect 25594 12960 25650 13016
rect 25778 14220 25780 14240
rect 25780 14220 25832 14240
rect 25832 14220 25834 14240
rect 25778 14184 25834 14220
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 26054 13232 26110 13288
rect 26974 20032 27030 20088
rect 26974 19760 27030 19816
rect 26698 16632 26754 16688
rect 26606 14048 26662 14104
rect 25778 13096 25834 13152
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25778 12416 25834 12472
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26514 11192 26570 11248
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 25962 10532 26018 10568
rect 25962 10512 25964 10532
rect 25964 10512 26016 10532
rect 26016 10512 26018 10532
rect 25870 10376 25926 10432
rect 25410 10240 25466 10296
rect 25502 9968 25558 10024
rect 25410 9696 25466 9752
rect 25778 8200 25834 8256
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 26698 12416 26754 12472
rect 26514 9036 26570 9072
rect 26514 9016 26516 9036
rect 26516 9016 26568 9036
rect 26568 9016 26570 9036
rect 26606 8336 26662 8392
rect 26974 16496 27030 16552
rect 26882 16360 26938 16416
rect 26974 15272 27030 15328
rect 26882 10240 26938 10296
rect 27434 13368 27490 13424
rect 27802 14048 27858 14104
rect 27618 13776 27674 13832
rect 27250 12552 27306 12608
rect 27066 10104 27122 10160
rect 26698 8200 26754 8256
rect 26514 7792 26570 7848
rect 26606 6840 26662 6896
rect 26698 6296 26754 6352
rect 26698 5636 26754 5672
rect 26698 5616 26700 5636
rect 26700 5616 26752 5636
rect 26752 5616 26754 5636
rect 25778 3440 25834 3496
rect 26422 5208 26478 5264
rect 26330 5108 26332 5128
rect 26332 5108 26384 5128
rect 26384 5108 26386 5128
rect 26330 5072 26386 5108
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26606 5072 26662 5128
rect 26606 2796 26608 2816
rect 26608 2796 26660 2816
rect 26660 2796 26662 2816
rect 26606 2760 26662 2796
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 1400 25926 1456
rect 1398 312 1454 368
rect 27526 12724 27528 12744
rect 27528 12724 27580 12744
rect 27580 12724 27582 12744
rect 27526 12688 27582 12724
rect 27526 9460 27528 9480
rect 27528 9460 27580 9480
rect 27580 9460 27582 9480
rect 27526 9424 27582 9460
rect 27710 9324 27712 9344
rect 27712 9324 27764 9344
rect 27764 9324 27766 9344
rect 27710 9288 27766 9324
rect 27710 8628 27766 8664
rect 27710 8608 27712 8628
rect 27712 8608 27764 8628
rect 27764 8608 27766 8628
rect 27526 8472 27582 8528
rect 27526 7384 27582 7440
rect 27710 7420 27712 7440
rect 27712 7420 27764 7440
rect 27764 7420 27766 7440
rect 27710 7384 27766 7420
rect 27802 3848 27858 3904
rect 26974 2080 27030 2136
rect 26882 856 26938 912
rect 26790 312 26846 368
<< metal3 >>
rect 0 23626 480 23656
rect 3509 23626 3575 23629
rect 0 23624 3575 23626
rect 0 23568 3514 23624
rect 3570 23568 3575 23624
rect 0 23566 3575 23568
rect 0 23536 480 23566
rect 3509 23563 3575 23566
rect 24945 23626 25011 23629
rect 29520 23626 30000 23656
rect 24945 23624 30000 23626
rect 24945 23568 24950 23624
rect 25006 23568 30000 23624
rect 24945 23566 30000 23568
rect 24945 23563 25011 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3509 23082 3575 23085
rect 0 23080 3575 23082
rect 0 23024 3514 23080
rect 3570 23024 3575 23080
rect 0 23022 3575 23024
rect 0 22992 480 23022
rect 3509 23019 3575 23022
rect 25313 23082 25379 23085
rect 29520 23082 30000 23112
rect 25313 23080 30000 23082
rect 25313 23024 25318 23080
rect 25374 23024 30000 23080
rect 25313 23022 30000 23024
rect 25313 23019 25379 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 3233 22402 3299 22405
rect 0 22400 3299 22402
rect 0 22344 3238 22400
rect 3294 22344 3299 22400
rect 0 22342 3299 22344
rect 0 22312 480 22342
rect 3233 22339 3299 22342
rect 25405 22402 25471 22405
rect 29520 22402 30000 22432
rect 25405 22400 30000 22402
rect 25405 22344 25410 22400
rect 25466 22344 30000 22400
rect 25405 22342 30000 22344
rect 25405 22339 25471 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 4061 21858 4127 21861
rect 29520 21858 30000 21888
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 480 21798
rect 4061 21795 4127 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25497 21586 25563 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25497 21584 26434 21586
rect 25497 21528 25502 21584
rect 25558 21528 26434 21584
rect 25497 21526 26434 21528
rect 25497 21523 25563 21526
rect 0 21314 480 21344
rect 4429 21314 4495 21317
rect 0 21312 4495 21314
rect 0 21256 4434 21312
rect 4490 21256 4495 21312
rect 0 21254 4495 21256
rect 0 21224 480 21254
rect 4429 21251 4495 21254
rect 25129 21314 25195 21317
rect 29520 21314 30000 21344
rect 25129 21312 30000 21314
rect 25129 21256 25134 21312
rect 25190 21256 30000 21312
rect 25129 21254 30000 21256
rect 25129 21251 25195 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3049 20634 3115 20637
rect 29520 20634 30000 20664
rect 0 20632 3115 20634
rect 0 20576 3054 20632
rect 3110 20576 3115 20632
rect 0 20574 3115 20576
rect 0 20544 480 20574
rect 3049 20571 3115 20574
rect 26374 20574 30000 20634
rect 9622 20362 9628 20364
rect 7606 20302 9628 20362
rect 2497 20226 2563 20229
rect 2773 20226 2839 20229
rect 2497 20224 2839 20226
rect 2497 20168 2502 20224
rect 2558 20168 2778 20224
rect 2834 20168 2839 20224
rect 2497 20166 2839 20168
rect 2497 20163 2563 20166
rect 2773 20163 2839 20166
rect 0 20090 480 20120
rect 7606 20090 7666 20302
rect 9622 20300 9628 20302
rect 9692 20300 9698 20364
rect 10944 20160 11264 20161
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 0 20030 7666 20090
rect 0 20000 480 20030
rect 1945 19954 2011 19957
rect 3785 19954 3851 19957
rect 1945 19952 3851 19954
rect 1945 19896 1950 19952
rect 2006 19896 3790 19952
rect 3846 19896 3851 19952
rect 1945 19894 3851 19896
rect 1945 19891 2011 19894
rect 3785 19891 3851 19894
rect 10225 19954 10291 19957
rect 12433 19954 12499 19957
rect 10225 19952 12499 19954
rect 10225 19896 10230 19952
rect 10286 19896 12438 19952
rect 12494 19896 12499 19952
rect 10225 19894 12499 19896
rect 10225 19891 10291 19894
rect 12433 19891 12499 19894
rect 18045 19954 18111 19957
rect 26374 19954 26434 20574
rect 29520 20544 30000 20574
rect 26969 20090 27035 20093
rect 29520 20090 30000 20120
rect 26969 20088 30000 20090
rect 26969 20032 26974 20088
rect 27030 20032 30000 20088
rect 26969 20030 30000 20032
rect 26969 20027 27035 20030
rect 29520 20000 30000 20030
rect 18045 19952 26434 19954
rect 18045 19896 18050 19952
rect 18106 19896 26434 19952
rect 18045 19894 26434 19896
rect 18045 19891 18111 19894
rect 1393 19818 1459 19821
rect 19425 19818 19491 19821
rect 26969 19818 27035 19821
rect 1393 19816 27035 19818
rect 1393 19760 1398 19816
rect 1454 19760 19430 19816
rect 19486 19760 26974 19816
rect 27030 19760 27035 19816
rect 1393 19758 27035 19760
rect 1393 19755 1459 19758
rect 19425 19755 19491 19758
rect 26969 19755 27035 19758
rect 9622 19620 9628 19684
rect 9692 19682 9698 19684
rect 9692 19622 14658 19682
rect 9692 19620 9698 19622
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 2405 19546 2471 19549
rect 4613 19546 4679 19549
rect 2405 19544 4679 19546
rect 2405 19488 2410 19544
rect 2466 19488 4618 19544
rect 4674 19488 4679 19544
rect 2405 19486 4679 19488
rect 2405 19483 2471 19486
rect 4613 19483 4679 19486
rect 9213 19546 9279 19549
rect 12157 19546 12223 19549
rect 9213 19544 12223 19546
rect 9213 19488 9218 19544
rect 9274 19488 12162 19544
rect 12218 19488 12223 19544
rect 9213 19486 12223 19488
rect 9213 19483 9279 19486
rect 12157 19483 12223 19486
rect 0 19410 480 19440
rect 14457 19410 14523 19413
rect 0 19408 14523 19410
rect 0 19352 14462 19408
rect 14518 19352 14523 19408
rect 0 19350 14523 19352
rect 14598 19410 14658 19622
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 18229 19410 18295 19413
rect 29520 19410 30000 19440
rect 14598 19408 18295 19410
rect 14598 19352 18234 19408
rect 18290 19352 18295 19408
rect 14598 19350 18295 19352
rect 0 19320 480 19350
rect 14457 19347 14523 19350
rect 18229 19347 18295 19350
rect 24902 19350 30000 19410
rect 16389 19276 16455 19277
rect 16389 19274 16436 19276
rect 16344 19272 16436 19274
rect 16500 19274 16506 19276
rect 16849 19274 16915 19277
rect 22553 19274 22619 19277
rect 24902 19274 24962 19350
rect 29520 19320 30000 19350
rect 25497 19274 25563 19277
rect 16500 19272 24962 19274
rect 16344 19216 16394 19272
rect 16500 19216 16854 19272
rect 16910 19216 22558 19272
rect 22614 19216 24962 19272
rect 16344 19214 16436 19216
rect 16389 19212 16436 19214
rect 16500 19214 24962 19216
rect 25040 19272 25563 19274
rect 25040 19216 25502 19272
rect 25558 19216 25563 19272
rect 25040 19214 25563 19216
rect 16500 19212 16506 19214
rect 16389 19211 16455 19212
rect 16849 19211 16915 19214
rect 22553 19211 22619 19214
rect 22461 19138 22527 19141
rect 25040 19138 25100 19214
rect 25497 19211 25563 19214
rect 22461 19136 25100 19138
rect 22461 19080 22466 19136
rect 22522 19080 25100 19136
rect 22461 19078 25100 19080
rect 22461 19075 22527 19078
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 25221 19002 25287 19005
rect 26417 19002 26483 19005
rect 25221 19000 26483 19002
rect 25221 18944 25226 19000
rect 25282 18944 26422 19000
rect 26478 18944 26483 19000
rect 25221 18942 26483 18944
rect 25221 18939 25287 18942
rect 26417 18939 26483 18942
rect 0 18866 480 18896
rect 11881 18866 11947 18869
rect 0 18864 11947 18866
rect 0 18808 11886 18864
rect 11942 18808 11947 18864
rect 0 18806 11947 18808
rect 0 18776 480 18806
rect 11881 18803 11947 18806
rect 25405 18866 25471 18869
rect 29520 18866 30000 18896
rect 25405 18864 30000 18866
rect 25405 18808 25410 18864
rect 25466 18808 30000 18864
rect 25405 18806 30000 18808
rect 25405 18803 25471 18806
rect 29520 18776 30000 18806
rect 10685 18730 10751 18733
rect 12433 18730 12499 18733
rect 10685 18728 12499 18730
rect 10685 18672 10690 18728
rect 10746 18672 12438 18728
rect 12494 18672 12499 18728
rect 10685 18670 12499 18672
rect 10685 18667 10751 18670
rect 12433 18667 12499 18670
rect 13353 18730 13419 18733
rect 20161 18730 20227 18733
rect 13353 18728 20227 18730
rect 13353 18672 13358 18728
rect 13414 18672 20166 18728
rect 20222 18672 20227 18728
rect 13353 18670 20227 18672
rect 13353 18667 13419 18670
rect 20161 18667 20227 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 0 18322 480 18352
rect 6545 18322 6611 18325
rect 0 18320 6611 18322
rect 0 18264 6550 18320
rect 6606 18264 6611 18320
rect 0 18262 6611 18264
rect 0 18232 480 18262
rect 6545 18259 6611 18262
rect 15009 18322 15075 18325
rect 15653 18322 15719 18325
rect 16849 18322 16915 18325
rect 29520 18322 30000 18352
rect 15009 18320 16915 18322
rect 15009 18264 15014 18320
rect 15070 18264 15658 18320
rect 15714 18264 16854 18320
rect 16910 18264 16915 18320
rect 15009 18262 16915 18264
rect 15009 18259 15075 18262
rect 15653 18259 15719 18262
rect 16849 18259 16915 18262
rect 25822 18262 30000 18322
rect 5809 18186 5875 18189
rect 21633 18186 21699 18189
rect 5809 18184 21699 18186
rect 5809 18128 5814 18184
rect 5870 18128 21638 18184
rect 21694 18128 21699 18184
rect 5809 18126 21699 18128
rect 5809 18123 5875 18126
rect 21633 18123 21699 18126
rect 13537 18050 13603 18053
rect 15377 18050 15443 18053
rect 13537 18048 15443 18050
rect 13537 17992 13542 18048
rect 13598 17992 15382 18048
rect 15438 17992 15443 18048
rect 13537 17990 15443 17992
rect 13537 17987 13603 17990
rect 15377 17987 15443 17990
rect 21357 18050 21423 18053
rect 24301 18050 24367 18053
rect 24853 18050 24919 18053
rect 21357 18048 24919 18050
rect 21357 17992 21362 18048
rect 21418 17992 24306 18048
rect 24362 17992 24858 18048
rect 24914 17992 24919 18048
rect 21357 17990 24919 17992
rect 21357 17987 21423 17990
rect 24301 17987 24367 17990
rect 24853 17987 24919 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 8293 17778 8359 17781
rect 614 17776 8359 17778
rect 614 17720 8298 17776
rect 8354 17720 8359 17776
rect 614 17718 8359 17720
rect 0 17642 480 17672
rect 614 17642 674 17718
rect 8293 17715 8359 17718
rect 8477 17778 8543 17781
rect 25129 17778 25195 17781
rect 25822 17778 25882 18262
rect 29520 18232 30000 18262
rect 8477 17776 25882 17778
rect 8477 17720 8482 17776
rect 8538 17720 25134 17776
rect 25190 17720 25882 17776
rect 8477 17718 25882 17720
rect 8477 17715 8543 17718
rect 25129 17715 25195 17718
rect 0 17582 674 17642
rect 4245 17642 4311 17645
rect 10317 17642 10383 17645
rect 17309 17642 17375 17645
rect 4245 17640 17375 17642
rect 4245 17584 4250 17640
rect 4306 17584 10322 17640
rect 10378 17584 17314 17640
rect 17370 17584 17375 17640
rect 4245 17582 17375 17584
rect 0 17552 480 17582
rect 4245 17579 4311 17582
rect 10317 17579 10383 17582
rect 17309 17579 17375 17582
rect 25681 17642 25747 17645
rect 29520 17642 30000 17672
rect 25681 17640 30000 17642
rect 25681 17584 25686 17640
rect 25742 17584 30000 17640
rect 25681 17582 30000 17584
rect 25681 17579 25747 17582
rect 29520 17552 30000 17582
rect 18229 17506 18295 17509
rect 25773 17506 25839 17509
rect 18229 17504 25839 17506
rect 18229 17448 18234 17504
rect 18290 17448 25778 17504
rect 25834 17448 25839 17504
rect 18229 17446 25839 17448
rect 18229 17443 18295 17446
rect 25773 17443 25839 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 0 17098 480 17128
rect 6637 17098 6703 17101
rect 0 17096 6703 17098
rect 0 17040 6642 17096
rect 6698 17040 6703 17096
rect 0 17038 6703 17040
rect 0 17008 480 17038
rect 6637 17035 6703 17038
rect 7925 17098 7991 17101
rect 16757 17098 16823 17101
rect 23933 17098 23999 17101
rect 7925 17096 23999 17098
rect 7925 17040 7930 17096
rect 7986 17040 16762 17096
rect 16818 17040 23938 17096
rect 23994 17040 23999 17096
rect 7925 17038 23999 17040
rect 7925 17035 7991 17038
rect 16757 17035 16823 17038
rect 23933 17035 23999 17038
rect 25773 17098 25839 17101
rect 29520 17098 30000 17128
rect 25773 17096 30000 17098
rect 25773 17040 25778 17096
rect 25834 17040 30000 17096
rect 25773 17038 30000 17040
rect 25773 17035 25839 17038
rect 29520 17008 30000 17038
rect 13169 16962 13235 16965
rect 18597 16962 18663 16965
rect 13169 16960 18663 16962
rect 13169 16904 13174 16960
rect 13230 16904 18602 16960
rect 18658 16904 18663 16960
rect 13169 16902 18663 16904
rect 13169 16899 13235 16902
rect 18597 16899 18663 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 8017 16826 8083 16829
rect 10409 16826 10475 16829
rect 8017 16824 10475 16826
rect 8017 16768 8022 16824
rect 8078 16768 10414 16824
rect 10470 16768 10475 16824
rect 8017 16766 10475 16768
rect 8017 16763 8083 16766
rect 10409 16763 10475 16766
rect 2037 16690 2103 16693
rect 5901 16690 5967 16693
rect 2037 16688 5967 16690
rect 2037 16632 2042 16688
rect 2098 16632 5906 16688
rect 5962 16632 5967 16688
rect 2037 16630 5967 16632
rect 2037 16627 2103 16630
rect 5901 16627 5967 16630
rect 17309 16690 17375 16693
rect 25037 16690 25103 16693
rect 26693 16690 26759 16693
rect 17309 16688 26759 16690
rect 17309 16632 17314 16688
rect 17370 16632 25042 16688
rect 25098 16632 26698 16688
rect 26754 16632 26759 16688
rect 17309 16630 26759 16632
rect 17309 16627 17375 16630
rect 25037 16627 25103 16630
rect 26693 16627 26759 16630
rect 2681 16554 2747 16557
rect 12525 16554 12591 16557
rect 2681 16552 12591 16554
rect 2681 16496 2686 16552
rect 2742 16496 12530 16552
rect 12586 16496 12591 16552
rect 2681 16494 12591 16496
rect 2681 16491 2747 16494
rect 12525 16491 12591 16494
rect 13169 16554 13235 16557
rect 26969 16554 27035 16557
rect 13169 16552 27035 16554
rect 13169 16496 13174 16552
rect 13230 16496 26974 16552
rect 27030 16496 27035 16552
rect 13169 16494 27035 16496
rect 13169 16491 13235 16494
rect 26969 16491 27035 16494
rect 0 16418 480 16448
rect 4981 16418 5047 16421
rect 0 16416 5047 16418
rect 0 16360 4986 16416
rect 5042 16360 5047 16416
rect 0 16358 5047 16360
rect 0 16328 480 16358
rect 4981 16355 5047 16358
rect 6545 16418 6611 16421
rect 14365 16418 14431 16421
rect 6545 16416 14431 16418
rect 6545 16360 6550 16416
rect 6606 16360 14370 16416
rect 14426 16360 14431 16416
rect 6545 16358 14431 16360
rect 6545 16355 6611 16358
rect 14365 16355 14431 16358
rect 16481 16418 16547 16421
rect 25773 16418 25839 16421
rect 16481 16416 25839 16418
rect 16481 16360 16486 16416
rect 16542 16360 25778 16416
rect 25834 16360 25839 16416
rect 16481 16358 25839 16360
rect 16481 16355 16547 16358
rect 25773 16355 25839 16358
rect 26877 16418 26943 16421
rect 29520 16418 30000 16448
rect 26877 16416 30000 16418
rect 26877 16360 26882 16416
rect 26938 16360 30000 16416
rect 26877 16358 30000 16360
rect 26877 16355 26943 16358
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 29520 16328 30000 16358
rect 25944 16287 26264 16288
rect 6637 16282 6703 16285
rect 14733 16282 14799 16285
rect 6637 16280 14799 16282
rect 6637 16224 6642 16280
rect 6698 16224 14738 16280
rect 14794 16224 14799 16280
rect 6637 16222 14799 16224
rect 6637 16219 6703 16222
rect 14733 16219 14799 16222
rect 19425 16282 19491 16285
rect 25681 16282 25747 16285
rect 19425 16280 25747 16282
rect 19425 16224 19430 16280
rect 19486 16224 25686 16280
rect 25742 16224 25747 16280
rect 19425 16222 25747 16224
rect 19425 16219 19491 16222
rect 25681 16219 25747 16222
rect 8293 16146 8359 16149
rect 12065 16146 12131 16149
rect 8293 16144 12131 16146
rect 8293 16088 8298 16144
rect 8354 16088 12070 16144
rect 12126 16088 12131 16144
rect 8293 16086 12131 16088
rect 8293 16083 8359 16086
rect 12065 16083 12131 16086
rect 24669 16146 24735 16149
rect 25405 16146 25471 16149
rect 24669 16144 25471 16146
rect 24669 16088 24674 16144
rect 24730 16088 25410 16144
rect 25466 16088 25471 16144
rect 24669 16086 25471 16088
rect 24669 16083 24735 16086
rect 25405 16083 25471 16086
rect 1945 16010 2011 16013
rect 3141 16010 3207 16013
rect 8569 16010 8635 16013
rect 12249 16010 12315 16013
rect 1945 16008 8635 16010
rect 1945 15952 1950 16008
rect 2006 15952 3146 16008
rect 3202 15952 8574 16008
rect 8630 15952 8635 16008
rect 1945 15950 8635 15952
rect 1945 15947 2011 15950
rect 3141 15947 3207 15950
rect 8569 15947 8635 15950
rect 10734 16008 12315 16010
rect 10734 15952 12254 16008
rect 12310 15952 12315 16008
rect 10734 15950 12315 15952
rect 0 15874 480 15904
rect 2681 15874 2747 15877
rect 0 15872 2747 15874
rect 0 15816 2686 15872
rect 2742 15816 2747 15872
rect 0 15814 2747 15816
rect 0 15784 480 15814
rect 2681 15811 2747 15814
rect 5625 15874 5691 15877
rect 10734 15874 10794 15950
rect 12249 15947 12315 15950
rect 14365 16010 14431 16013
rect 26233 16010 26299 16013
rect 14365 16008 26299 16010
rect 14365 15952 14370 16008
rect 14426 15952 26238 16008
rect 26294 15952 26299 16008
rect 14365 15950 26299 15952
rect 14365 15947 14431 15950
rect 26233 15947 26299 15950
rect 5625 15872 10794 15874
rect 5625 15816 5630 15872
rect 5686 15816 10794 15872
rect 5625 15814 10794 15816
rect 24945 15874 25011 15877
rect 29520 15874 30000 15904
rect 24945 15872 30000 15874
rect 24945 15816 24950 15872
rect 25006 15816 30000 15872
rect 24945 15814 30000 15816
rect 5625 15811 5691 15814
rect 24945 15811 25011 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 12617 15738 12683 15741
rect 13629 15738 13695 15741
rect 21725 15738 21791 15741
rect 25589 15738 25655 15741
rect 12617 15736 19074 15738
rect 12617 15680 12622 15736
rect 12678 15680 13634 15736
rect 13690 15680 19074 15736
rect 12617 15678 19074 15680
rect 12617 15675 12683 15678
rect 13629 15675 13695 15678
rect 5533 15602 5599 15605
rect 18873 15602 18939 15605
rect 5533 15600 18939 15602
rect 5533 15544 5538 15600
rect 5594 15544 18878 15600
rect 18934 15544 18939 15600
rect 5533 15542 18939 15544
rect 19014 15602 19074 15678
rect 21725 15736 25655 15738
rect 21725 15680 21730 15736
rect 21786 15680 25594 15736
rect 25650 15680 25655 15736
rect 21725 15678 25655 15680
rect 21725 15675 21791 15678
rect 25589 15675 25655 15678
rect 24393 15602 24459 15605
rect 24669 15602 24735 15605
rect 19014 15600 24735 15602
rect 19014 15544 24398 15600
rect 24454 15544 24674 15600
rect 24730 15544 24735 15600
rect 19014 15542 24735 15544
rect 5533 15539 5599 15542
rect 18873 15539 18939 15542
rect 24393 15539 24459 15542
rect 24669 15539 24735 15542
rect 25037 15600 25103 15605
rect 25037 15544 25042 15600
rect 25098 15544 25103 15600
rect 25037 15539 25103 15544
rect 10593 15466 10659 15469
rect 21357 15466 21423 15469
rect 10593 15464 21423 15466
rect 10593 15408 10598 15464
rect 10654 15408 21362 15464
rect 21418 15408 21423 15464
rect 10593 15406 21423 15408
rect 10593 15403 10659 15406
rect 21357 15403 21423 15406
rect 0 15330 480 15360
rect 2037 15330 2103 15333
rect 0 15328 2103 15330
rect 0 15272 2042 15328
rect 2098 15272 2103 15328
rect 0 15270 2103 15272
rect 25040 15330 25100 15539
rect 25773 15330 25839 15333
rect 25040 15328 25839 15330
rect 25040 15272 25778 15328
rect 25834 15272 25839 15328
rect 25040 15270 25839 15272
rect 0 15240 480 15270
rect 2037 15267 2103 15270
rect 25773 15267 25839 15270
rect 26969 15330 27035 15333
rect 29520 15330 30000 15360
rect 26969 15328 30000 15330
rect 26969 15272 26974 15328
rect 27030 15272 30000 15328
rect 26969 15270 30000 15272
rect 26969 15267 27035 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 3233 15194 3299 15197
rect 3366 15194 3372 15196
rect 3233 15192 3372 15194
rect 3233 15136 3238 15192
rect 3294 15136 3372 15192
rect 3233 15134 3372 15136
rect 3233 15131 3299 15134
rect 3366 15132 3372 15134
rect 3436 15132 3442 15196
rect 8477 15194 8543 15197
rect 15745 15194 15811 15197
rect 8477 15192 15811 15194
rect 8477 15136 8482 15192
rect 8538 15136 15750 15192
rect 15806 15136 15811 15192
rect 8477 15134 15811 15136
rect 8477 15131 8543 15134
rect 15745 15131 15811 15134
rect 24577 15194 24643 15197
rect 25497 15194 25563 15197
rect 24577 15192 25563 15194
rect 24577 15136 24582 15192
rect 24638 15136 25502 15192
rect 25558 15136 25563 15192
rect 24577 15134 25563 15136
rect 24577 15131 24643 15134
rect 25497 15131 25563 15134
rect 8017 15058 8083 15061
rect 11145 15058 11211 15061
rect 8017 15056 11211 15058
rect 8017 15000 8022 15056
rect 8078 15000 11150 15056
rect 11206 15000 11211 15056
rect 8017 14998 11211 15000
rect 8017 14995 8083 14998
rect 11145 14995 11211 14998
rect 20161 15058 20227 15061
rect 23749 15058 23815 15061
rect 20161 15056 23815 15058
rect 20161 15000 20166 15056
rect 20222 15000 23754 15056
rect 23810 15000 23815 15056
rect 20161 14998 23815 15000
rect 20161 14995 20227 14998
rect 23749 14995 23815 14998
rect 9213 14922 9279 14925
rect 11237 14922 11303 14925
rect 9213 14920 11303 14922
rect 9213 14864 9218 14920
rect 9274 14864 11242 14920
rect 11298 14864 11303 14920
rect 9213 14862 11303 14864
rect 9213 14859 9279 14862
rect 11237 14859 11303 14862
rect 19701 14922 19767 14925
rect 23473 14922 23539 14925
rect 19701 14920 23539 14922
rect 19701 14864 19706 14920
rect 19762 14864 23478 14920
rect 23534 14864 23539 14920
rect 19701 14862 23539 14864
rect 19701 14859 19767 14862
rect 23473 14859 23539 14862
rect 21909 14786 21975 14789
rect 24025 14786 24091 14789
rect 21909 14784 24091 14786
rect 21909 14728 21914 14784
rect 21970 14728 24030 14784
rect 24086 14728 24091 14784
rect 21909 14726 24091 14728
rect 21909 14723 21975 14726
rect 24025 14723 24091 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 3969 14650 4035 14653
rect 0 14648 4035 14650
rect 0 14592 3974 14648
rect 4030 14592 4035 14648
rect 0 14590 4035 14592
rect 0 14560 480 14590
rect 3969 14587 4035 14590
rect 16665 14650 16731 14653
rect 20437 14650 20503 14653
rect 16665 14648 20503 14650
rect 16665 14592 16670 14648
rect 16726 14592 20442 14648
rect 20498 14592 20503 14648
rect 16665 14590 20503 14592
rect 16665 14587 16731 14590
rect 20437 14587 20503 14590
rect 25589 14650 25655 14653
rect 29520 14650 30000 14680
rect 25589 14648 30000 14650
rect 25589 14592 25594 14648
rect 25650 14592 30000 14648
rect 25589 14590 30000 14592
rect 25589 14587 25655 14590
rect 29520 14560 30000 14590
rect 9489 14514 9555 14517
rect 12433 14514 12499 14517
rect 9489 14512 12499 14514
rect 9489 14456 9494 14512
rect 9550 14456 12438 14512
rect 12494 14456 12499 14512
rect 9489 14454 12499 14456
rect 9489 14451 9555 14454
rect 12433 14451 12499 14454
rect 20253 14514 20319 14517
rect 24117 14514 24183 14517
rect 20253 14512 24183 14514
rect 20253 14456 20258 14512
rect 20314 14456 24122 14512
rect 24178 14456 24183 14512
rect 20253 14454 24183 14456
rect 20253 14451 20319 14454
rect 24117 14451 24183 14454
rect 10409 14378 10475 14381
rect 13997 14378 14063 14381
rect 10409 14376 14063 14378
rect 10409 14320 10414 14376
rect 10470 14320 14002 14376
rect 14058 14320 14063 14376
rect 10409 14318 14063 14320
rect 10409 14315 10475 14318
rect 13997 14315 14063 14318
rect 16757 14378 16823 14381
rect 20161 14378 20227 14381
rect 16757 14376 20227 14378
rect 16757 14320 16762 14376
rect 16818 14320 20166 14376
rect 20222 14320 20227 14376
rect 16757 14318 20227 14320
rect 16757 14315 16823 14318
rect 20161 14315 20227 14318
rect 23657 14378 23723 14381
rect 25221 14378 25287 14381
rect 23657 14376 25287 14378
rect 23657 14320 23662 14376
rect 23718 14320 25226 14376
rect 25282 14320 25287 14376
rect 23657 14318 25287 14320
rect 23657 14315 23723 14318
rect 25221 14315 25287 14318
rect 7649 14242 7715 14245
rect 10869 14242 10935 14245
rect 7649 14240 10935 14242
rect 7649 14184 7654 14240
rect 7710 14184 10874 14240
rect 10930 14184 10935 14240
rect 7649 14182 10935 14184
rect 7649 14179 7715 14182
rect 10869 14179 10935 14182
rect 19241 14242 19307 14245
rect 25773 14242 25839 14245
rect 19241 14240 25839 14242
rect 19241 14184 19246 14240
rect 19302 14184 25778 14240
rect 25834 14184 25839 14240
rect 19241 14182 25839 14184
rect 19241 14179 19307 14182
rect 25773 14179 25839 14182
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 11881 14106 11947 14109
rect 0 14046 3066 14106
rect 0 14016 480 14046
rect 3006 13837 3066 14046
rect 10734 14104 11947 14106
rect 10734 14048 11886 14104
rect 11942 14048 11947 14104
rect 10734 14046 11947 14048
rect 5533 13970 5599 13973
rect 10734 13970 10794 14046
rect 11881 14043 11947 14046
rect 16849 14106 16915 14109
rect 20069 14106 20135 14109
rect 16849 14104 20135 14106
rect 16849 14048 16854 14104
rect 16910 14048 20074 14104
rect 20130 14048 20135 14104
rect 16849 14046 20135 14048
rect 16849 14043 16915 14046
rect 20069 14043 20135 14046
rect 26601 14106 26667 14109
rect 27797 14106 27863 14109
rect 29520 14106 30000 14136
rect 26601 14104 30000 14106
rect 26601 14048 26606 14104
rect 26662 14048 27802 14104
rect 27858 14048 30000 14104
rect 26601 14046 30000 14048
rect 26601 14043 26667 14046
rect 27797 14043 27863 14046
rect 29520 14016 30000 14046
rect 5533 13968 10794 13970
rect 5533 13912 5538 13968
rect 5594 13912 10794 13968
rect 5533 13910 10794 13912
rect 10869 13970 10935 13973
rect 15745 13970 15811 13973
rect 10869 13968 15811 13970
rect 10869 13912 10874 13968
rect 10930 13912 15750 13968
rect 15806 13912 15811 13968
rect 10869 13910 15811 13912
rect 5533 13907 5599 13910
rect 10869 13907 10935 13910
rect 15745 13907 15811 13910
rect 17902 13908 17908 13972
rect 17972 13970 17978 13972
rect 18045 13970 18111 13973
rect 23473 13970 23539 13973
rect 17972 13968 23539 13970
rect 17972 13912 18050 13968
rect 18106 13912 23478 13968
rect 23534 13912 23539 13968
rect 17972 13910 23539 13912
rect 17972 13908 17978 13910
rect 18045 13907 18111 13910
rect 23473 13907 23539 13910
rect 3006 13832 3115 13837
rect 3006 13776 3054 13832
rect 3110 13776 3115 13832
rect 3006 13774 3115 13776
rect 3049 13771 3115 13774
rect 8753 13834 8819 13837
rect 14825 13834 14891 13837
rect 8753 13832 14891 13834
rect 8753 13776 8758 13832
rect 8814 13776 14830 13832
rect 14886 13776 14891 13832
rect 8753 13774 14891 13776
rect 8753 13771 8819 13774
rect 14825 13771 14891 13774
rect 15561 13834 15627 13837
rect 19517 13834 19583 13837
rect 19885 13834 19951 13837
rect 23657 13834 23723 13837
rect 15561 13832 19810 13834
rect 15561 13776 15566 13832
rect 15622 13776 19522 13832
rect 19578 13776 19810 13832
rect 15561 13774 19810 13776
rect 15561 13771 15627 13774
rect 19517 13771 19583 13774
rect 3969 13698 4035 13701
rect 7005 13698 7071 13701
rect 3969 13696 7071 13698
rect 3969 13640 3974 13696
rect 4030 13640 7010 13696
rect 7066 13640 7071 13696
rect 3969 13638 7071 13640
rect 3969 13635 4035 13638
rect 7005 13635 7071 13638
rect 12801 13698 12867 13701
rect 18505 13698 18571 13701
rect 12801 13696 18571 13698
rect 12801 13640 12806 13696
rect 12862 13640 18510 13696
rect 18566 13640 18571 13696
rect 12801 13638 18571 13640
rect 19750 13698 19810 13774
rect 19885 13832 23723 13834
rect 19885 13776 19890 13832
rect 19946 13776 23662 13832
rect 23718 13776 23723 13832
rect 19885 13774 23723 13776
rect 19885 13771 19951 13774
rect 23657 13771 23723 13774
rect 24761 13834 24827 13837
rect 27613 13834 27679 13837
rect 24761 13832 27679 13834
rect 24761 13776 24766 13832
rect 24822 13776 27618 13832
rect 27674 13776 27679 13832
rect 24761 13774 27679 13776
rect 24761 13771 24827 13774
rect 27613 13771 27679 13774
rect 20805 13698 20871 13701
rect 19750 13696 20871 13698
rect 19750 13640 20810 13696
rect 20866 13640 20871 13696
rect 19750 13638 20871 13640
rect 12801 13635 12867 13638
rect 18505 13635 18571 13638
rect 20805 13635 20871 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 13261 13562 13327 13565
rect 19057 13562 19123 13565
rect 13261 13560 19123 13562
rect 13261 13504 13266 13560
rect 13322 13504 19062 13560
rect 19118 13504 19123 13560
rect 13261 13502 19123 13504
rect 13261 13499 13327 13502
rect 19057 13499 19123 13502
rect 0 13426 480 13456
rect 2957 13426 3023 13429
rect 0 13424 3023 13426
rect 0 13368 2962 13424
rect 3018 13368 3023 13424
rect 0 13366 3023 13368
rect 0 13336 480 13366
rect 2957 13363 3023 13366
rect 9581 13426 9647 13429
rect 12433 13426 12499 13429
rect 9581 13424 12499 13426
rect 9581 13368 9586 13424
rect 9642 13368 12438 13424
rect 12494 13368 12499 13424
rect 9581 13366 12499 13368
rect 9581 13363 9647 13366
rect 12433 13363 12499 13366
rect 22001 13426 22067 13429
rect 27429 13426 27495 13429
rect 29520 13426 30000 13456
rect 22001 13424 30000 13426
rect 22001 13368 22006 13424
rect 22062 13368 27434 13424
rect 27490 13368 30000 13424
rect 22001 13366 30000 13368
rect 22001 13363 22067 13366
rect 27429 13363 27495 13366
rect 29520 13336 30000 13366
rect 3049 13290 3115 13293
rect 4613 13290 4679 13293
rect 10777 13290 10843 13293
rect 13997 13290 14063 13293
rect 3049 13288 6424 13290
rect 3049 13232 3054 13288
rect 3110 13232 4618 13288
rect 4674 13232 6424 13288
rect 3049 13230 6424 13232
rect 3049 13227 3115 13230
rect 4613 13227 4679 13230
rect 6364 13154 6424 13230
rect 10777 13288 14063 13290
rect 10777 13232 10782 13288
rect 10838 13232 14002 13288
rect 14058 13232 14063 13288
rect 10777 13230 14063 13232
rect 10777 13227 10843 13230
rect 13997 13227 14063 13230
rect 14273 13290 14339 13293
rect 17033 13290 17099 13293
rect 19333 13290 19399 13293
rect 24669 13290 24735 13293
rect 26049 13290 26115 13293
rect 14273 13288 24594 13290
rect 14273 13232 14278 13288
rect 14334 13232 17038 13288
rect 17094 13232 19338 13288
rect 19394 13232 24594 13288
rect 14273 13230 24594 13232
rect 14273 13227 14339 13230
rect 17033 13227 17099 13230
rect 19333 13227 19399 13230
rect 12249 13154 12315 13157
rect 6364 13152 12315 13154
rect 6364 13096 12254 13152
rect 12310 13096 12315 13152
rect 6364 13094 12315 13096
rect 12249 13091 12315 13094
rect 16389 13154 16455 13157
rect 22461 13154 22527 13157
rect 16389 13152 22527 13154
rect 16389 13096 16394 13152
rect 16450 13096 22466 13152
rect 22522 13096 22527 13152
rect 16389 13094 22527 13096
rect 24534 13154 24594 13230
rect 24669 13288 26115 13290
rect 24669 13232 24674 13288
rect 24730 13232 26054 13288
rect 26110 13232 26115 13288
rect 24669 13230 26115 13232
rect 24669 13227 24735 13230
rect 26049 13227 26115 13230
rect 24853 13154 24919 13157
rect 25773 13154 25839 13157
rect 24534 13152 25839 13154
rect 24534 13096 24858 13152
rect 24914 13096 25778 13152
rect 25834 13096 25839 13152
rect 24534 13094 25839 13096
rect 16389 13091 16455 13094
rect 22461 13091 22527 13094
rect 24853 13091 24919 13094
rect 25773 13091 25839 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 1945 13018 2011 13021
rect 5625 13018 5691 13021
rect 1945 13016 5691 13018
rect 1945 12960 1950 13016
rect 2006 12960 5630 13016
rect 5686 12960 5691 13016
rect 1945 12958 5691 12960
rect 1945 12955 2011 12958
rect 5625 12955 5691 12958
rect 8569 13018 8635 13021
rect 9305 13018 9371 13021
rect 14549 13018 14615 13021
rect 22093 13018 22159 13021
rect 25589 13018 25655 13021
rect 8569 13016 15762 13018
rect 8569 12960 8574 13016
rect 8630 12960 9310 13016
rect 9366 12960 14554 13016
rect 14610 12960 15762 13016
rect 8569 12958 15762 12960
rect 8569 12955 8635 12958
rect 9305 12955 9371 12958
rect 14549 12955 14615 12958
rect 0 12882 480 12912
rect 3233 12882 3299 12885
rect 4797 12882 4863 12885
rect 11605 12882 11671 12885
rect 0 12880 11671 12882
rect 0 12824 3238 12880
rect 3294 12824 4802 12880
rect 4858 12824 11610 12880
rect 11666 12824 11671 12880
rect 0 12822 11671 12824
rect 15702 12882 15762 12958
rect 22093 13016 25655 13018
rect 22093 12960 22098 13016
rect 22154 12960 25594 13016
rect 25650 12960 25655 13016
rect 22093 12958 25655 12960
rect 22093 12955 22159 12958
rect 25589 12955 25655 12958
rect 21357 12882 21423 12885
rect 15702 12880 21423 12882
rect 15702 12824 21362 12880
rect 21418 12824 21423 12880
rect 15702 12822 21423 12824
rect 0 12792 480 12822
rect 3233 12819 3299 12822
rect 4797 12819 4863 12822
rect 11605 12819 11671 12822
rect 21357 12819 21423 12822
rect 25129 12882 25195 12885
rect 29520 12882 30000 12912
rect 25129 12880 30000 12882
rect 25129 12824 25134 12880
rect 25190 12824 30000 12880
rect 25129 12822 30000 12824
rect 25129 12819 25195 12822
rect 29520 12792 30000 12822
rect 5625 12746 5691 12749
rect 7741 12746 7807 12749
rect 10041 12746 10107 12749
rect 5625 12744 10107 12746
rect 5625 12688 5630 12744
rect 5686 12688 7746 12744
rect 7802 12688 10046 12744
rect 10102 12688 10107 12744
rect 5625 12686 10107 12688
rect 5625 12683 5691 12686
rect 7741 12683 7807 12686
rect 10041 12683 10107 12686
rect 12801 12746 12867 12749
rect 17861 12746 17927 12749
rect 12801 12744 17927 12746
rect 12801 12688 12806 12744
rect 12862 12688 17866 12744
rect 17922 12688 17927 12744
rect 12801 12686 17927 12688
rect 12801 12683 12867 12686
rect 17861 12683 17927 12686
rect 18413 12746 18479 12749
rect 24025 12746 24091 12749
rect 27521 12746 27587 12749
rect 18413 12744 27587 12746
rect 18413 12688 18418 12744
rect 18474 12688 24030 12744
rect 24086 12688 27526 12744
rect 27582 12688 27587 12744
rect 18413 12686 27587 12688
rect 18413 12683 18479 12686
rect 24025 12683 24091 12686
rect 27521 12683 27587 12686
rect 5165 12610 5231 12613
rect 7741 12610 7807 12613
rect 5165 12608 7807 12610
rect 5165 12552 5170 12608
rect 5226 12552 7746 12608
rect 7802 12552 7807 12608
rect 5165 12550 7807 12552
rect 5165 12547 5231 12550
rect 7741 12547 7807 12550
rect 22369 12610 22435 12613
rect 27245 12610 27311 12613
rect 22369 12608 27311 12610
rect 22369 12552 22374 12608
rect 22430 12552 27250 12608
rect 27306 12552 27311 12608
rect 22369 12550 27311 12552
rect 22369 12547 22435 12550
rect 27245 12547 27311 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 1945 12474 2011 12477
rect 1350 12472 2011 12474
rect 1350 12416 1950 12472
rect 2006 12416 2011 12472
rect 1350 12414 2011 12416
rect 0 12338 480 12368
rect 1350 12338 1410 12414
rect 1945 12411 2011 12414
rect 3601 12474 3667 12477
rect 8845 12474 8911 12477
rect 3601 12472 8911 12474
rect 3601 12416 3606 12472
rect 3662 12416 8850 12472
rect 8906 12416 8911 12472
rect 3601 12414 8911 12416
rect 3601 12411 3667 12414
rect 8845 12411 8911 12414
rect 15837 12474 15903 12477
rect 16430 12474 16436 12476
rect 15837 12472 16436 12474
rect 15837 12416 15842 12472
rect 15898 12416 16436 12472
rect 15837 12414 16436 12416
rect 15837 12411 15903 12414
rect 16430 12412 16436 12414
rect 16500 12412 16506 12476
rect 23749 12474 23815 12477
rect 25773 12474 25839 12477
rect 26693 12474 26759 12477
rect 23749 12472 25330 12474
rect 23749 12416 23754 12472
rect 23810 12416 25330 12472
rect 23749 12414 25330 12416
rect 23749 12411 23815 12414
rect 0 12278 1410 12338
rect 1577 12338 1643 12341
rect 4245 12338 4311 12341
rect 1577 12336 4311 12338
rect 1577 12280 1582 12336
rect 1638 12280 4250 12336
rect 4306 12280 4311 12336
rect 1577 12278 4311 12280
rect 0 12248 480 12278
rect 1577 12275 1643 12278
rect 4245 12275 4311 12278
rect 4429 12338 4495 12341
rect 13077 12338 13143 12341
rect 4429 12336 13143 12338
rect 4429 12280 4434 12336
rect 4490 12280 13082 12336
rect 13138 12280 13143 12336
rect 4429 12278 13143 12280
rect 4429 12275 4495 12278
rect 13077 12275 13143 12278
rect 16757 12338 16823 12341
rect 25037 12338 25103 12341
rect 16757 12336 25103 12338
rect 16757 12280 16762 12336
rect 16818 12280 25042 12336
rect 25098 12280 25103 12336
rect 16757 12278 25103 12280
rect 25270 12338 25330 12414
rect 25773 12472 26759 12474
rect 25773 12416 25778 12472
rect 25834 12416 26698 12472
rect 26754 12416 26759 12472
rect 25773 12414 26759 12416
rect 25773 12411 25839 12414
rect 26693 12411 26759 12414
rect 29520 12338 30000 12368
rect 25270 12278 30000 12338
rect 16757 12275 16823 12278
rect 25037 12275 25103 12278
rect 29520 12248 30000 12278
rect 4153 12202 4219 12205
rect 11237 12202 11303 12205
rect 4153 12200 11303 12202
rect 4153 12144 4158 12200
rect 4214 12144 11242 12200
rect 11298 12144 11303 12200
rect 4153 12142 11303 12144
rect 4153 12139 4219 12142
rect 11237 12139 11303 12142
rect 16665 12202 16731 12205
rect 25129 12202 25195 12205
rect 16665 12200 25195 12202
rect 16665 12144 16670 12200
rect 16726 12144 25134 12200
rect 25190 12144 25195 12200
rect 16665 12142 25195 12144
rect 16665 12139 16731 12142
rect 25129 12139 25195 12142
rect 3417 12066 3483 12069
rect 3734 12066 3740 12068
rect 3417 12064 3740 12066
rect 3417 12008 3422 12064
rect 3478 12008 3740 12064
rect 3417 12006 3740 12008
rect 3417 12003 3483 12006
rect 3734 12004 3740 12006
rect 3804 12004 3810 12068
rect 21817 12066 21883 12069
rect 18462 12064 21883 12066
rect 18462 12008 21822 12064
rect 21878 12008 21883 12064
rect 18462 12006 21883 12008
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 1393 11794 1459 11797
rect 3141 11794 3207 11797
rect 1393 11792 3207 11794
rect 1393 11736 1398 11792
rect 1454 11736 3146 11792
rect 3202 11736 3207 11792
rect 1393 11734 3207 11736
rect 1393 11731 1459 11734
rect 3141 11731 3207 11734
rect 5533 11794 5599 11797
rect 8293 11794 8359 11797
rect 5533 11792 8359 11794
rect 5533 11736 5538 11792
rect 5594 11736 8298 11792
rect 8354 11736 8359 11792
rect 5533 11734 8359 11736
rect 5533 11731 5599 11734
rect 8293 11731 8359 11734
rect 0 11658 480 11688
rect 3233 11658 3299 11661
rect 0 11656 3299 11658
rect 0 11600 3238 11656
rect 3294 11600 3299 11656
rect 0 11598 3299 11600
rect 0 11568 480 11598
rect 3233 11595 3299 11598
rect 4981 11658 5047 11661
rect 18462 11658 18522 12006
rect 21817 12003 21883 12006
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 18873 11930 18939 11933
rect 19609 11930 19675 11933
rect 23473 11930 23539 11933
rect 18873 11928 23539 11930
rect 18873 11872 18878 11928
rect 18934 11872 19614 11928
rect 19670 11872 23478 11928
rect 23534 11872 23539 11928
rect 18873 11870 23539 11872
rect 18873 11867 18939 11870
rect 19609 11867 19675 11870
rect 23473 11867 23539 11870
rect 18597 11794 18663 11797
rect 21357 11794 21423 11797
rect 23749 11794 23815 11797
rect 18597 11792 23815 11794
rect 18597 11736 18602 11792
rect 18658 11736 21362 11792
rect 21418 11736 23754 11792
rect 23810 11736 23815 11792
rect 18597 11734 23815 11736
rect 18597 11731 18663 11734
rect 21357 11731 21423 11734
rect 23749 11731 23815 11734
rect 4981 11656 18522 11658
rect 4981 11600 4986 11656
rect 5042 11600 18522 11656
rect 4981 11598 18522 11600
rect 21449 11658 21515 11661
rect 29520 11658 30000 11688
rect 21449 11656 30000 11658
rect 21449 11600 21454 11656
rect 21510 11600 30000 11656
rect 21449 11598 30000 11600
rect 4981 11595 5047 11598
rect 21449 11595 21515 11598
rect 29520 11568 30000 11598
rect 5165 11522 5231 11525
rect 7465 11522 7531 11525
rect 5165 11520 7531 11522
rect 5165 11464 5170 11520
rect 5226 11464 7470 11520
rect 7526 11464 7531 11520
rect 5165 11462 7531 11464
rect 5165 11459 5231 11462
rect 7465 11459 7531 11462
rect 19241 11522 19307 11525
rect 20805 11522 20871 11525
rect 19241 11520 20871 11522
rect 19241 11464 19246 11520
rect 19302 11464 20810 11520
rect 20866 11464 20871 11520
rect 19241 11462 20871 11464
rect 19241 11459 19307 11462
rect 20805 11459 20871 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 6269 11386 6335 11389
rect 9673 11386 9739 11389
rect 6269 11384 9739 11386
rect 6269 11328 6274 11384
rect 6330 11328 9678 11384
rect 9734 11328 9739 11384
rect 6269 11326 9739 11328
rect 6269 11323 6335 11326
rect 9673 11323 9739 11326
rect 16297 11386 16363 11389
rect 20253 11386 20319 11389
rect 16297 11384 20319 11386
rect 16297 11328 16302 11384
rect 16358 11328 20258 11384
rect 20314 11328 20319 11384
rect 16297 11326 20319 11328
rect 16297 11323 16363 11326
rect 20253 11323 20319 11326
rect 10409 11250 10475 11253
rect 22093 11250 22159 11253
rect 10409 11248 22159 11250
rect 10409 11192 10414 11248
rect 10470 11192 22098 11248
rect 22154 11192 22159 11248
rect 10409 11190 22159 11192
rect 10409 11187 10475 11190
rect 22093 11187 22159 11190
rect 25037 11250 25103 11253
rect 26509 11250 26575 11253
rect 25037 11248 26575 11250
rect 25037 11192 25042 11248
rect 25098 11192 26514 11248
rect 26570 11192 26575 11248
rect 25037 11190 26575 11192
rect 25037 11187 25103 11190
rect 26509 11187 26575 11190
rect 0 11114 480 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 0 11024 480 11054
rect 4061 11051 4127 11054
rect 13302 11052 13308 11116
rect 13372 11114 13378 11116
rect 13445 11114 13511 11117
rect 13372 11112 13511 11114
rect 13372 11056 13450 11112
rect 13506 11056 13511 11112
rect 13372 11054 13511 11056
rect 13372 11052 13378 11054
rect 13445 11051 13511 11054
rect 24945 11114 25011 11117
rect 29520 11114 30000 11144
rect 24945 11112 30000 11114
rect 24945 11056 24950 11112
rect 25006 11056 30000 11112
rect 24945 11054 30000 11056
rect 24945 11051 25011 11054
rect 29520 11024 30000 11054
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 6361 10842 6427 10845
rect 15469 10842 15535 10845
rect 6361 10840 15535 10842
rect 6361 10784 6366 10840
rect 6422 10784 15474 10840
rect 15530 10784 15535 10840
rect 6361 10782 15535 10784
rect 6361 10779 6427 10782
rect 15469 10779 15535 10782
rect 14825 10706 14891 10709
rect 18413 10706 18479 10709
rect 14825 10704 18479 10706
rect 14825 10648 14830 10704
rect 14886 10648 18418 10704
rect 18474 10648 18479 10704
rect 14825 10646 18479 10648
rect 14825 10643 14891 10646
rect 18413 10643 18479 10646
rect 7925 10570 7991 10573
rect 17401 10570 17467 10573
rect 25957 10570 26023 10573
rect 7925 10568 17467 10570
rect 7925 10512 7930 10568
rect 7986 10512 17406 10568
rect 17462 10512 17467 10568
rect 7925 10510 17467 10512
rect 7925 10507 7991 10510
rect 17401 10507 17467 10510
rect 19750 10568 26023 10570
rect 19750 10512 25962 10568
rect 26018 10512 26023 10568
rect 19750 10510 26023 10512
rect 0 10434 480 10464
rect 3969 10434 4035 10437
rect 0 10432 4035 10434
rect 0 10376 3974 10432
rect 4030 10376 4035 10432
rect 0 10374 4035 10376
rect 0 10344 480 10374
rect 3969 10371 4035 10374
rect 4429 10434 4495 10437
rect 9581 10434 9647 10437
rect 4429 10432 9647 10434
rect 4429 10376 4434 10432
rect 4490 10376 9586 10432
rect 9642 10376 9647 10432
rect 4429 10374 9647 10376
rect 4429 10371 4495 10374
rect 9581 10371 9647 10374
rect 16849 10434 16915 10437
rect 19609 10434 19675 10437
rect 16849 10432 19675 10434
rect 16849 10376 16854 10432
rect 16910 10376 19614 10432
rect 19670 10376 19675 10432
rect 16849 10374 19675 10376
rect 16849 10371 16915 10374
rect 19609 10371 19675 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 13629 10298 13695 10301
rect 11470 10296 13695 10298
rect 11470 10240 13634 10296
rect 13690 10240 13695 10296
rect 11470 10238 13695 10240
rect 3325 10162 3391 10165
rect 11470 10162 11530 10238
rect 13629 10235 13695 10238
rect 11697 10162 11763 10165
rect 19750 10162 19810 10510
rect 25957 10507 26023 10510
rect 25865 10434 25931 10437
rect 29520 10434 30000 10464
rect 25865 10432 30000 10434
rect 25865 10376 25870 10432
rect 25926 10376 30000 10432
rect 25865 10374 30000 10376
rect 25865 10371 25931 10374
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 25405 10298 25471 10301
rect 26877 10298 26943 10301
rect 25405 10296 26943 10298
rect 25405 10240 25410 10296
rect 25466 10240 26882 10296
rect 26938 10240 26943 10296
rect 25405 10238 26943 10240
rect 25405 10235 25471 10238
rect 26877 10235 26943 10238
rect 3325 10160 11530 10162
rect 3325 10104 3330 10160
rect 3386 10104 11530 10160
rect 3325 10102 11530 10104
rect 11654 10160 19810 10162
rect 11654 10104 11702 10160
rect 11758 10104 19810 10160
rect 11654 10102 19810 10104
rect 24209 10162 24275 10165
rect 27061 10162 27127 10165
rect 24209 10160 27127 10162
rect 24209 10104 24214 10160
rect 24270 10104 27066 10160
rect 27122 10104 27127 10160
rect 24209 10102 27127 10104
rect 3325 10099 3391 10102
rect 11654 10099 11763 10102
rect 24209 10099 24275 10102
rect 27061 10099 27127 10102
rect 3417 10026 3483 10029
rect 9581 10026 9647 10029
rect 11654 10026 11714 10099
rect 25497 10026 25563 10029
rect 3417 10024 6562 10026
rect 3417 9968 3422 10024
rect 3478 9968 6562 10024
rect 3417 9966 6562 9968
rect 3417 9963 3483 9966
rect 0 9890 480 9920
rect 1945 9890 2011 9893
rect 0 9888 2011 9890
rect 0 9832 1950 9888
rect 2006 9832 2011 9888
rect 0 9830 2011 9832
rect 0 9800 480 9830
rect 1945 9827 2011 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 6502 9754 6562 9966
rect 9581 10024 11714 10026
rect 9581 9968 9586 10024
rect 9642 9968 11714 10024
rect 9581 9966 11714 9968
rect 14552 9966 16452 10026
rect 9581 9963 9647 9966
rect 14552 9754 14612 9966
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 6502 9694 14612 9754
rect 16392 9754 16452 9966
rect 25497 10024 26434 10026
rect 25497 9968 25502 10024
rect 25558 9968 26434 10024
rect 25497 9966 26434 9968
rect 25497 9963 25563 9966
rect 20069 9890 20135 9893
rect 24117 9890 24183 9893
rect 20069 9888 24183 9890
rect 20069 9832 20074 9888
rect 20130 9832 24122 9888
rect 24178 9832 24183 9888
rect 20069 9830 24183 9832
rect 26374 9890 26434 9966
rect 29520 9890 30000 9920
rect 26374 9830 30000 9890
rect 20069 9827 20135 9830
rect 24117 9827 24183 9830
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 25405 9754 25471 9757
rect 16392 9752 25471 9754
rect 16392 9696 25410 9752
rect 25466 9696 25471 9752
rect 16392 9694 25471 9696
rect 25405 9691 25471 9694
rect 5533 9618 5599 9621
rect 17769 9618 17835 9621
rect 5533 9616 17835 9618
rect 5533 9560 5538 9616
rect 5594 9560 17774 9616
rect 17830 9560 17835 9616
rect 5533 9558 17835 9560
rect 5533 9555 5599 9558
rect 17769 9555 17835 9558
rect 12985 9482 13051 9485
rect 21357 9482 21423 9485
rect 27521 9482 27587 9485
rect 12985 9480 27587 9482
rect 12985 9424 12990 9480
rect 13046 9424 21362 9480
rect 21418 9424 27526 9480
rect 27582 9424 27587 9480
rect 12985 9422 27587 9424
rect 12985 9419 13051 9422
rect 21357 9419 21423 9422
rect 27521 9419 27587 9422
rect 0 9346 480 9376
rect 2589 9346 2655 9349
rect 0 9344 2655 9346
rect 0 9288 2594 9344
rect 2650 9288 2655 9344
rect 0 9286 2655 9288
rect 0 9256 480 9286
rect 2589 9283 2655 9286
rect 4061 9346 4127 9349
rect 6269 9346 6335 9349
rect 4061 9344 6335 9346
rect 4061 9288 4066 9344
rect 4122 9288 6274 9344
rect 6330 9288 6335 9344
rect 4061 9286 6335 9288
rect 4061 9283 4127 9286
rect 6269 9283 6335 9286
rect 7833 9346 7899 9349
rect 10777 9346 10843 9349
rect 7833 9344 10843 9346
rect 7833 9288 7838 9344
rect 7894 9288 10782 9344
rect 10838 9288 10843 9344
rect 7833 9286 10843 9288
rect 7833 9283 7899 9286
rect 10777 9283 10843 9286
rect 27705 9346 27771 9349
rect 29520 9346 30000 9376
rect 27705 9344 30000 9346
rect 27705 9288 27710 9344
rect 27766 9288 30000 9344
rect 27705 9286 30000 9288
rect 27705 9283 27771 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 13445 9210 13511 9213
rect 13445 9208 17418 9210
rect 13445 9152 13450 9208
rect 13506 9152 17418 9208
rect 13445 9150 17418 9152
rect 13445 9147 13511 9150
rect 4061 9074 4127 9077
rect 17358 9074 17418 9150
rect 26509 9074 26575 9077
rect 4061 9072 17234 9074
rect 4061 9016 4066 9072
rect 4122 9016 17234 9072
rect 4061 9014 17234 9016
rect 17358 9072 26575 9074
rect 17358 9016 26514 9072
rect 26570 9016 26575 9072
rect 17358 9014 26575 9016
rect 4061 9011 4127 9014
rect 5901 8938 5967 8941
rect 17174 8938 17234 9014
rect 26509 9011 26575 9014
rect 23933 8938 23999 8941
rect 5901 8936 17050 8938
rect 5901 8880 5906 8936
rect 5962 8880 17050 8936
rect 5901 8878 17050 8880
rect 17174 8936 23999 8938
rect 17174 8880 23938 8936
rect 23994 8880 23999 8936
rect 17174 8878 23999 8880
rect 5901 8875 5967 8878
rect 16990 8802 17050 8878
rect 23933 8875 23999 8878
rect 22001 8802 22067 8805
rect 16990 8800 22067 8802
rect 16990 8744 22006 8800
rect 22062 8744 22067 8800
rect 16990 8742 22067 8744
rect 22001 8739 22067 8742
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 2681 8666 2747 8669
rect 0 8664 2747 8666
rect 0 8608 2686 8664
rect 2742 8608 2747 8664
rect 0 8606 2747 8608
rect 0 8576 480 8606
rect 2681 8603 2747 8606
rect 27705 8666 27771 8669
rect 29520 8666 30000 8696
rect 27705 8664 30000 8666
rect 27705 8608 27710 8664
rect 27766 8608 30000 8664
rect 27705 8606 30000 8608
rect 27705 8603 27771 8606
rect 29520 8576 30000 8606
rect 5901 8530 5967 8533
rect 7557 8530 7623 8533
rect 5901 8528 7623 8530
rect 5901 8472 5906 8528
rect 5962 8472 7562 8528
rect 7618 8472 7623 8528
rect 5901 8470 7623 8472
rect 5901 8467 5967 8470
rect 7557 8467 7623 8470
rect 18413 8530 18479 8533
rect 27521 8530 27587 8533
rect 18413 8528 27587 8530
rect 18413 8472 18418 8528
rect 18474 8472 27526 8528
rect 27582 8472 27587 8528
rect 18413 8470 27587 8472
rect 18413 8467 18479 8470
rect 27521 8467 27587 8470
rect 2773 8394 2839 8397
rect 4337 8394 4403 8397
rect 2773 8392 4403 8394
rect 2773 8336 2778 8392
rect 2834 8336 4342 8392
rect 4398 8336 4403 8392
rect 2773 8334 4403 8336
rect 2773 8331 2839 8334
rect 4337 8331 4403 8334
rect 26601 8394 26667 8397
rect 26601 8392 27584 8394
rect 26601 8336 26606 8392
rect 26662 8336 27584 8392
rect 26601 8334 27584 8336
rect 26601 8331 26667 8334
rect 7373 8258 7439 8261
rect 10409 8258 10475 8261
rect 7373 8256 10475 8258
rect 7373 8200 7378 8256
rect 7434 8200 10414 8256
rect 10470 8200 10475 8256
rect 7373 8198 10475 8200
rect 7373 8195 7439 8198
rect 10409 8195 10475 8198
rect 25773 8258 25839 8261
rect 26693 8258 26759 8261
rect 25773 8256 26759 8258
rect 25773 8200 25778 8256
rect 25834 8200 26698 8256
rect 26754 8200 26759 8256
rect 25773 8198 26759 8200
rect 25773 8195 25839 8198
rect 26693 8195 26759 8198
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 27524 8122 27584 8334
rect 29520 8122 30000 8152
rect 27524 8062 30000 8122
rect 0 8032 480 8062
rect 1577 8059 1643 8062
rect 29520 8032 30000 8062
rect 3601 7986 3667 7989
rect 13353 7986 13419 7989
rect 3601 7984 13419 7986
rect 3601 7928 3606 7984
rect 3662 7928 13358 7984
rect 13414 7928 13419 7984
rect 3601 7926 13419 7928
rect 3601 7923 3667 7926
rect 13353 7923 13419 7926
rect 1761 7850 1827 7853
rect 13261 7850 13327 7853
rect 1761 7848 13327 7850
rect 1761 7792 1766 7848
rect 1822 7792 13266 7848
rect 13322 7792 13327 7848
rect 1761 7790 13327 7792
rect 1761 7787 1827 7790
rect 13261 7787 13327 7790
rect 18965 7850 19031 7853
rect 26509 7850 26575 7853
rect 18965 7848 26575 7850
rect 18965 7792 18970 7848
rect 19026 7792 26514 7848
rect 26570 7792 26575 7848
rect 18965 7790 26575 7792
rect 18965 7787 19031 7790
rect 26509 7787 26575 7790
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 2037 7442 2103 7445
rect 15837 7442 15903 7445
rect 2037 7440 15903 7442
rect 2037 7384 2042 7440
rect 2098 7384 15842 7440
rect 15898 7384 15903 7440
rect 2037 7382 15903 7384
rect 2037 7379 2103 7382
rect 15837 7379 15903 7382
rect 22461 7442 22527 7445
rect 27521 7442 27587 7445
rect 22461 7440 27587 7442
rect 22461 7384 22466 7440
rect 22522 7384 27526 7440
rect 27582 7384 27587 7440
rect 22461 7382 27587 7384
rect 22461 7379 22527 7382
rect 27521 7379 27587 7382
rect 27705 7442 27771 7445
rect 29520 7442 30000 7472
rect 27705 7440 30000 7442
rect 27705 7384 27710 7440
rect 27766 7384 30000 7440
rect 27705 7382 30000 7384
rect 27705 7379 27771 7382
rect 29520 7352 30000 7382
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 26601 6898 26667 6901
rect 29520 6898 30000 6928
rect 26601 6896 30000 6898
rect 26601 6840 26606 6896
rect 26662 6840 30000 6896
rect 26601 6838 30000 6840
rect 26601 6835 26667 6838
rect 29520 6808 30000 6838
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 3233 6354 3299 6357
rect 6269 6354 6335 6357
rect 3233 6352 6335 6354
rect 3233 6296 3238 6352
rect 3294 6296 6274 6352
rect 6330 6296 6335 6352
rect 3233 6294 6335 6296
rect 3233 6291 3299 6294
rect 6269 6291 6335 6294
rect 26693 6354 26759 6357
rect 29520 6354 30000 6384
rect 26693 6352 30000 6354
rect 26693 6296 26698 6352
rect 26754 6296 30000 6352
rect 26693 6294 30000 6296
rect 26693 6291 26759 6294
rect 29520 6264 30000 6294
rect 14733 6218 14799 6221
rect 24761 6218 24827 6221
rect 14733 6216 24827 6218
rect 14733 6160 14738 6216
rect 14794 6160 24766 6216
rect 24822 6160 24827 6216
rect 14733 6158 24827 6160
rect 14733 6155 14799 6158
rect 24761 6155 24827 6158
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 26693 5674 26759 5677
rect 29520 5674 30000 5704
rect 26693 5672 30000 5674
rect 26693 5616 26698 5672
rect 26754 5616 30000 5672
rect 26693 5614 30000 5616
rect 26693 5611 26759 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 2037 5402 2103 5405
rect 4613 5402 4679 5405
rect 2037 5400 4679 5402
rect 2037 5344 2042 5400
rect 2098 5344 4618 5400
rect 4674 5344 4679 5400
rect 2037 5342 4679 5344
rect 2037 5339 2103 5342
rect 4613 5339 4679 5342
rect 9673 5266 9739 5269
rect 26417 5266 26483 5269
rect 9673 5264 26483 5266
rect 9673 5208 9678 5264
rect 9734 5208 26422 5264
rect 26478 5208 26483 5264
rect 9673 5206 26483 5208
rect 9673 5203 9739 5206
rect 26417 5203 26483 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 24761 5130 24827 5133
rect 26325 5130 26391 5133
rect 24761 5128 26391 5130
rect 24761 5072 24766 5128
rect 24822 5072 26330 5128
rect 26386 5072 26391 5128
rect 24761 5070 26391 5072
rect 24761 5067 24827 5070
rect 26325 5067 26391 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 24853 4586 24919 4589
rect 24853 4584 26434 4586
rect 24853 4528 24858 4584
rect 24914 4528 26434 4584
rect 24853 4526 26434 4528
rect 24853 4523 24919 4526
rect 0 4450 480 4480
rect 3693 4450 3759 4453
rect 0 4448 3759 4450
rect 0 4392 3698 4448
rect 3754 4392 3759 4448
rect 0 4390 3759 4392
rect 26374 4450 26434 4526
rect 29520 4450 30000 4480
rect 26374 4390 30000 4450
rect 0 4360 480 4390
rect 3693 4387 3759 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 0 3906 480 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 480 3846
rect 1485 3843 1551 3846
rect 27797 3906 27863 3909
rect 29520 3906 30000 3936
rect 27797 3904 30000 3906
rect 27797 3848 27802 3904
rect 27858 3848 30000 3904
rect 27797 3846 30000 3848
rect 27797 3843 27863 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 2037 3498 2103 3501
rect 7373 3498 7439 3501
rect 2037 3496 7439 3498
rect 2037 3440 2042 3496
rect 2098 3440 7378 3496
rect 7434 3440 7439 3496
rect 2037 3438 7439 3440
rect 2037 3435 2103 3438
rect 7373 3435 7439 3438
rect 25773 3498 25839 3501
rect 25773 3496 26434 3498
rect 25773 3440 25778 3496
rect 25834 3440 26434 3496
rect 25773 3438 26434 3440
rect 25773 3435 25839 3438
rect 0 3362 480 3392
rect 3785 3362 3851 3365
rect 0 3360 3851 3362
rect 0 3304 3790 3360
rect 3846 3304 3851 3360
rect 0 3302 3851 3304
rect 26374 3362 26434 3438
rect 29520 3362 30000 3392
rect 26374 3302 30000 3362
rect 0 3272 480 3302
rect 3785 3299 3851 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 26601 2818 26667 2821
rect 26601 2816 26802 2818
rect 26601 2760 26606 2816
rect 26662 2760 26802 2816
rect 26601 2758 26802 2760
rect 26601 2755 26667 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 26742 2682 26802 2758
rect 29520 2682 30000 2712
rect 26742 2622 30000 2682
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 29520 2592 30000 2622
rect 7189 2410 7255 2413
rect 14917 2410 14983 2413
rect 7189 2408 14983 2410
rect 7189 2352 7194 2408
rect 7250 2352 14922 2408
rect 14978 2352 14983 2408
rect 7189 2350 14983 2352
rect 7189 2347 7255 2350
rect 14917 2347 14983 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 4061 2138 4127 2141
rect 0 2136 4127 2138
rect 0 2080 4066 2136
rect 4122 2080 4127 2136
rect 0 2078 4127 2080
rect 0 2048 480 2078
rect 4061 2075 4127 2078
rect 26969 2138 27035 2141
rect 29520 2138 30000 2168
rect 26969 2136 30000 2138
rect 26969 2080 26974 2136
rect 27030 2080 30000 2136
rect 26969 2078 30000 2080
rect 26969 2075 27035 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 2681 1458 2747 1461
rect 0 1456 2747 1458
rect 0 1400 2686 1456
rect 2742 1400 2747 1456
rect 0 1398 2747 1400
rect 0 1368 480 1398
rect 2681 1395 2747 1398
rect 25865 1458 25931 1461
rect 29520 1458 30000 1488
rect 25865 1456 30000 1458
rect 25865 1400 25870 1456
rect 25926 1400 30000 1456
rect 25865 1398 30000 1400
rect 25865 1395 25931 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 3969 914 4035 917
rect 0 912 4035 914
rect 0 856 3974 912
rect 4030 856 4035 912
rect 0 854 4035 856
rect 0 824 480 854
rect 3969 851 4035 854
rect 26877 914 26943 917
rect 29520 914 30000 944
rect 26877 912 30000 914
rect 26877 856 26882 912
rect 26938 856 30000 912
rect 26877 854 30000 856
rect 26877 851 26943 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 1393 370 1459 373
rect 0 368 1459 370
rect 0 312 1398 368
rect 1454 312 1459 368
rect 0 310 1459 312
rect 0 280 480 310
rect 1393 307 1459 310
rect 26785 370 26851 373
rect 29520 370 30000 400
rect 26785 368 30000 370
rect 26785 312 26790 368
rect 26846 312 30000 368
rect 26785 310 30000 312
rect 26785 307 26851 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 9628 20300 9692 20364
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 9628 19620 9692 19684
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 16436 19272 16500 19276
rect 16436 19216 16450 19272
rect 16450 19216 16500 19272
rect 16436 19212 16500 19216
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 3372 15132 3436 15196
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 17908 13908 17972 13972
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 16436 12412 16500 12476
rect 3740 12004 3804 12068
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 13308 11052 13372 11116
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 9627 20364 9693 20365
rect 9627 20300 9628 20364
rect 9692 20300 9693 20364
rect 9627 20299 9693 20300
rect 9630 19685 9690 20299
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 9627 19684 9693 19685
rect 9627 19620 9628 19684
rect 9692 19620 9693 19684
rect 9627 19619 9693 19620
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 3371 15196 3437 15197
rect 3371 15132 3372 15196
rect 3436 15132 3437 15196
rect 3371 15131 3437 15132
rect 3374 14738 3434 15131
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 3739 12068 3805 12069
rect 3739 12004 3740 12068
rect 3804 12004 3805 12068
rect 3739 12003 3805 12004
rect 3742 11338 3802 12003
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 16438 12477 16498 19211
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 17910 13973 17970 14502
rect 17907 13972 17973 13973
rect 17907 13908 17908 13972
rect 17972 13908 17973 13972
rect 17907 13907 17973 13908
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 16435 12476 16501 12477
rect 16435 12412 16436 12476
rect 16500 12412 16501 12476
rect 16435 12411 16501 12412
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 13307 11052 13308 11102
rect 13372 11052 13373 11102
rect 13307 11051 13373 11052
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 3286 14502 3522 14738
rect 3654 11102 3890 11338
rect 17822 14502 18058 14738
rect 13222 11116 13458 11338
rect 13222 11102 13308 11116
rect 13308 11102 13372 11116
rect 13372 11102 13458 11116
<< metal5 >>
rect 3244 14738 18100 14780
rect 3244 14502 3286 14738
rect 3522 14502 17822 14738
rect 18058 14502 18100 14738
rect 3244 14460 18100 14502
rect 3612 11338 13500 11380
rect 3612 11102 3654 11338
rect 3890 11102 13222 11338
rect 13458 11102 13500 11338
rect 3612 11060 13500 11102
use sky130_fd_sc_hd__buf_2  _47_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_11
timestamp 1604666999
transform 1 0 2116 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_23
timestamp 1604666999
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35
timestamp 1604666999
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604666999
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_47
timestamp 1604666999
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604666999
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1604666999
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604666999
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604666999
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604666999
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604666999
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604666999
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604666999
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604666999
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604666999
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604666999
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604666999
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604666999
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604666999
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604666999
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604666999
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604666999
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_269
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604666999
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604666999
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1604666999
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_292
timestamp 1604666999
transform 1 0 27968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604666999
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_283
timestamp 1604666999
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604666999
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 28520 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604666999
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604666999
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604666999
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604666999
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604666999
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604666999
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604666999
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604666999
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_288
timestamp 1604666999
transform 1 0 27600 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp 1604666999
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604666999
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604666999
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604666999
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604666999
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604666999
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604666999
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1604666999
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1604666999
transform 1 0 28060 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604666999
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_7
timestamp 1604666999
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_19
timestamp 1604666999
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604666999
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604666999
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604666999
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604666999
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604666999
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604666999
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604666999
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_288
timestamp 1604666999
transform 1 0 27600 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_296
timestamp 1604666999
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604666999
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604666999
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1604666999
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_17
timestamp 1604666999
transform 1 0 2668 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_29
timestamp 1604666999
transform 1 0 3772 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_41
timestamp 1604666999
transform 1 0 4876 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1604666999
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604666999
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604666999
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604666999
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604666999
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604666999
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604666999
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604666999
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604666999
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604666999
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604666999
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604666999
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_283
timestamp 1604666999
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_287
timestamp 1604666999
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604666999
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1604666999
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604666999
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604666999
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1604666999
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604666999
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604666999
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_19
timestamp 1604666999
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1604666999
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604666999
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1604666999
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604666999
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604666999
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604666999
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604666999
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_35
timestamp 1604666999
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 1604666999
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604666999
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_56
timestamp 1604666999
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1604666999
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604666999
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604666999
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604666999
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604666999
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604666999
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604666999
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604666999
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604666999
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604666999
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604666999
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604666999
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604666999
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604666999
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604666999
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604666999
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604666999
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604666999
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604666999
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_269
timestamp 1604666999
transform 1 0 25852 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604666999
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604666999
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604666999
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604666999
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_283
timestamp 1604666999
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1604666999
transform 1 0 28244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604666999
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604666999
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604666999
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1604666999
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1604666999
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604666999
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_36
timestamp 1604666999
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_40
timestamp 1604666999
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_44
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_59
timestamp 1604666999
transform 1 0 6532 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_71
timestamp 1604666999
transform 1 0 7636 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_83
timestamp 1604666999
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604666999
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604666999
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604666999
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604666999
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604666999
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604666999
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604666999
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604666999
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604666999
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604666999
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604666999
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604666999
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604666999
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604666999
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604666999
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604666999
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604666999
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1604666999
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604666999
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604666999
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604666999
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604666999
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604666999
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604666999
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1604666999
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1604666999
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1604666999
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_51
timestamp 1604666999
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_55
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604666999
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1604666999
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1604666999
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1604666999
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_106
timestamp 1604666999
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1604666999
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604666999
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604666999
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604666999
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604666999
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604666999
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604666999
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604666999
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_257
timestamp 1604666999
transform 1 0 24748 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604666999
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604666999
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_265
timestamp 1604666999
transform 1 0 25484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_273
timestamp 1604666999
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604666999
transform 1 0 27508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604666999
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604666999
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604666999
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604666999
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1604666999
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_291
timestamp 1604666999
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1604666999
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_7
timestamp 1604666999
transform 1 0 1748 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp 1604666999
transform 1 0 2208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 1604666999
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1604666999
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1604666999
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1604666999
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1604666999
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1604666999
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1604666999
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6716 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp 1604666999
transform 1 0 7544 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_78
timestamp 1604666999
transform 1 0 8280 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_81
timestamp 1604666999
transform 1 0 8556 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1604666999
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604666999
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604666999
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604666999
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604666999
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604666999
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604666999
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604666999
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604666999
transform 1 0 25300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1604666999
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604666999
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604666999
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604666999
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_18
timestamp 1604666999
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1604666999
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1604666999
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_40
timestamp 1604666999
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604666999
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604666999
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_88
timestamp 1604666999
transform 1 0 9200 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_100
timestamp 1604666999
transform 1 0 10304 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_112
timestamp 1604666999
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604666999
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604666999
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604666999
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604666999
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604666999
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604666999
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_255
timestamp 1604666999
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604666999
transform 1 0 25300 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604666999
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_259
timestamp 1604666999
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_267
timestamp 1604666999
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_271
timestamp 1604666999
transform 1 0 26036 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604666999
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604666999
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604666999
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604666999
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1604666999
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_283
timestamp 1604666999
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_291
timestamp 1604666999
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1604666999
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1604666999
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1604666999
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4324 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1604666999
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1604666999
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5888 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_44
timestamp 1604666999
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1604666999
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1604666999
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1604666999
transform 1 0 8004 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_81
timestamp 1604666999
transform 1 0 8556 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1604666999
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604666999
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604666999
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604666999
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604666999
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_178
timestamp 1604666999
transform 1 0 17480 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_186
timestamp 1604666999
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_190
timestamp 1604666999
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_198
timestamp 1604666999
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_203
timestamp 1604666999
transform 1 0 19780 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1604666999
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_215
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 21528 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1604666999
transform 1 0 21436 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1604666999
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_228
timestamp 1604666999
transform 1 0 22080 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l3_in_0_
timestamp 1604666999
transform 1 0 24380 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23552 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 23920 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_240
timestamp 1604666999
transform 1 0 23184 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_246
timestamp 1604666999
transform 1 0 23736 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_250
timestamp 1604666999
transform 1 0 24104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_262
timestamp 1604666999
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604666999
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604666999
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604666999
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604666999
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1604666999
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604666999
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1604666999
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1604666999
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1604666999
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_36
timestamp 1604666999
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_40
timestamp 1604666999
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp 1604666999
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 1604666999
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604666999
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1604666999
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6532 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7452 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1604666999
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1604666999
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1604666999
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1604666999
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1604666999
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1604666999
transform 1 0 8648 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 1604666999
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_89
timestamp 1604666999
transform 1 0 9292 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_101
timestamp 1604666999
transform 1 0 10396 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1604666999
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_100
timestamp 1604666999
transform 1 0 10304 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_112
timestamp 1604666999
transform 1 0 11408 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1604666999
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604666999
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_124
timestamp 1604666999
transform 1 0 12512 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_136
timestamp 1604666999
transform 1 0 13616 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604666999
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1604666999
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604666999
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604666999
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1604666999
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604666999
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604666999
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_180
timestamp 1604666999
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604666999
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_3_
timestamp 1604666999
transform 1 0 17848 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1604666999
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp 1604666999
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1604666999
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604666999
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1604666999
transform 1 0 20148 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1604666999
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1604666999
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_210
timestamp 1604666999
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_211
timestamp 1604666999
transform 1 0 20516 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_214
timestamp 1604666999
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_215
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1604666999
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_220
timestamp 1604666999
transform 1 0 21344 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_3_
timestamp 1604666999
transform 1 0 21528 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_2_
timestamp 1604666999
transform 1 0 21528 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_235
timestamp 1604666999
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1604666999
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_235
timestamp 1604666999
transform 1 0 22724 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_231
timestamp 1604666999
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23552 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23828 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604666999
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_256
timestamp 1604666999
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_239
timestamp 1604666999
transform 1 0 23092 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_263
timestamp 1604666999
transform 1 0 25300 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_260
timestamp 1604666999
transform 1 0 25024 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604666999
transform 1 0 25392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604666999
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_271
timestamp 1604666999
transform 1 0 26036 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_267
timestamp 1604666999
transform 1 0 25668 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 26128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604666999
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604666999
transform 1 0 26404 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1604666999
transform 1 0 27232 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_280
timestamp 1604666999
transform 1 0 26864 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_283
timestamp 1604666999
transform 1 0 27140 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_279
timestamp 1604666999
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604666999
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_291
timestamp 1604666999
transform 1 0 27876 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_295
timestamp 1604666999
transform 1 0 28244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_291
timestamp 1604666999
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604666999
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604666999
transform 1 0 27508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604666999
transform 1 0 27600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1604666999
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1604666999
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1604666999
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604666999
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604666999
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604666999
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604666999
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7452 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1604666999
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1604666999
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9016 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1604666999
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1604666999
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1604666999
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_103
timestamp 1604666999
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1604666999
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604666999
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1604666999
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1604666999
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1604666999
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1604666999
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604666999
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_171
timestamp 1604666999
transform 1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_176
timestamp 1604666999
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1604666999
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604666999
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1604666999
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l3_in_1_
timestamp 1604666999
transform 1 0 21160 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604666999
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_210
timestamp 1604666999
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1604666999
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_227
timestamp 1604666999
transform 1 0 21988 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_233
timestamp 1604666999
transform 1 0 22540 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1604666999
transform 1 0 22908 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604666999
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_1_
timestamp 1604666999
transform 1 0 26128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604666999
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604666999
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 27508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1604666999
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_285
timestamp 1604666999
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1604666999
transform 1 0 27692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1604666999
transform 1 0 28060 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604666999
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1604666999
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1604666999
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4232 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1604666999
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1604666999
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_57
timestamp 1604666999
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7084 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 1604666999
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604666999
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604666999
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1604666999
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1604666999
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_126
timestamp 1604666999
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_138
timestamp 1604666999
transform 1 0 13800 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_146
timestamp 1604666999
transform 1 0 14536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_154
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15916 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l4_in_0_
timestamp 1604666999
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_160
timestamp 1604666999
transform 1 0 15824 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1604666999
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1604666999
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_1_
timestamp 1604666999
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1604666999
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_191
timestamp 1604666999
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_196
timestamp 1604666999
transform 1 0 19136 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604666999
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1604666999
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604666999
transform 1 0 21252 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l3_in_1_
timestamp 1604666999
transform 1 0 22356 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21804 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22172 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_223
timestamp 1604666999
transform 1 0 21620 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_227
timestamp 1604666999
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_3_
timestamp 1604666999
transform 1 0 23920 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_240
timestamp 1604666999
transform 1 0 23184 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_244
timestamp 1604666999
transform 1 0 23552 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_247
timestamp 1604666999
transform 1 0 23828 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_257
timestamp 1604666999
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 24932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_261
timestamp 1604666999
transform 1 0 25116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_265
timestamp 1604666999
transform 1 0 25484 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_271
timestamp 1604666999
transform 1 0 26036 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604666999
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_285
timestamp 1604666999
transform 1 0 27324 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1604666999
transform 1 0 28428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604666999
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1604666999
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604666999
transform 1 0 4048 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604666999
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1604666999
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp 1604666999
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1604666999
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604666999
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604666999
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604666999
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1604666999
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1604666999
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8556 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_100
timestamp 1604666999
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_104
timestamp 1604666999
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_108
timestamp 1604666999
transform 1 0 11040 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1604666999
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1604666999
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604666999
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604666999
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604666999
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l3_in_1_
timestamp 1604666999
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604666999
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18952 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1604666999
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604666999
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604666999
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_230
timestamp 1604666999
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_234
timestamp 1604666999
transform 1 0 22632 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_2_
timestamp 1604666999
transform 1 0 24012 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26128 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604666999
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1604666999
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_268
timestamp 1604666999
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 28060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_291
timestamp 1604666999
transform 1 0 27876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1604666999
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 1604666999
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_10
timestamp 1604666999
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4508 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604666999
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1604666999
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1604666999
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_60
timestamp 1604666999
transform 1 0 6624 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1604666999
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1604666999
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_83
timestamp 1604666999
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1604666999
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604666999
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11316 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_102
timestamp 1604666999
transform 1 0 10488 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_108
timestamp 1604666999
transform 1 0 11040 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1604666999
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_134
timestamp 1604666999
transform 1 0 13432 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_142
timestamp 1604666999
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1604666999
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604666999
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1604666999
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16284 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_162
timestamp 1604666999
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_174
timestamp 1604666999
transform 1 0 17112 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 17848 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_201
timestamp 1604666999
transform 1 0 19596 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_207
timestamp 1604666999
transform 1 0 20148 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1604666999
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1604666999
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_238
timestamp 1604666999
transform 1 0 23000 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604666999
transform 1 0 23736 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1604666999
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_254
timestamp 1604666999
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_2_
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 25852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_267
timestamp 1604666999
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_271
timestamp 1604666999
transform 1 0 26036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_285
timestamp 1604666999
transform 1 0 27324 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1604666999
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1656 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1604666999
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_10
timestamp 1604666999
transform 1 0 2024 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_20
timestamp 1604666999
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_24
timestamp 1604666999
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1604666999
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1604666999
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1604666999
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_33
timestamp 1604666999
transform 1 0 4140 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_36
timestamp 1604666999
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1604666999
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4876 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1604666999
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_50
timestamp 1604666999
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_55
timestamp 1604666999
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_51
timestamp 1604666999
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6440 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1604666999
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1604666999
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 7268 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1604666999
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_76
timestamp 1604666999
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1604666999
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1604666999
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_87
timestamp 1604666999
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1604666999
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604666999
transform 1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1604666999
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1604666999
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9844 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1604666999
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1604666999
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1604666999
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_125
timestamp 1604666999
transform 1 0 12604 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1604666999
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1604666999
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_136
timestamp 1604666999
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604666999
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_139
timestamp 1604666999
transform 1 0 13892 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_148
timestamp 1604666999
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1604666999
transform 1 0 14352 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1604666999
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1604666999
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14996 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_167
timestamp 1604666999
transform 1 0 16468 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1604666999
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1604666999
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1604666999
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1604666999
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1604666999
transform 1 0 17020 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_176
timestamp 1604666999
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1604666999
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 17112 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18584 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_180
timestamp 1604666999
transform 1 0 17664 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_193
timestamp 1604666999
transform 1 0 18860 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604666999
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1604666999
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_203
timestamp 1604666999
transform 1 0 19780 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1604666999
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604666999
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604666999
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1604666999
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l4_in_0_
timestamp 1604666999
transform 1 0 20332 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 21160 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l1_in_1_
timestamp 1604666999
transform 1 0 21896 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1604666999
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1604666999
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_237
timestamp 1604666999
transform 1 0 22908 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_245
timestamp 1604666999
transform 1 0 23644 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_241
timestamp 1604666999
transform 1 0 23276 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_239
timestamp 1604666999
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 23092 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23736 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_256
timestamp 1604666999
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_252
timestamp 1604666999
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604666999
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604666999
transform 1 0 23920 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23920 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 25024 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l3_in_1_
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1604666999
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_271
timestamp 1604666999
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_285
timestamp 1604666999
transform 1 0 27324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_283
timestamp 1604666999
transform 1 0 27140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_279
timestamp 1604666999
transform 1 0 26772 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 27324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_289
timestamp 1604666999
transform 1 0 27692 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1604666999
transform 1 0 28244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_291
timestamp 1604666999
transform 1 0 27876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 27508 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604666999
transform 1 0 28060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604666999
transform 1 0 27508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1604666999
transform 1 0 28428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 1840 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1604666999
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604666999
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_31
timestamp 1604666999
transform 1 0 3956 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_34
timestamp 1604666999
transform 1 0 4232 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604666999
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604666999
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604666999
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604666999
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_79
timestamp 1604666999
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1604666999
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1604666999
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604666999
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604666999
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604666999
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604666999
transform 1 0 13984 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_143
timestamp 1604666999
transform 1 0 14260 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_160
timestamp 1604666999
transform 1 0 15824 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_168
timestamp 1604666999
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_172
timestamp 1604666999
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18676 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1604666999
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1604666999
transform 1 0 18400 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20240 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1604666999
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_204
timestamp 1604666999
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604666999
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21804 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604666999
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_234
timestamp 1604666999
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1604666999
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 24380 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_251
timestamp 1604666999
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_272
timestamp 1604666999
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_276
timestamp 1604666999
transform 1 0 26496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_3_
timestamp 1604666999
transform 1 0 26864 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 26680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 27876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 28244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_289
timestamp 1604666999
transform 1 0 27692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_293
timestamp 1604666999
transform 1 0 28060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1604666999
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 1472 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604666999
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 5428 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1604666999
transform 1 0 4784 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_46
timestamp 1604666999
transform 1 0 5336 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1604666999
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_70
timestamp 1604666999
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 10120 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604666999
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_117
timestamp 1604666999
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12604 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1604666999
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_144
timestamp 1604666999
transform 1 0 14352 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_158
timestamp 1604666999
transform 1 0 15640 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16376 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_185
timestamp 1604666999
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1604666999
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1604666999
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604666999
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1604666999
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21528 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 21344 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1604666999
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l1_in_2_
timestamp 1604666999
transform 1 0 24012 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_241
timestamp 1604666999
transform 1 0 23276 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_266
timestamp 1604666999
transform 1 0 25576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_262
timestamp 1604666999
transform 1 0 25208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_258
timestamp 1604666999
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604666999
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_270
timestamp 1604666999
transform 1 0 25944 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 26128 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l4_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_285
timestamp 1604666999
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1604666999
transform 1 0 27692 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1604666999
transform 1 0 28428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1604666999
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1604666999
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604666999
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1604666999
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1604666999
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_77
timestamp 1604666999
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1604666999
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8280 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1604666999
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l4_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604666999
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604666999
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604666999
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604666999
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_136
timestamp 1604666999
transform 1 0 13616 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 14812 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_141
timestamp 1604666999
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1604666999
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1604666999
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1604666999
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604666999
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19044 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604666999
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1604666999
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1604666999
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_214
timestamp 1604666999
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21712 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_220
timestamp 1604666999
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_233
timestamp 1604666999
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1604666999
transform 1 0 22908 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_241
timestamp 1604666999
transform 1 0 23276 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_254
timestamp 1604666999
transform 1 0 24472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26128 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_260
timestamp 1604666999
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1604666999
transform 1 0 25392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604666999
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 28060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_291
timestamp 1604666999
transform 1 0 27876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1604666999
transform 1 0 28244 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1604666999
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_20
timestamp 1604666999
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_24
timestamp 1604666999
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1604666999
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 4876 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_40
timestamp 1604666999
transform 1 0 4784 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_60
timestamp 1604666999
transform 1 0 6624 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1604666999
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1604666999
transform 1 0 7452 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 10212 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604666999
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11776 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_108
timestamp 1604666999
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1604666999
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 1604666999
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_139
timestamp 1604666999
transform 1 0 13892 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1604666999
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1604666999
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_177
timestamp 1604666999
transform 1 0 17388 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18400 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_185
timestamp 1604666999
transform 1 0 18124 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1604666999
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1604666999
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1604666999
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 21896 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1604666999
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_222
timestamp 1604666999
transform 1 0 21528 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_245
timestamp 1604666999
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_249
timestamp 1604666999
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1604666999
transform 1 0 24380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24840 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l3_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 26128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_267
timestamp 1604666999
transform 1 0 25668 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_271
timestamp 1604666999
transform 1 0 26036 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604666999
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_285
timestamp 1604666999
transform 1 0 27324 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1604666999
transform 1 0 28428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1604666999
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1604666999
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp 1604666999
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_35
timestamp 1604666999
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_39
timestamp 1604666999
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604666999
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604666999
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_72
timestamp 1604666999
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_77
timestamp 1604666999
transform 1 0 8188 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8464 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1604666999
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1604666999
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1604666999
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1604666999
transform 1 0 11500 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604666999
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12788 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 15272 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_146
timestamp 1604666999
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp 1604666999
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_163
timestamp 1604666999
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_167
timestamp 1604666999
transform 1 0 16468 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_173
timestamp 1604666999
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1604666999
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18400 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_207
timestamp 1604666999
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_211
timestamp 1604666999
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1604666999
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l3_in_1_
timestamp 1604666999
transform 1 0 21804 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604666999
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1604666999
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604666999
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26128 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1604666999
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_268
timestamp 1604666999
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 28060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_291
timestamp 1604666999
transform 1 0 27876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1604666999
transform 1 0 28244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1564 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1604666999
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1604666999
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_28
timestamp 1604666999
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1604666999
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_46
timestamp 1604666999
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_41
timestamp 1604666999
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_55
timestamp 1604666999
transform 1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 1604666999
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_50
timestamp 1604666999
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_67
timestamp 1604666999
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604666999
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1604666999
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604666999
transform 1 0 6992 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1604666999
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1604666999
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 8004 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1604666999
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1604666999
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1604666999
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1604666999
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10580 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l3_in_1_
timestamp 1604666999
transform 1 0 10488 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_111
timestamp 1604666999
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_115
timestamp 1604666999
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 1604666999
transform 1 0 12052 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_126
timestamp 1604666999
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1604666999
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1604666999
transform 1 0 13616 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1604666999
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13064 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 14812 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_139
timestamp 1604666999
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_144
timestamp 1604666999
transform 1 0 14352 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1604666999
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_168
timestamp 1604666999
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1604666999
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_176
timestamp 1604666999
transform 1 0 17296 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18584 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18584 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_180
timestamp 1604666999
transform 1 0 17664 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604666999
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_203
timestamp 1604666999
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1604666999
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1604666999
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1604666999
transform 1 0 20148 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1604666999
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1604666999
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604666999
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1604666999
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_219
timestamp 1604666999
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l4_in_0_
timestamp 1604666999
transform 1 0 21804 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1604666999
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_234
timestamp 1604666999
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21620 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_27_245
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_246
timestamp 1604666999
transform 1 0 23736 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_242
timestamp 1604666999
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23552 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_254
timestamp 1604666999
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1604666999
transform 1 0 24104 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23920 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23920 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1604666999
transform 1 0 25668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_267
timestamp 1604666999
transform 1 0 25668 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24840 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_271
timestamp 1604666999
transform 1 0 26036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604666999
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_271
timestamp 1604666999
transform 1 0 26036 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 25852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 26220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_1_
timestamp 1604666999
transform 1 0 26404 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l1_in_2_
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 27416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 27784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 28152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_285
timestamp 1604666999
transform 1 0 27324 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1604666999
transform 1 0 28428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_284
timestamp 1604666999
transform 1 0 27232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_288
timestamp 1604666999
transform 1 0 27600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_292
timestamp 1604666999
transform 1 0 27968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_296
timestamp 1604666999
transform 1 0 28336 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604666999
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1604666999
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_39
timestamp 1604666999
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5060 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_62
timestamp 1604666999
transform 1 0 6808 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_70
timestamp 1604666999
transform 1 0 7544 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_3_
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_84
timestamp 1604666999
transform 1 0 8832 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11500 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1604666999
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1604666999
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_110
timestamp 1604666999
transform 1 0 11224 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_132
timestamp 1604666999
transform 1 0 13248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1604666999
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_148
timestamp 1604666999
transform 1 0 14720 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604666999
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_157
timestamp 1604666999
transform 1 0 15548 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16652 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_167
timestamp 1604666999
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19136 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_188
timestamp 1604666999
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_192
timestamp 1604666999
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604666999
transform 1 0 21160 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20332 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1604666999
transform 1 0 19964 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1604666999
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 22172 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 21620 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1604666999
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1604666999
transform 1 0 21804 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_248
timestamp 1604666999
transform 1 0 23920 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_252
timestamp 1604666999
transform 1 0 24288 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l1_in_1_
timestamp 1604666999
transform 1 0 24840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_1_
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_267
timestamp 1604666999
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1604666999
transform 1 0 26036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_285
timestamp 1604666999
transform 1 0 27324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1604666999
transform 1 0 28428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1472 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1604666999
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1604666999
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604666999
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1604666999
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1604666999
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_51
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_55
timestamp 1604666999
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_65
timestamp 1604666999
transform 1 0 7084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp 1604666999
transform 1 0 7452 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_72
timestamp 1604666999
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1604666999
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8464 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1604666999
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1604666999
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1604666999
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1604666999
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1604666999
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604666999
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 15180 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_140
timestamp 1604666999
transform 1 0 13984 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_146
timestamp 1604666999
transform 1 0 14536 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1604666999
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1604666999
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_176
timestamp 1604666999
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 18768 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1604666999
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1604666999
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 20332 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1604666999
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1604666999
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_218
timestamp 1604666999
transform 1 0 21160 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_3_
timestamp 1604666999
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_223
timestamp 1604666999
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604666999
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24104 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604666999
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 25668 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 25484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1604666999
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_263
timestamp 1604666999
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 27600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 27968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_286
timestamp 1604666999
transform 1 0 27416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_290
timestamp 1604666999
transform 1 0 27784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1604666999
transform 1 0 28152 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1604666999
transform 1 0 28520 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 1564 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_14
timestamp 1604666999
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1604666999
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1604666999
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1604666999
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1604666999
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4968 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1604666999
transform 1 0 5796 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_59
timestamp 1604666999
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l4_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_64
timestamp 1604666999
transform 1 0 6992 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_72
timestamp 1604666999
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l4_in_0_
timestamp 1604666999
transform 1 0 10212 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_84
timestamp 1604666999
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 11776 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_108
timestamp 1604666999
transform 1 0 11040 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_135
timestamp 1604666999
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1604666999
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_158
timestamp 1604666999
transform 1 0 15640 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16284 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_162
timestamp 1604666999
transform 1 0 16008 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_174
timestamp 1604666999
transform 1 0 17112 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 17848 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20332 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1604666999
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_205
timestamp 1604666999
transform 1 0 19964 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1604666999
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_218
timestamp 1604666999
transform 1 0 21160 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_2_
timestamp 1604666999
transform 1 0 22080 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_237
timestamp 1604666999
transform 1 0 22908 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23920 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 23368 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_241
timestamp 1604666999
transform 1 0 23276 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_244
timestamp 1604666999
transform 1 0 23552 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_2_
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1604666999
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_285
timestamp 1604666999
transform 1 0 27324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1604666999
transform 1 0 28428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604666999
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_11
timestamp 1604666999
transform 1 0 2116 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2208 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1604666999
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1604666999
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_35
timestamp 1604666999
transform 1 0 4324 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 4784 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_49
timestamp 1604666999
transform 1 0 5612 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_74
timestamp 1604666999
transform 1 0 7912 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_77
timestamp 1604666999
transform 1 0 8188 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_85
timestamp 1604666999
transform 1 0 8924 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1604666999
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_93
timestamp 1604666999
transform 1 0 9660 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l3_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604666999
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_114
timestamp 1604666999
transform 1 0 11592 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604666999
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1604666999
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_140
timestamp 1604666999
transform 1 0 13984 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1604666999
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1604666999
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1604666999
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_175
timestamp 1604666999
transform 1 0 17204 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1604666999
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1604666999
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 19504 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21988 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_219
timestamp 1604666999
transform 1 0 21252 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_230
timestamp 1604666999
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_234
timestamp 1604666999
transform 1 0 22632 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l4_in_0_
timestamp 1604666999
transform 1 0 24656 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 24104 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_242
timestamp 1604666999
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_249
timestamp 1604666999
transform 1 0 24012 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_252
timestamp 1604666999
transform 1 0 24288 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_3_
timestamp 1604666999
transform 1 0 26312 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_265
timestamp 1604666999
transform 1 0 25484 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_270
timestamp 1604666999
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 27324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_283
timestamp 1604666999
transform 1 0 27140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_287
timestamp 1604666999
transform 1 0 27508 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1604666999
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_19
timestamp 1604666999
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1604666999
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1604666999
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1604666999
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_78
timestamp 1604666999
transform 1 0 8280 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1604666999
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_1_
timestamp 1604666999
transform 1 0 11960 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_107
timestamp 1604666999
transform 1 0 10948 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_115
timestamp 1604666999
transform 1 0 11684 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1604666999
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_131
timestamp 1604666999
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_143
timestamp 1604666999
transform 1 0 14260 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1604666999
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_163
timestamp 1604666999
transform 1 0 16100 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1604666999
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 17848 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1604666999
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_191
timestamp 1604666999
transform 1 0 18676 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1604666999
transform 1 0 19228 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_200
timestamp 1604666999
transform 1 0 19504 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1604666999
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604666999
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 23920 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_239
timestamp 1604666999
transform 1 0 23092 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_247
timestamp 1604666999
transform 1 0 23828 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1604666999
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_254
timestamp 1604666999
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l3_in_0_
timestamp 1604666999
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 25852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_267
timestamp 1604666999
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1604666999
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_279
timestamp 1604666999
transform 1 0 26772 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_291
timestamp 1604666999
transform 1 0 27876 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_6
timestamp 1604666999
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_10
timestamp 1604666999
transform 1 0 2024 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_22
timestamp 1604666999
transform 1 0 3128 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_34
timestamp 1604666999
transform 1 0 4232 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_46
timestamp 1604666999
transform 1 0 5336 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_58
timestamp 1604666999
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604666999
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604666999
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 6992 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_67
timestamp 1604666999
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_71
timestamp 1604666999
transform 1 0 7636 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604666999
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9384 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_83
timestamp 1604666999
transform 1 0 8740 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_89
timestamp 1604666999
transform 1 0 9292 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1604666999
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_97
timestamp 1604666999
transform 1 0 10028 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_109
timestamp 1604666999
transform 1 0 11132 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604666999
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_126
timestamp 1604666999
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_130
timestamp 1604666999
transform 1 0 13064 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14536 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1604666999
transform 1 0 14168 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1604666999
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_153
timestamp 1604666999
transform 1 0 15180 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604666999
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16928 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_165
timestamp 1604666999
transform 1 0 16284 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_171
timestamp 1604666999
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604666999
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604666999
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1604666999
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1604666999
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_190
timestamp 1604666999
transform 1 0 18584 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1604666999
transform 1 0 19044 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1604666999
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 19320 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 19320 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20884 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_207
timestamp 1604666999
transform 1 0 20148 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_218
timestamp 1604666999
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1604666999
transform 1 0 19504 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604666999
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_222
timestamp 1604666999
transform 1 0 21528 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_234
timestamp 1604666999
transform 1 0 22632 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604666999
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1604666999
transform 1 0 24380 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_247
timestamp 1604666999
transform 1 0 23828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_253
timestamp 1604666999
transform 1 0 24380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1604666999
transform 1 0 25392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_260
timestamp 1604666999
transform 1 0 25024 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 25576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 25392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25116 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l3_in_1_
timestamp 1604666999
transform 1 0 25576 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_272
timestamp 1604666999
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_268
timestamp 1604666999
transform 1 0 25760 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25944 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_275
timestamp 1604666999
transform 1 0 26404 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_287
timestamp 1604666999
transform 1 0 27508 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604666999
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604666999
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604666999
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604666999
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604666999
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604666999
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604666999
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604666999
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604666999
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604666999
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604666999
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604666999
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604666999
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604666999
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604666999
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604666999
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604666999
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604666999
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604666999
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604666999
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604666999
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604666999
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604666999
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604666999
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604666999
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604666999
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604666999
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14922 0 14978 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 24950 0 25006 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 prog_clk
port 82 nsew default input
rlabel metal2 s 938 23520 994 24000 6 top_grid_pin_16_
port 83 nsew default tristate
rlabel metal2 s 2778 23520 2834 24000 6 top_grid_pin_17_
port 84 nsew default tristate
rlabel metal2 s 4618 23520 4674 24000 6 top_grid_pin_18_
port 85 nsew default tristate
rlabel metal2 s 6550 23520 6606 24000 6 top_grid_pin_19_
port 86 nsew default tristate
rlabel metal2 s 8390 23520 8446 24000 6 top_grid_pin_20_
port 87 nsew default tristate
rlabel metal2 s 10230 23520 10286 24000 6 top_grid_pin_21_
port 88 nsew default tristate
rlabel metal2 s 12162 23520 12218 24000 6 top_grid_pin_22_
port 89 nsew default tristate
rlabel metal2 s 14002 23520 14058 24000 6 top_grid_pin_23_
port 90 nsew default tristate
rlabel metal2 s 15934 23520 15990 24000 6 top_grid_pin_24_
port 91 nsew default tristate
rlabel metal2 s 17774 23520 17830 24000 6 top_grid_pin_25_
port 92 nsew default tristate
rlabel metal2 s 19614 23520 19670 24000 6 top_grid_pin_26_
port 93 nsew default tristate
rlabel metal2 s 21546 23520 21602 24000 6 top_grid_pin_27_
port 94 nsew default tristate
rlabel metal2 s 23386 23520 23442 24000 6 top_grid_pin_28_
port 95 nsew default tristate
rlabel metal2 s 25226 23520 25282 24000 6 top_grid_pin_29_
port 96 nsew default tristate
rlabel metal2 s 27158 23520 27214 24000 6 top_grid_pin_30_
port 97 nsew default tristate
rlabel metal2 s 28998 23520 29054 24000 6 top_grid_pin_31_
port 98 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 99 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
