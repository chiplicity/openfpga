magic
tech EFS8A
magscale 1 2
timestamp 1604337983
<< locali >>
rect 3433 33303 3467 33405
rect 12081 31195 12115 31365
rect 9689 4063 9723 4233
<< viali >>
rect 11345 36873 11379 36907
rect 11161 36669 11195 36703
rect 11713 36669 11747 36703
rect 10977 36329 11011 36363
rect 12081 36329 12115 36363
rect 10793 36193 10827 36227
rect 11897 36193 11931 36227
rect 4353 35989 4387 36023
rect 8033 35785 8067 35819
rect 9137 35785 9171 35819
rect 10241 35785 10275 35819
rect 11345 35785 11379 35819
rect 12633 35785 12667 35819
rect 4077 35717 4111 35751
rect 1593 35649 1627 35683
rect 3525 35649 3559 35683
rect 4537 35649 4571 35683
rect 4629 35649 4663 35683
rect 1409 35581 1443 35615
rect 7849 35581 7883 35615
rect 8401 35581 8435 35615
rect 8953 35581 8987 35615
rect 9505 35581 9539 35615
rect 10057 35581 10091 35615
rect 11161 35581 11195 35615
rect 12449 35581 12483 35615
rect 2237 35445 2271 35479
rect 3893 35445 3927 35479
rect 4537 35445 4571 35479
rect 9873 35445 9907 35479
rect 10793 35445 10827 35479
rect 11989 35445 12023 35479
rect 13093 35445 13127 35479
rect 7665 35241 7699 35275
rect 9873 35241 9907 35275
rect 10977 35241 11011 35275
rect 11345 35241 11379 35275
rect 12081 35241 12115 35275
rect 13369 35241 13403 35275
rect 2053 35173 2087 35207
rect 2697 35173 2731 35207
rect 5264 35173 5298 35207
rect 7481 35105 7515 35139
rect 9689 35105 9723 35139
rect 10793 35105 10827 35139
rect 11897 35105 11931 35139
rect 13185 35105 13219 35139
rect 2605 35037 2639 35071
rect 2789 35037 2823 35071
rect 4997 35037 5031 35071
rect 1685 34901 1719 34935
rect 2237 34901 2271 34935
rect 3249 34901 3283 34935
rect 4353 34901 4387 34935
rect 6377 34901 6411 34935
rect 7021 34901 7055 34935
rect 8493 34901 8527 34935
rect 2513 34697 2547 34731
rect 4077 34697 4111 34731
rect 7849 34697 7883 34731
rect 10149 34697 10183 34731
rect 11253 34697 11287 34731
rect 13645 34697 13679 34731
rect 6929 34629 6963 34663
rect 8493 34629 8527 34663
rect 2329 34561 2363 34595
rect 2973 34561 3007 34595
rect 3525 34561 3559 34595
rect 4445 34561 4479 34595
rect 5549 34561 5583 34595
rect 9045 34561 9079 34595
rect 10517 34561 10551 34595
rect 1961 34493 1995 34527
rect 3065 34493 3099 34527
rect 4629 34493 4663 34527
rect 5457 34493 5491 34527
rect 6285 34493 6319 34527
rect 7205 34493 7239 34527
rect 8309 34493 8343 34527
rect 8769 34493 8803 34527
rect 9965 34493 9999 34527
rect 11069 34493 11103 34527
rect 11621 34493 11655 34527
rect 12081 34493 12115 34527
rect 13185 34493 13219 34527
rect 13461 34493 13495 34527
rect 7389 34425 7423 34459
rect 7481 34425 7515 34459
rect 14013 34425 14047 34459
rect 2973 34357 3007 34391
rect 3893 34357 3927 34391
rect 4537 34357 4571 34391
rect 5089 34357 5123 34391
rect 6653 34357 6687 34391
rect 8953 34357 8987 34391
rect 9781 34357 9815 34391
rect 10885 34357 10919 34391
rect 2237 34153 2271 34187
rect 3433 34153 3467 34187
rect 8217 34153 8251 34187
rect 12909 34153 12943 34187
rect 2329 34085 2363 34119
rect 4620 34085 4654 34119
rect 7082 34085 7116 34119
rect 2053 34017 2087 34051
rect 4353 34017 4387 34051
rect 9689 34017 9723 34051
rect 9956 34017 9990 34051
rect 12725 34017 12759 34051
rect 2789 33949 2823 33983
rect 3065 33949 3099 33983
rect 6837 33949 6871 33983
rect 1777 33881 1811 33915
rect 5733 33813 5767 33847
rect 8861 33813 8895 33847
rect 11069 33813 11103 33847
rect 2973 33609 3007 33643
rect 7113 33609 7147 33643
rect 11253 33609 11287 33643
rect 13645 33609 13679 33643
rect 1593 33405 1627 33439
rect 3433 33405 3467 33439
rect 3617 33405 3651 33439
rect 3985 33405 4019 33439
rect 4077 33405 4111 33439
rect 4344 33405 4378 33439
rect 8033 33405 8067 33439
rect 8493 33405 8527 33439
rect 8585 33405 8619 33439
rect 11069 33405 11103 33439
rect 13461 33405 13495 33439
rect 14013 33405 14047 33439
rect 1860 33337 1894 33371
rect 7389 33337 7423 33371
rect 7573 33337 7607 33371
rect 7665 33337 7699 33371
rect 8852 33337 8886 33371
rect 3433 33269 3467 33303
rect 5457 33269 5491 33303
rect 6193 33269 6227 33303
rect 6653 33269 6687 33303
rect 9965 33269 9999 33303
rect 10517 33269 10551 33303
rect 11621 33269 11655 33303
rect 12725 33269 12759 33303
rect 2053 33065 2087 33099
rect 4629 33065 4663 33099
rect 5089 33065 5123 33099
rect 5549 33065 5583 33099
rect 7481 33065 7515 33099
rect 8677 33065 8711 33099
rect 9505 33065 9539 33099
rect 11529 33065 11563 33099
rect 1777 32997 1811 33031
rect 2881 32997 2915 33031
rect 6561 32997 6595 33031
rect 8125 32997 8159 33031
rect 8217 32997 8251 33031
rect 9965 32997 9999 33031
rect 2973 32929 3007 32963
rect 3893 32929 3927 32963
rect 4721 32929 4755 32963
rect 10149 32929 10183 32963
rect 10416 32929 10450 32963
rect 2881 32861 2915 32895
rect 4629 32861 4663 32895
rect 6561 32861 6595 32895
rect 6653 32861 6687 32895
rect 8125 32861 8159 32895
rect 2421 32793 2455 32827
rect 3433 32793 3467 32827
rect 4169 32793 4203 32827
rect 5917 32793 5951 32827
rect 7665 32793 7699 32827
rect 6101 32725 6135 32759
rect 7113 32725 7147 32759
rect 3157 32521 3191 32555
rect 4537 32521 4571 32555
rect 8309 32521 8343 32555
rect 9229 32521 9263 32555
rect 9505 32521 9539 32555
rect 10425 32521 10459 32555
rect 10793 32521 10827 32555
rect 11161 32521 11195 32555
rect 2421 32453 2455 32487
rect 4169 32453 4203 32487
rect 5273 32453 5307 32487
rect 8861 32453 8895 32487
rect 1593 32385 1627 32419
rect 3617 32385 3651 32419
rect 5733 32385 5767 32419
rect 6285 32385 6319 32419
rect 10057 32385 10091 32419
rect 1409 32317 1443 32351
rect 2789 32317 2823 32351
rect 5089 32317 5123 32351
rect 5825 32317 5859 32351
rect 6653 32317 6687 32351
rect 6929 32317 6963 32351
rect 7196 32317 7230 32351
rect 10977 32317 11011 32351
rect 11529 32317 11563 32351
rect 3617 32249 3651 32283
rect 3709 32249 3743 32283
rect 9781 32249 9815 32283
rect 9965 32249 9999 32283
rect 5733 32181 5767 32215
rect 1593 31977 1627 32011
rect 2053 31977 2087 32011
rect 2421 31977 2455 32011
rect 3065 31977 3099 32011
rect 3525 31977 3559 32011
rect 5273 31977 5307 32011
rect 6101 31977 6135 32011
rect 6469 31977 6503 32011
rect 6911 31977 6945 32011
rect 8401 31977 8435 32011
rect 9413 31977 9447 32011
rect 10793 31977 10827 32011
rect 11069 31977 11103 32011
rect 4261 31909 4295 31943
rect 7205 31909 7239 31943
rect 7389 31909 7423 31943
rect 7481 31909 7515 31943
rect 7941 31909 7975 31943
rect 10241 31909 10275 31943
rect 11805 31909 11839 31943
rect 11897 31909 11931 31943
rect 8217 31841 8251 31875
rect 10333 31841 10367 31875
rect 11327 31841 11361 31875
rect 10241 31773 10275 31807
rect 11805 31773 11839 31807
rect 9781 31637 9815 31671
rect 12541 31637 12575 31671
rect 12909 31637 12943 31671
rect 6653 31433 6687 31467
rect 7113 31433 7147 31467
rect 10241 31433 10275 31467
rect 7389 31365 7423 31399
rect 9321 31365 9355 31399
rect 10885 31365 10919 31399
rect 12081 31365 12115 31399
rect 12541 31365 12575 31399
rect 8769 31297 8803 31331
rect 9781 31297 9815 31331
rect 11437 31297 11471 31331
rect 9137 31229 9171 31263
rect 9873 31229 9907 31263
rect 11161 31229 11195 31263
rect 11805 31229 11839 31263
rect 12909 31297 12943 31331
rect 13461 31297 13495 31331
rect 13093 31229 13127 31263
rect 12081 31161 12115 31195
rect 13001 31161 13035 31195
rect 9781 31093 9815 31127
rect 10609 31093 10643 31127
rect 11345 31093 11379 31127
rect 12173 31093 12207 31127
rect 9965 30889 9999 30923
rect 10241 30889 10275 30923
rect 12449 30889 12483 30923
rect 1685 30821 1719 30855
rect 10793 30821 10827 30855
rect 1409 30753 1443 30787
rect 11336 30753 11370 30787
rect 11069 30685 11103 30719
rect 6929 30549 6963 30583
rect 9321 30549 9355 30583
rect 1685 30345 1719 30379
rect 9873 30345 9907 30379
rect 6929 30277 6963 30311
rect 11345 30209 11379 30243
rect 3341 30141 3375 30175
rect 3433 30141 3467 30175
rect 6653 30141 6687 30175
rect 7481 30141 7515 30175
rect 9689 30141 9723 30175
rect 11161 30141 11195 30175
rect 3678 30073 3712 30107
rect 6285 30073 6319 30107
rect 7205 30073 7239 30107
rect 7389 30073 7423 30107
rect 9321 30073 9355 30107
rect 10149 30073 10183 30107
rect 10425 30073 10459 30107
rect 4813 30005 4847 30039
rect 10333 30005 10367 30039
rect 11897 30005 11931 30039
rect 10323 29801 10357 29835
rect 12357 29801 12391 29835
rect 5448 29733 5482 29767
rect 8217 29733 8251 29767
rect 10609 29733 10643 29767
rect 10793 29733 10827 29767
rect 5181 29665 5215 29699
rect 8309 29665 8343 29699
rect 12173 29665 12207 29699
rect 8125 29597 8159 29631
rect 10885 29597 10919 29631
rect 12449 29597 12483 29631
rect 7757 29529 7791 29563
rect 11897 29529 11931 29563
rect 3433 29461 3467 29495
rect 6561 29461 6595 29495
rect 7113 29461 7147 29495
rect 7481 29461 7515 29495
rect 8677 29461 8711 29495
rect 9965 29461 9999 29495
rect 6929 29257 6963 29291
rect 9965 29257 9999 29291
rect 12633 29257 12667 29291
rect 10609 29189 10643 29223
rect 4169 29121 4203 29155
rect 4261 29121 4295 29155
rect 6653 29121 6687 29155
rect 7389 29121 7423 29155
rect 10885 29121 10919 29155
rect 8401 29053 8435 29087
rect 8585 29053 8619 29087
rect 4506 28985 4540 29019
rect 6285 28985 6319 29019
rect 7481 28985 7515 29019
rect 7941 28985 7975 29019
rect 8830 28985 8864 29019
rect 11897 28985 11931 29019
rect 5641 28917 5675 28951
rect 7389 28917 7423 28951
rect 12265 28917 12299 28951
rect 6929 28713 6963 28747
rect 8493 28713 8527 28747
rect 10241 28713 10275 28747
rect 12357 28713 12391 28747
rect 1685 28645 1719 28679
rect 5365 28645 5399 28679
rect 11222 28645 11256 28679
rect 1409 28577 1443 28611
rect 4353 28577 4387 28611
rect 6561 28577 6595 28611
rect 7380 28577 7414 28611
rect 10977 28577 11011 28611
rect 5273 28509 5307 28543
rect 5457 28509 5491 28543
rect 7113 28509 7147 28543
rect 4721 28373 4755 28407
rect 4905 28373 4939 28407
rect 5825 28373 5859 28407
rect 10609 28373 10643 28407
rect 5917 28169 5951 28203
rect 7665 28169 7699 28203
rect 7941 28169 7975 28203
rect 10149 28169 10183 28203
rect 10425 28169 10459 28203
rect 10701 28169 10735 28203
rect 11621 28169 11655 28203
rect 4997 28101 5031 28135
rect 7113 28033 7147 28067
rect 8125 28033 8159 28067
rect 11253 28033 11287 28067
rect 2421 27965 2455 27999
rect 2666 27897 2700 27931
rect 4445 27897 4479 27931
rect 5273 27897 5307 27931
rect 5457 27897 5491 27931
rect 5549 27897 5583 27931
rect 6285 27897 6319 27931
rect 8370 27897 8404 27931
rect 10977 27897 11011 27931
rect 1685 27829 1719 27863
rect 2329 27829 2363 27863
rect 3801 27829 3835 27863
rect 4813 27829 4847 27863
rect 9505 27829 9539 27863
rect 11161 27829 11195 27863
rect 11069 27625 11103 27659
rect 5549 27557 5583 27591
rect 7113 27557 7147 27591
rect 8217 27557 8251 27591
rect 10241 27557 10275 27591
rect 10333 27557 10367 27591
rect 5365 27489 5399 27523
rect 5641 27421 5675 27455
rect 6469 27421 6503 27455
rect 7021 27421 7055 27455
rect 7205 27421 7239 27455
rect 10149 27421 10183 27455
rect 6653 27353 6687 27387
rect 9781 27353 9815 27387
rect 2513 27285 2547 27319
rect 4813 27285 4847 27319
rect 5089 27285 5123 27319
rect 7665 27285 7699 27319
rect 4353 27081 4387 27115
rect 6653 27081 6687 27115
rect 9781 27081 9815 27115
rect 10425 27081 10459 27115
rect 4629 27013 4663 27047
rect 6929 27013 6963 27047
rect 10057 27013 10091 27047
rect 5089 26945 5123 26979
rect 5917 26945 5951 26979
rect 7389 26945 7423 26979
rect 8217 26945 8251 26979
rect 4077 26877 4111 26911
rect 5181 26877 5215 26911
rect 3709 26809 3743 26843
rect 5089 26809 5123 26843
rect 7481 26809 7515 26843
rect 5549 26741 5583 26775
rect 7389 26741 7423 26775
rect 7849 26741 7883 26775
rect 6561 26537 6595 26571
rect 4813 26469 4847 26503
rect 7573 26469 7607 26503
rect 10241 26469 10275 26503
rect 6929 26401 6963 26435
rect 10333 26401 10367 26435
rect 4813 26333 4847 26367
rect 4905 26333 4939 26367
rect 7481 26333 7515 26367
rect 7665 26333 7699 26367
rect 10149 26333 10183 26367
rect 4353 26265 4387 26299
rect 5365 26265 5399 26299
rect 7113 26265 7147 26299
rect 9781 26265 9815 26299
rect 2789 26197 2823 26231
rect 8033 26197 8067 26231
rect 2237 25993 2271 26027
rect 4077 25993 4111 26027
rect 4997 25993 5031 26027
rect 7389 25993 7423 26027
rect 4721 25925 4755 25959
rect 7113 25925 7147 25959
rect 9689 25925 9723 25959
rect 9965 25925 9999 25959
rect 1593 25857 1627 25891
rect 6285 25857 6319 25891
rect 7849 25857 7883 25891
rect 10333 25857 10367 25891
rect 1409 25789 1443 25823
rect 2697 25789 2731 25823
rect 9045 25789 9079 25823
rect 2964 25721 2998 25755
rect 6653 25721 6687 25755
rect 7849 25721 7883 25755
rect 7941 25721 7975 25755
rect 10517 25721 10551 25755
rect 2605 25653 2639 25687
rect 5365 25653 5399 25687
rect 8401 25653 8435 25687
rect 9321 25653 9355 25687
rect 10425 25653 10459 25687
rect 10977 25653 11011 25687
rect 2973 25449 3007 25483
rect 5181 25449 5215 25483
rect 8033 25449 8067 25483
rect 9965 25449 9999 25483
rect 4629 25381 4663 25415
rect 6070 25381 6104 25415
rect 4721 25313 4755 25347
rect 5825 25313 5859 25347
rect 10793 25313 10827 25347
rect 11060 25313 11094 25347
rect 2973 25245 3007 25279
rect 3065 25245 3099 25279
rect 4629 25245 4663 25279
rect 1961 25177 1995 25211
rect 2513 25177 2547 25211
rect 2329 25109 2363 25143
rect 3525 25109 3559 25143
rect 4169 25109 4203 25143
rect 7205 25109 7239 25143
rect 10333 25109 10367 25143
rect 12173 25109 12207 25143
rect 12817 25109 12851 25143
rect 2513 24905 2547 24939
rect 4169 24905 4203 24939
rect 5641 24905 5675 24939
rect 6561 24905 6595 24939
rect 7389 24905 7423 24939
rect 8033 24905 8067 24939
rect 10793 24905 10827 24939
rect 12541 24905 12575 24939
rect 2789 24837 2823 24871
rect 6285 24837 6319 24871
rect 9597 24837 9631 24871
rect 3341 24769 3375 24803
rect 7113 24769 7147 24803
rect 12173 24769 12207 24803
rect 1409 24701 1443 24735
rect 3065 24701 3099 24735
rect 3709 24701 3743 24735
rect 4261 24701 4295 24735
rect 4528 24701 4562 24735
rect 8309 24701 8343 24735
rect 8953 24701 8987 24735
rect 9873 24701 9907 24735
rect 11805 24701 11839 24735
rect 13093 24701 13127 24735
rect 1685 24633 1719 24667
rect 3249 24633 3283 24667
rect 8585 24633 8619 24667
rect 10149 24633 10183 24667
rect 12817 24633 12851 24667
rect 7849 24565 7883 24599
rect 8493 24565 8527 24599
rect 9413 24565 9447 24599
rect 10057 24565 10091 24599
rect 11161 24565 11195 24599
rect 13001 24565 13035 24599
rect 1593 24361 1627 24395
rect 2035 24361 2069 24395
rect 2973 24361 3007 24395
rect 4077 24361 4111 24395
rect 4629 24361 4663 24395
rect 4905 24361 4939 24395
rect 5917 24361 5951 24395
rect 8493 24361 8527 24395
rect 12541 24361 12575 24395
rect 2513 24293 2547 24327
rect 2605 24293 2639 24327
rect 3341 24293 3375 24327
rect 7358 24293 7392 24327
rect 2329 24225 2363 24259
rect 7113 24225 7147 24259
rect 11161 24225 11195 24259
rect 11428 24225 11462 24259
rect 5917 24157 5951 24191
rect 6009 24157 6043 24191
rect 9873 24157 9907 24191
rect 5457 24021 5491 24055
rect 10885 24021 10919 24055
rect 2329 23817 2363 23851
rect 3617 23817 3651 23851
rect 4813 23817 4847 23851
rect 5825 23817 5859 23851
rect 7297 23817 7331 23851
rect 7941 23817 7975 23851
rect 11805 23817 11839 23851
rect 2053 23749 2087 23783
rect 4629 23749 4663 23783
rect 7665 23749 7699 23783
rect 10609 23749 10643 23783
rect 10885 23749 10919 23783
rect 12541 23749 12575 23783
rect 2789 23681 2823 23715
rect 3249 23681 3283 23715
rect 5365 23681 5399 23715
rect 8493 23681 8527 23715
rect 8861 23681 8895 23715
rect 13093 23681 13127 23715
rect 2881 23613 2915 23647
rect 4261 23613 4295 23647
rect 6101 23613 6135 23647
rect 8217 23613 8251 23647
rect 11161 23613 11195 23647
rect 12265 23613 12299 23647
rect 12817 23613 12851 23647
rect 1685 23545 1719 23579
rect 2789 23545 2823 23579
rect 5089 23545 5123 23579
rect 5273 23545 5307 23579
rect 6837 23545 6871 23579
rect 11437 23545 11471 23579
rect 8401 23477 8435 23511
rect 10241 23477 10275 23511
rect 11345 23477 11379 23511
rect 13001 23477 13035 23511
rect 1961 23273 1995 23307
rect 5089 23273 5123 23307
rect 5439 23273 5473 23307
rect 5917 23273 5951 23307
rect 7205 23273 7239 23307
rect 7941 23273 7975 23307
rect 9965 23273 9999 23307
rect 12081 23273 12115 23307
rect 12541 23273 12575 23307
rect 13001 23273 13035 23307
rect 2973 23205 3007 23239
rect 8585 23205 8619 23239
rect 11069 23205 11103 23239
rect 2329 23137 2363 23171
rect 2789 23137 2823 23171
rect 4813 23137 4847 23171
rect 8401 23137 8435 23171
rect 11161 23137 11195 23171
rect 3065 23069 3099 23103
rect 5917 23069 5951 23103
rect 6009 23069 6043 23103
rect 8677 23069 8711 23103
rect 11069 23069 11103 23103
rect 2513 23001 2547 23035
rect 11529 23001 11563 23035
rect 8125 22933 8159 22967
rect 10609 22933 10643 22967
rect 2513 22729 2547 22763
rect 2881 22729 2915 22763
rect 5825 22729 5859 22763
rect 6101 22729 6135 22763
rect 7205 22729 7239 22763
rect 7849 22729 7883 22763
rect 8125 22729 8159 22763
rect 9045 22729 9079 22763
rect 10701 22729 10735 22763
rect 11345 22729 11379 22763
rect 5457 22661 5491 22695
rect 9689 22661 9723 22695
rect 9505 22593 9539 22627
rect 10241 22593 10275 22627
rect 11069 22593 11103 22627
rect 7573 22525 7607 22559
rect 8401 22525 8435 22559
rect 9965 22525 9999 22559
rect 8677 22457 8711 22491
rect 10149 22457 10183 22491
rect 3157 22389 3191 22423
rect 8585 22389 8619 22423
rect 4629 22185 4663 22219
rect 8309 22185 8343 22219
rect 8677 22185 8711 22219
rect 9965 22185 9999 22219
rect 10333 22185 10367 22219
rect 2973 22117 3007 22151
rect 6193 22117 6227 22151
rect 7757 22117 7791 22151
rect 11130 22117 11164 22151
rect 7573 22049 7607 22083
rect 10885 22049 10919 22083
rect 2973 21981 3007 22015
rect 3065 21981 3099 22015
rect 4537 21981 4571 22015
rect 4721 21981 4755 22015
rect 6101 21981 6135 22015
rect 6285 21981 6319 22015
rect 7849 21981 7883 22015
rect 2513 21913 2547 21947
rect 4169 21913 4203 21947
rect 3893 21845 3927 21879
rect 5733 21845 5767 21879
rect 7297 21845 7331 21879
rect 12265 21845 12299 21879
rect 2145 21641 2179 21675
rect 4905 21641 4939 21675
rect 6193 21641 6227 21675
rect 6653 21641 6687 21675
rect 10977 21641 11011 21675
rect 11253 21641 11287 21675
rect 5917 21573 5951 21607
rect 8217 21573 8251 21607
rect 9781 21573 9815 21607
rect 3065 21505 3099 21539
rect 5549 21505 5583 21539
rect 7941 21505 7975 21539
rect 10241 21505 10275 21539
rect 3525 21437 3559 21471
rect 3792 21437 3826 21471
rect 9597 21437 9631 21471
rect 10333 21437 10367 21471
rect 8493 21369 8527 21403
rect 8769 21369 8803 21403
rect 9229 21369 9263 21403
rect 10241 21369 10275 21403
rect 2421 21301 2455 21335
rect 3341 21301 3375 21335
rect 7297 21301 7331 21335
rect 7573 21301 7607 21335
rect 8677 21301 8711 21335
rect 2513 21097 2547 21131
rect 5457 21097 5491 21131
rect 1685 21029 1719 21063
rect 7113 21029 7147 21063
rect 9956 21029 9990 21063
rect 1409 20961 1443 20995
rect 4344 20961 4378 20995
rect 7205 20961 7239 20995
rect 9689 20961 9723 20995
rect 3617 20893 3651 20927
rect 4077 20893 4111 20927
rect 6377 20893 6411 20927
rect 7113 20893 7147 20927
rect 6653 20825 6687 20859
rect 6009 20757 6043 20791
rect 8217 20757 8251 20791
rect 8585 20757 8619 20791
rect 11069 20757 11103 20791
rect 5273 20553 5307 20587
rect 8033 20553 8067 20587
rect 10517 20553 10551 20587
rect 3709 20485 3743 20519
rect 10241 20485 10275 20519
rect 2237 20417 2271 20451
rect 5733 20417 5767 20451
rect 6837 20417 6871 20451
rect 8217 20417 8251 20451
rect 1409 20349 1443 20383
rect 8484 20349 8518 20383
rect 1685 20281 1719 20315
rect 3525 20281 3559 20315
rect 3985 20281 4019 20315
rect 4169 20281 4203 20315
rect 4261 20281 4295 20315
rect 5733 20281 5767 20315
rect 5825 20281 5859 20315
rect 6285 20281 6319 20315
rect 7757 20281 7791 20315
rect 3157 20213 3191 20247
rect 4629 20213 4663 20247
rect 5089 20213 5123 20247
rect 6653 20213 6687 20247
rect 7389 20213 7423 20247
rect 9597 20213 9631 20247
rect 1593 20009 1627 20043
rect 3709 20009 3743 20043
rect 4353 20009 4387 20043
rect 6193 20009 6227 20043
rect 6837 20009 6871 20043
rect 9413 20009 9447 20043
rect 12081 20009 12115 20043
rect 4721 19941 4755 19975
rect 5080 19941 5114 19975
rect 7849 19941 7883 19975
rect 7941 19941 7975 19975
rect 10701 19873 10735 19907
rect 10968 19873 11002 19907
rect 4813 19805 4847 19839
rect 7849 19805 7883 19839
rect 7389 19737 7423 19771
rect 5273 19465 5307 19499
rect 6653 19465 6687 19499
rect 10701 19465 10735 19499
rect 2237 19261 2271 19295
rect 2329 19261 2363 19295
rect 4905 19261 4939 19295
rect 6837 19261 6871 19295
rect 9395 19261 9429 19295
rect 9965 19261 9999 19295
rect 2596 19193 2630 19227
rect 7082 19193 7116 19227
rect 8769 19193 8803 19227
rect 9689 19193 9723 19227
rect 3709 19125 3743 19159
rect 8217 19125 8251 19159
rect 9229 19125 9263 19159
rect 9873 19125 9907 19159
rect 11069 19125 11103 19159
rect 4813 18921 4847 18955
rect 6837 18921 6871 18955
rect 7297 18921 7331 18955
rect 8493 18921 8527 18955
rect 9321 18921 9355 18955
rect 7757 18853 7791 18887
rect 7941 18853 7975 18887
rect 10241 18853 10275 18887
rect 8033 18785 8067 18819
rect 4077 18717 4111 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 7481 18649 7515 18683
rect 2421 18581 2455 18615
rect 9781 18581 9815 18615
rect 1961 18377 1995 18411
rect 6653 18377 6687 18411
rect 9965 18377 9999 18411
rect 10885 18377 10919 18411
rect 11253 18377 11287 18411
rect 4905 18309 4939 18343
rect 7297 18309 7331 18343
rect 8309 18309 8343 18343
rect 2053 18241 2087 18275
rect 5273 18241 5307 18275
rect 7665 18241 7699 18275
rect 8861 18241 8895 18275
rect 4353 18173 4387 18207
rect 5457 18173 5491 18207
rect 8585 18173 8619 18207
rect 9413 18173 9447 18207
rect 10517 18173 10551 18207
rect 2298 18105 2332 18139
rect 4721 18105 4755 18139
rect 5365 18105 5399 18139
rect 8033 18105 8067 18139
rect 8769 18105 8803 18139
rect 10241 18105 10275 18139
rect 3433 18037 3467 18071
rect 9689 18037 9723 18071
rect 10425 18037 10459 18071
rect 5365 17833 5399 17867
rect 7481 17833 7515 17867
rect 9873 17833 9907 17867
rect 12265 17833 12299 17867
rect 2973 17765 3007 17799
rect 5457 17765 5491 17799
rect 8585 17765 8619 17799
rect 5181 17697 5215 17731
rect 8401 17697 8435 17731
rect 10333 17697 10367 17731
rect 10793 17697 10827 17731
rect 11152 17697 11186 17731
rect 2973 17629 3007 17663
rect 3065 17629 3099 17663
rect 8677 17629 8711 17663
rect 10885 17629 10919 17663
rect 1777 17561 1811 17595
rect 2053 17493 2087 17527
rect 2513 17493 2547 17527
rect 4905 17493 4939 17527
rect 8125 17493 8159 17527
rect 9321 17493 9355 17527
rect 1685 17289 1719 17323
rect 2053 17289 2087 17323
rect 3525 17289 3559 17323
rect 5089 17289 5123 17323
rect 7389 17289 7423 17323
rect 7757 17289 7791 17323
rect 9321 17289 9355 17323
rect 10885 17289 10919 17323
rect 2237 17221 2271 17255
rect 8125 17221 8159 17255
rect 3709 17153 3743 17187
rect 9137 17153 9171 17187
rect 9873 17153 9907 17187
rect 2513 17085 2547 17119
rect 3976 17085 4010 17119
rect 11161 17085 11195 17119
rect 2789 17017 2823 17051
rect 8769 17017 8803 17051
rect 9597 17017 9631 17051
rect 9781 17017 9815 17051
rect 10333 17017 10367 17051
rect 11437 17017 11471 17051
rect 11897 17017 11931 17051
rect 12449 17017 12483 17051
rect 2697 16949 2731 16983
rect 3157 16949 3191 16983
rect 5733 16949 5767 16983
rect 10701 16949 10735 16983
rect 11345 16949 11379 16983
rect 12173 16949 12207 16983
rect 1685 16745 1719 16779
rect 3801 16745 3835 16779
rect 5457 16745 5491 16779
rect 9321 16745 9355 16779
rect 12173 16745 12207 16779
rect 2329 16677 2363 16711
rect 4629 16677 4663 16711
rect 4721 16677 4755 16711
rect 5089 16677 5123 16711
rect 5886 16677 5920 16711
rect 4445 16609 4479 16643
rect 5641 16609 5675 16643
rect 8125 16609 8159 16643
rect 11049 16609 11083 16643
rect 2237 16541 2271 16575
rect 2421 16541 2455 16575
rect 10793 16541 10827 16575
rect 1869 16405 1903 16439
rect 3157 16405 3191 16439
rect 4169 16405 4203 16439
rect 7021 16405 7055 16439
rect 7665 16405 7699 16439
rect 2237 16201 2271 16235
rect 2513 16201 2547 16235
rect 3157 16201 3191 16235
rect 4169 16201 4203 16235
rect 5641 16201 5675 16235
rect 6009 16201 6043 16235
rect 9413 16201 9447 16235
rect 11253 16201 11287 16235
rect 4721 16133 4755 16167
rect 7389 16133 7423 16167
rect 1593 16065 1627 16099
rect 2973 16065 3007 16099
rect 3617 16065 3651 16099
rect 5273 16065 5307 16099
rect 7849 16065 7883 16099
rect 8309 16065 8343 16099
rect 9965 16065 9999 16099
rect 1409 15997 1443 16031
rect 4997 15997 5031 16031
rect 6377 15997 6411 16031
rect 7205 15997 7239 16031
rect 7941 15997 7975 16031
rect 3709 15929 3743 15963
rect 5181 15929 5215 15963
rect 7849 15929 7883 15963
rect 9229 15929 9263 15963
rect 9689 15929 9723 15963
rect 3617 15861 3651 15895
rect 4445 15861 4479 15895
rect 9873 15861 9907 15895
rect 10885 15861 10919 15895
rect 3433 15657 3467 15691
rect 4353 15657 4387 15691
rect 5365 15657 5399 15691
rect 8493 15657 8527 15691
rect 2605 15589 2639 15623
rect 3157 15589 3191 15623
rect 4721 15589 4755 15623
rect 5089 15589 5123 15623
rect 10241 15589 10275 15623
rect 7380 15521 7414 15555
rect 10333 15521 10367 15555
rect 11520 15521 11554 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 7113 15453 7147 15487
rect 10149 15453 10183 15487
rect 11253 15453 11287 15487
rect 1869 15385 1903 15419
rect 2145 15385 2179 15419
rect 9781 15385 9815 15419
rect 9413 15317 9447 15351
rect 12633 15317 12667 15351
rect 2145 15113 2179 15147
rect 6653 15113 6687 15147
rect 7113 15113 7147 15147
rect 7849 15113 7883 15147
rect 10057 15113 10091 15147
rect 11621 15113 11655 15147
rect 2973 15045 3007 15079
rect 4721 15045 4755 15079
rect 3433 14977 3467 15011
rect 4537 14977 4571 15011
rect 5089 14977 5123 15011
rect 5273 14977 5307 15011
rect 2789 14909 2823 14943
rect 3525 14909 3559 14943
rect 5641 14909 5675 14943
rect 8125 14909 8159 14943
rect 8769 14909 8803 14943
rect 5181 14841 5215 14875
rect 8401 14841 8435 14875
rect 9137 14841 9171 14875
rect 1685 14773 1719 14807
rect 3433 14773 3467 14807
rect 3893 14773 3927 14807
rect 7665 14773 7699 14807
rect 8309 14773 8343 14807
rect 9781 14773 9815 14807
rect 10425 14773 10459 14807
rect 11253 14773 11287 14807
rect 1593 14569 1627 14603
rect 2145 14569 2179 14603
rect 6653 14569 6687 14603
rect 7481 14569 7515 14603
rect 8401 14569 8435 14603
rect 13461 14569 13495 14603
rect 3249 14501 3283 14535
rect 5089 14501 5123 14535
rect 5917 14501 5951 14535
rect 6745 14501 6779 14535
rect 8217 14501 8251 14535
rect 10057 14501 10091 14535
rect 10241 14501 10275 14535
rect 12348 14501 12382 14535
rect 12081 14433 12115 14467
rect 4997 14365 5031 14399
rect 5181 14365 5215 14399
rect 6653 14365 6687 14399
rect 8493 14365 8527 14399
rect 10333 14365 10367 14399
rect 5641 14297 5675 14331
rect 6193 14297 6227 14331
rect 7941 14297 7975 14331
rect 9781 14297 9815 14331
rect 2973 14229 3007 14263
rect 4629 14229 4663 14263
rect 7205 14229 7239 14263
rect 3341 14025 3375 14059
rect 6193 14025 6227 14059
rect 8033 14025 8067 14059
rect 8309 14025 8343 14059
rect 9321 14025 9355 14059
rect 9781 14025 9815 14059
rect 11253 14025 11287 14059
rect 12173 14025 12207 14059
rect 5273 13957 5307 13991
rect 7021 13957 7055 13991
rect 12633 13957 12667 13991
rect 2237 13889 2271 13923
rect 3893 13889 3927 13923
rect 5733 13889 5767 13923
rect 7389 13889 7423 13923
rect 7573 13889 7607 13923
rect 1409 13821 1443 13855
rect 1685 13821 1719 13855
rect 3617 13821 3651 13855
rect 4629 13821 4663 13855
rect 5089 13821 5123 13855
rect 6653 13821 6687 13855
rect 8677 13821 8711 13855
rect 9873 13821 9907 13855
rect 3157 13753 3191 13787
rect 3801 13753 3835 13787
rect 5825 13753 5859 13787
rect 10140 13753 10174 13787
rect 2789 13685 2823 13719
rect 5733 13685 5767 13719
rect 7481 13685 7515 13719
rect 4629 13481 4663 13515
rect 4997 13481 5031 13515
rect 7941 13481 7975 13515
rect 10333 13481 10367 13515
rect 10609 13481 10643 13515
rect 2881 13413 2915 13447
rect 5702 13413 5736 13447
rect 11336 13413 11370 13447
rect 2973 13345 3007 13379
rect 5457 13345 5491 13379
rect 2881 13277 2915 13311
rect 11069 13277 11103 13311
rect 2237 13209 2271 13243
rect 3341 13209 3375 13243
rect 1685 13141 1719 13175
rect 2421 13141 2455 13175
rect 5365 13141 5399 13175
rect 6837 13141 6871 13175
rect 7389 13141 7423 13175
rect 9873 13141 9907 13175
rect 12449 13141 12483 13175
rect 1593 12937 1627 12971
rect 6929 12937 6963 12971
rect 7941 12937 7975 12971
rect 9965 12937 9999 12971
rect 11529 12937 11563 12971
rect 2973 12869 3007 12903
rect 5825 12869 5859 12903
rect 6561 12869 6595 12903
rect 6193 12801 6227 12835
rect 7297 12801 7331 12835
rect 3065 12733 3099 12767
rect 3321 12733 3355 12767
rect 5549 12733 5583 12767
rect 7481 12733 7515 12767
rect 8585 12733 8619 12767
rect 11069 12733 11103 12767
rect 1869 12665 1903 12699
rect 2145 12665 2179 12699
rect 8830 12665 8864 12699
rect 2053 12597 2087 12631
rect 2513 12597 2547 12631
rect 4445 12597 4479 12631
rect 7389 12597 7423 12631
rect 8401 12597 8435 12631
rect 1961 12393 1995 12427
rect 2311 12393 2345 12427
rect 3249 12393 3283 12427
rect 6929 12393 6963 12427
rect 8585 12393 8619 12427
rect 1685 12325 1719 12359
rect 2789 12325 2823 12359
rect 4997 12325 5031 12359
rect 7849 12325 7883 12359
rect 10333 12325 10367 12359
rect 4813 12257 4847 12291
rect 7665 12257 7699 12291
rect 10425 12257 10459 12291
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 5089 12189 5123 12223
rect 7941 12189 7975 12223
rect 10241 12189 10275 12223
rect 10793 12189 10827 12223
rect 7389 12121 7423 12155
rect 11161 12121 11195 12155
rect 4537 12053 4571 12087
rect 9873 12053 9907 12087
rect 2697 11849 2731 11883
rect 4353 11849 4387 11883
rect 4905 11849 4939 11883
rect 5273 11849 5307 11883
rect 6285 11849 6319 11883
rect 7757 11849 7791 11883
rect 9229 11849 9263 11883
rect 10425 11781 10459 11815
rect 1593 11713 1627 11747
rect 7849 11713 7883 11747
rect 1409 11645 1443 11679
rect 2973 11645 3007 11679
rect 10701 11645 10735 11679
rect 3240 11577 3274 11611
rect 7389 11577 7423 11611
rect 8094 11577 8128 11611
rect 10149 11577 10183 11611
rect 10977 11577 11011 11611
rect 2329 11509 2363 11543
rect 6653 11509 6687 11543
rect 9873 11509 9907 11543
rect 10885 11509 10919 11543
rect 11345 11509 11379 11543
rect 12449 11509 12483 11543
rect 1593 11305 1627 11339
rect 2329 11305 2363 11339
rect 3065 11305 3099 11339
rect 4537 11305 4571 11339
rect 6837 11305 6871 11339
rect 7665 11305 7699 11339
rect 8493 11305 8527 11339
rect 9965 11305 9999 11339
rect 5724 11237 5758 11271
rect 10977 11237 11011 11271
rect 12063 11237 12097 11271
rect 12541 11237 12575 11271
rect 12633 11237 12667 11271
rect 5457 11169 5491 11203
rect 11069 11169 11103 11203
rect 8401 11101 8435 11135
rect 8585 11101 8619 11135
rect 10885 11101 10919 11135
rect 12541 11101 12575 11135
rect 3341 11033 3375 11067
rect 8033 11033 8067 11067
rect 10517 11033 10551 11067
rect 11897 11033 11931 11067
rect 11437 10965 11471 10999
rect 13093 10965 13127 10999
rect 5549 10761 5583 10795
rect 6101 10761 6135 10795
rect 8953 10761 8987 10795
rect 9781 10761 9815 10795
rect 12081 10761 12115 10795
rect 10149 10693 10183 10727
rect 10425 10693 10459 10727
rect 10793 10693 10827 10727
rect 12541 10693 12575 10727
rect 7573 10625 7607 10659
rect 11253 10625 11287 10659
rect 11345 10625 11379 10659
rect 13093 10625 13127 10659
rect 12817 10557 12851 10591
rect 13461 10557 13495 10591
rect 7113 10489 7147 10523
rect 7840 10489 7874 10523
rect 11253 10489 11287 10523
rect 4537 10421 4571 10455
rect 5641 10421 5675 10455
rect 7389 10421 7423 10455
rect 13001 10421 13035 10455
rect 1685 10217 1719 10251
rect 8401 10217 8435 10251
rect 8677 10217 8711 10251
rect 10425 10217 10459 10251
rect 10977 10217 11011 10251
rect 4629 10149 4663 10183
rect 6644 10149 6678 10183
rect 11253 10149 11287 10183
rect 11989 10149 12023 10183
rect 12081 10149 12115 10183
rect 13369 10149 13403 10183
rect 13553 10149 13587 10183
rect 4445 10081 4479 10115
rect 6377 10081 6411 10115
rect 10517 10081 10551 10115
rect 13645 10081 13679 10115
rect 4721 10013 4755 10047
rect 10333 10013 10367 10047
rect 11897 10013 11931 10047
rect 3893 9945 3927 9979
rect 9965 9945 9999 9979
rect 13093 9945 13127 9979
rect 2973 9877 3007 9911
rect 4169 9877 4203 9911
rect 5181 9877 5215 9911
rect 7757 9877 7791 9911
rect 11529 9877 11563 9911
rect 12449 9877 12483 9911
rect 12817 9877 12851 9911
rect 6101 9673 6135 9707
rect 8493 9673 8527 9707
rect 9873 9673 9907 9707
rect 10241 9673 10275 9707
rect 10609 9673 10643 9707
rect 11437 9673 11471 9707
rect 12725 9673 12759 9707
rect 2973 9605 3007 9639
rect 4537 9605 4571 9639
rect 6377 9605 6411 9639
rect 7481 9605 7515 9639
rect 11805 9605 11839 9639
rect 12173 9605 12207 9639
rect 13001 9605 13035 9639
rect 1593 9537 1627 9571
rect 3525 9537 3559 9571
rect 4997 9537 5031 9571
rect 8033 9537 8067 9571
rect 1409 9469 1443 9503
rect 2421 9469 2455 9503
rect 8769 9469 8803 9503
rect 13369 9469 13403 9503
rect 13921 9469 13955 9503
rect 2789 9401 2823 9435
rect 3249 9401 3283 9435
rect 4997 9401 5031 9435
rect 5089 9401 5123 9435
rect 7757 9401 7791 9435
rect 7941 9401 7975 9435
rect 3433 9333 3467 9367
rect 4169 9333 4203 9367
rect 5457 9333 5491 9367
rect 7205 9333 7239 9367
rect 13553 9333 13587 9367
rect 2053 9129 2087 9163
rect 2973 9129 3007 9163
rect 5641 9129 5675 9163
rect 6929 9129 6963 9163
rect 11897 9129 11931 9163
rect 13645 9129 13679 9163
rect 1685 9061 1719 9095
rect 3065 9061 3099 9095
rect 4506 9061 4540 9095
rect 8033 9061 8067 9095
rect 10241 9061 10275 9095
rect 11989 9061 12023 9095
rect 13185 9061 13219 9095
rect 3893 8993 3927 9027
rect 4261 8993 4295 9027
rect 10057 8993 10091 9027
rect 11713 8993 11747 9027
rect 12898 8993 12932 9027
rect 2973 8925 3007 8959
rect 7941 8925 7975 8959
rect 8125 8925 8159 8959
rect 10333 8925 10367 8959
rect 7573 8857 7607 8891
rect 8861 8857 8895 8891
rect 11437 8857 11471 8891
rect 2513 8789 2547 8823
rect 9781 8789 9815 8823
rect 3893 8585 3927 8619
rect 5273 8585 5307 8619
rect 6929 8585 6963 8619
rect 8217 8585 8251 8619
rect 9873 8585 9907 8619
rect 11161 8585 11195 8619
rect 12909 8585 12943 8619
rect 5089 8517 5123 8551
rect 8953 8517 8987 8551
rect 11437 8517 11471 8551
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 7481 8449 7515 8483
rect 7849 8449 7883 8483
rect 8677 8449 8711 8483
rect 1961 8381 1995 8415
rect 2217 8381 2251 8415
rect 7205 8381 7239 8415
rect 9229 8381 9263 8415
rect 11253 8381 11287 8415
rect 11805 8381 11839 8415
rect 13093 8381 13127 8415
rect 13645 8381 13679 8415
rect 6653 8313 6687 8347
rect 7389 8313 7423 8347
rect 9413 8313 9447 8347
rect 9505 8313 9539 8347
rect 1869 8245 1903 8279
rect 3341 8245 3375 8279
rect 4353 8245 4387 8279
rect 4721 8245 4755 8279
rect 5733 8245 5767 8279
rect 10241 8245 10275 8279
rect 10609 8245 10643 8279
rect 12265 8245 12299 8279
rect 13277 8245 13311 8279
rect 1961 8041 1995 8075
rect 2973 8041 3007 8075
rect 3525 8041 3559 8075
rect 6377 8041 6411 8075
rect 6929 8041 6963 8075
rect 7573 8041 7607 8075
rect 9137 8041 9171 8075
rect 11437 8041 11471 8075
rect 2237 7973 2271 8007
rect 5264 7973 5298 8007
rect 8401 7973 8435 8007
rect 8585 7973 8619 8007
rect 8677 7973 8711 8007
rect 10241 7973 10275 8007
rect 10333 7973 10367 8007
rect 3065 7905 3099 7939
rect 7941 7905 7975 7939
rect 10057 7905 10091 7939
rect 12072 7905 12106 7939
rect 2973 7837 3007 7871
rect 4997 7837 5031 7871
rect 11805 7837 11839 7871
rect 9781 7769 9815 7803
rect 13185 7769 13219 7803
rect 2513 7701 2547 7735
rect 4353 7701 4387 7735
rect 8125 7701 8159 7735
rect 9505 7701 9539 7735
rect 10701 7701 10735 7735
rect 2513 7497 2547 7531
rect 3157 7497 3191 7531
rect 4353 7497 4387 7531
rect 8769 7497 8803 7531
rect 9137 7429 9171 7463
rect 9781 7429 9815 7463
rect 1593 7361 1627 7395
rect 4813 7361 4847 7395
rect 1409 7293 1443 7327
rect 3801 7293 3835 7327
rect 4905 7293 4939 7327
rect 5641 7293 5675 7327
rect 6837 7293 6871 7327
rect 9873 7293 9907 7327
rect 11805 7293 11839 7327
rect 12725 7293 12759 7327
rect 4077 7225 4111 7259
rect 4813 7225 4847 7259
rect 7082 7225 7116 7259
rect 10118 7225 10152 7259
rect 13277 7225 13311 7259
rect 2789 7157 2823 7191
rect 5273 7157 5307 7191
rect 6561 7157 6595 7191
rect 8217 7157 8251 7191
rect 11253 7157 11287 7191
rect 12265 7157 12299 7191
rect 12909 7157 12943 7191
rect 5457 6953 5491 6987
rect 6929 6953 6963 6987
rect 8493 6953 8527 6987
rect 9965 6953 9999 6987
rect 9505 6885 9539 6919
rect 10578 6885 10612 6919
rect 1409 6817 1443 6851
rect 2697 6817 2731 6851
rect 3801 6817 3835 6851
rect 4344 6817 4378 6851
rect 7380 6817 7414 6851
rect 9045 6817 9079 6851
rect 12817 6817 12851 6851
rect 1593 6749 1627 6783
rect 2881 6749 2915 6783
rect 4077 6749 4111 6783
rect 7113 6749 7147 6783
rect 10333 6749 10367 6783
rect 2237 6613 2271 6647
rect 2513 6613 2547 6647
rect 3433 6613 3467 6647
rect 11713 6613 11747 6647
rect 13001 6613 13035 6647
rect 8401 6409 8435 6443
rect 10701 6409 10735 6443
rect 11897 6409 11931 6443
rect 13369 6409 13403 6443
rect 9045 6341 9079 6375
rect 8861 6273 8895 6307
rect 1961 6205 1995 6239
rect 2228 6205 2262 6239
rect 7849 6205 7883 6239
rect 9321 6205 9355 6239
rect 9597 6205 9631 6239
rect 11253 6205 11287 6239
rect 12449 6205 12483 6239
rect 13001 6205 13035 6239
rect 1869 6137 1903 6171
rect 4445 6137 4479 6171
rect 9459 6137 9493 6171
rect 3341 6069 3375 6103
rect 4169 6069 4203 6103
rect 7113 6069 7147 6103
rect 7573 6069 7607 6103
rect 8033 6069 8067 6103
rect 10333 6069 10367 6103
rect 11437 6069 11471 6103
rect 12633 6069 12667 6103
rect 2329 5865 2363 5899
rect 8953 5865 8987 5899
rect 10241 5865 10275 5899
rect 12909 5865 12943 5899
rect 8309 5797 8343 5831
rect 10057 5797 10091 5831
rect 10333 5797 10367 5831
rect 11796 5797 11830 5831
rect 2145 5729 2179 5763
rect 4537 5729 4571 5763
rect 6653 5729 6687 5763
rect 8125 5729 8159 5763
rect 2421 5661 2455 5695
rect 4077 5661 4111 5695
rect 7665 5661 7699 5695
rect 8401 5661 8435 5695
rect 11529 5661 11563 5695
rect 1869 5593 1903 5627
rect 3801 5593 3835 5627
rect 9781 5593 9815 5627
rect 1685 5525 1719 5559
rect 2881 5525 2915 5559
rect 3433 5525 3467 5559
rect 6837 5525 6871 5559
rect 7849 5525 7883 5559
rect 10701 5525 10735 5559
rect 1777 5321 1811 5355
rect 1961 5321 1995 5355
rect 6653 5321 6687 5355
rect 7113 5321 7147 5355
rect 7481 5321 7515 5355
rect 10885 5321 10919 5355
rect 11989 5321 12023 5355
rect 3525 5253 3559 5287
rect 4813 5253 4847 5287
rect 7757 5253 7791 5287
rect 9965 5253 9999 5287
rect 2421 5185 2455 5219
rect 3985 5185 4019 5219
rect 10425 5185 10459 5219
rect 2513 5117 2547 5151
rect 5733 5117 5767 5151
rect 8033 5117 8067 5151
rect 8677 5117 8711 5151
rect 9413 5117 9447 5151
rect 9781 5117 9815 5151
rect 10517 5117 10551 5151
rect 12449 5117 12483 5151
rect 13001 5117 13035 5151
rect 4077 5049 4111 5083
rect 8217 5049 8251 5083
rect 8309 5049 8343 5083
rect 10425 5049 10459 5083
rect 2421 4981 2455 5015
rect 2881 4981 2915 5015
rect 3341 4981 3375 5015
rect 3985 4981 4019 5015
rect 4445 4981 4479 5015
rect 5273 4981 5307 5015
rect 5641 4981 5675 5015
rect 6285 4981 6319 5015
rect 11529 4981 11563 5015
rect 12633 4981 12667 5015
rect 1961 4777 1995 4811
rect 2697 4777 2731 4811
rect 3525 4777 3559 4811
rect 6009 4777 6043 4811
rect 6837 4777 6871 4811
rect 7481 4777 7515 4811
rect 7941 4777 7975 4811
rect 9873 4777 9907 4811
rect 10977 4777 11011 4811
rect 2789 4709 2823 4743
rect 4629 4709 4663 4743
rect 7573 4709 7607 4743
rect 10793 4709 10827 4743
rect 4445 4641 4479 4675
rect 5825 4641 5859 4675
rect 8493 4641 8527 4675
rect 10333 4641 10367 4675
rect 11989 4641 12023 4675
rect 13093 4641 13127 4675
rect 2697 4573 2731 4607
rect 4721 4573 4755 4607
rect 7481 4573 7515 4607
rect 9505 4573 9539 4607
rect 11069 4573 11103 4607
rect 2237 4505 2271 4539
rect 4169 4505 4203 4539
rect 5733 4505 5767 4539
rect 8401 4505 8435 4539
rect 10517 4505 10551 4539
rect 3801 4437 3835 4471
rect 5273 4437 5307 4471
rect 6469 4437 6503 4471
rect 7021 4437 7055 4471
rect 8677 4437 8711 4471
rect 9137 4437 9171 4471
rect 12173 4437 12207 4471
rect 13277 4437 13311 4471
rect 3709 4233 3743 4267
rect 4353 4233 4387 4267
rect 5273 4233 5307 4267
rect 6193 4233 6227 4267
rect 7849 4233 7883 4267
rect 8309 4233 8343 4267
rect 9689 4233 9723 4267
rect 10977 4233 11011 4267
rect 11989 4233 12023 4267
rect 13185 4233 13219 4267
rect 6653 4165 6687 4199
rect 5641 4097 5675 4131
rect 6911 4097 6945 4131
rect 7481 4097 7515 4131
rect 8953 4097 8987 4131
rect 10057 4165 10091 4199
rect 10609 4097 10643 4131
rect 11345 4097 11379 4131
rect 2329 4029 2363 4063
rect 8475 4029 8509 4063
rect 9689 4029 9723 4063
rect 12449 4029 12483 4063
rect 1869 3961 1903 3995
rect 2574 3961 2608 3995
rect 5825 3961 5859 3995
rect 7205 3961 7239 3995
rect 8953 3961 8987 3995
rect 9045 3961 9079 3995
rect 10333 3961 10367 3995
rect 13553 3961 13587 3995
rect 2237 3893 2271 3927
rect 4721 3893 4755 3927
rect 4997 3893 5031 3927
rect 5733 3893 5767 3927
rect 7389 3893 7423 3927
rect 9505 3893 9539 3927
rect 9781 3893 9815 3927
rect 10517 3893 10551 3927
rect 12633 3893 12667 3927
rect 1961 3689 1995 3723
rect 7573 3689 7607 3723
rect 8217 3689 8251 3723
rect 8769 3689 8803 3723
rect 11621 3689 11655 3723
rect 2973 3621 3007 3655
rect 5448 3621 5482 3655
rect 7113 3621 7147 3655
rect 8033 3621 8067 3655
rect 9045 3621 9079 3655
rect 9413 3621 9447 3655
rect 10057 3621 10091 3655
rect 10486 3621 10520 3655
rect 13277 3621 13311 3655
rect 4077 3553 4111 3587
rect 4629 3553 4663 3587
rect 5181 3553 5215 3587
rect 8309 3553 8343 3587
rect 13093 3553 13127 3587
rect 13369 3553 13403 3587
rect 2973 3485 3007 3519
rect 3065 3485 3099 3519
rect 10241 3485 10275 3519
rect 12449 3485 12483 3519
rect 2513 3417 2547 3451
rect 7757 3417 7791 3451
rect 12817 3417 12851 3451
rect 2329 3349 2363 3383
rect 3433 3349 3467 3383
rect 3893 3349 3927 3383
rect 4261 3349 4295 3383
rect 4997 3349 5031 3383
rect 6561 3349 6595 3383
rect 2789 3145 2823 3179
rect 3709 3145 3743 3179
rect 6929 3145 6963 3179
rect 7941 3145 7975 3179
rect 10057 3145 10091 3179
rect 10977 3145 11011 3179
rect 13369 3145 13403 3179
rect 6285 3077 6319 3111
rect 8493 3077 8527 3111
rect 12173 3077 12207 3111
rect 13737 3077 13771 3111
rect 1593 3009 1627 3043
rect 2605 3009 2639 3043
rect 3157 3009 3191 3043
rect 6653 3009 6687 3043
rect 7481 3009 7515 3043
rect 8677 3009 8711 3043
rect 1409 2941 1443 2975
rect 4077 2941 4111 2975
rect 4261 2941 4295 2975
rect 4528 2941 4562 2975
rect 7205 2941 7239 2975
rect 11161 2941 11195 2975
rect 11713 2941 11747 2975
rect 12449 2941 12483 2975
rect 13001 2941 13035 2975
rect 2237 2873 2271 2907
rect 3249 2873 3283 2907
rect 3341 2873 3375 2907
rect 7389 2873 7423 2907
rect 8922 2873 8956 2907
rect 5641 2805 5675 2839
rect 10609 2805 10643 2839
rect 11345 2805 11379 2839
rect 12633 2805 12667 2839
rect 5549 2601 5583 2635
rect 6377 2601 6411 2635
rect 7481 2601 7515 2635
rect 7941 2601 7975 2635
rect 10425 2601 10459 2635
rect 11069 2601 11103 2635
rect 11529 2601 11563 2635
rect 2973 2533 3007 2567
rect 3525 2533 3559 2567
rect 4414 2533 4448 2567
rect 11161 2533 11195 2567
rect 2789 2465 2823 2499
rect 3893 2465 3927 2499
rect 4169 2465 4203 2499
rect 8493 2465 8527 2499
rect 9045 2465 9079 2499
rect 10057 2465 10091 2499
rect 10885 2465 10919 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 3065 2397 3099 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 7573 2397 7607 2431
rect 8401 2397 8435 2431
rect 9413 2397 9447 2431
rect 2237 2329 2271 2363
rect 2513 2329 2547 2363
rect 7021 2329 7055 2363
rect 8677 2329 8711 2363
rect 10609 2329 10643 2363
rect 1961 2261 1995 2295
rect 12817 2261 12851 2295
<< metal1 >>
rect 5534 37680 5540 37732
rect 5592 37720 5598 37732
rect 6362 37720 6368 37732
rect 5592 37692 6368 37720
rect 5592 37680 5598 37692
rect 6362 37680 6368 37692
rect 6420 37680 6426 37732
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 11333 36907 11391 36913
rect 11333 36873 11345 36907
rect 11379 36904 11391 36907
rect 12342 36904 12348 36916
rect 11379 36876 12348 36904
rect 11379 36873 11391 36876
rect 11333 36867 11391 36873
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 11149 36703 11207 36709
rect 11149 36669 11161 36703
rect 11195 36700 11207 36703
rect 11330 36700 11336 36712
rect 11195 36672 11336 36700
rect 11195 36669 11207 36672
rect 11149 36663 11207 36669
rect 11330 36660 11336 36672
rect 11388 36700 11394 36712
rect 11701 36703 11759 36709
rect 11701 36700 11713 36703
rect 11388 36672 11713 36700
rect 11388 36660 11394 36672
rect 11701 36669 11713 36672
rect 11747 36669 11759 36703
rect 11701 36663 11759 36669
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 10962 36360 10968 36372
rect 10923 36332 10968 36360
rect 10962 36320 10968 36332
rect 11020 36320 11026 36372
rect 12069 36363 12127 36369
rect 12069 36329 12081 36363
rect 12115 36360 12127 36363
rect 13446 36360 13452 36372
rect 12115 36332 13452 36360
rect 12115 36329 12127 36332
rect 12069 36323 12127 36329
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 10778 36224 10784 36236
rect 10739 36196 10784 36224
rect 10778 36184 10784 36196
rect 10836 36184 10842 36236
rect 11885 36227 11943 36233
rect 11885 36193 11897 36227
rect 11931 36224 11943 36227
rect 12250 36224 12256 36236
rect 11931 36196 12256 36224
rect 11931 36193 11943 36196
rect 11885 36187 11943 36193
rect 12250 36184 12256 36196
rect 12308 36184 12314 36236
rect 4338 36020 4344 36032
rect 4251 35992 4344 36020
rect 4338 35980 4344 35992
rect 4396 36020 4402 36032
rect 4614 36020 4620 36032
rect 4396 35992 4620 36020
rect 4396 35980 4402 35992
rect 4614 35980 4620 35992
rect 4672 35980 4678 36032
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 8021 35819 8079 35825
rect 8021 35785 8033 35819
rect 8067 35816 8079 35819
rect 8202 35816 8208 35828
rect 8067 35788 8208 35816
rect 8067 35785 8079 35788
rect 8021 35779 8079 35785
rect 8202 35776 8208 35788
rect 8260 35776 8266 35828
rect 9125 35819 9183 35825
rect 9125 35785 9137 35819
rect 9171 35816 9183 35819
rect 9306 35816 9312 35828
rect 9171 35788 9312 35816
rect 9171 35785 9183 35788
rect 9125 35779 9183 35785
rect 9306 35776 9312 35788
rect 9364 35776 9370 35828
rect 10229 35819 10287 35825
rect 10229 35785 10241 35819
rect 10275 35816 10287 35819
rect 10686 35816 10692 35828
rect 10275 35788 10692 35816
rect 10275 35785 10287 35788
rect 10229 35779 10287 35785
rect 10686 35776 10692 35788
rect 10744 35776 10750 35828
rect 11054 35776 11060 35828
rect 11112 35816 11118 35828
rect 11333 35819 11391 35825
rect 11333 35816 11345 35819
rect 11112 35788 11345 35816
rect 11112 35776 11118 35788
rect 11333 35785 11345 35788
rect 11379 35785 11391 35819
rect 11333 35779 11391 35785
rect 12621 35819 12679 35825
rect 12621 35785 12633 35819
rect 12667 35816 12679 35819
rect 13722 35816 13728 35828
rect 12667 35788 13728 35816
rect 12667 35785 12679 35788
rect 12621 35779 12679 35785
rect 13722 35776 13728 35788
rect 13780 35776 13786 35828
rect 3970 35708 3976 35760
rect 4028 35748 4034 35760
rect 4065 35751 4123 35757
rect 4065 35748 4077 35751
rect 4028 35720 4077 35748
rect 4028 35708 4034 35720
rect 4065 35717 4077 35720
rect 4111 35717 4123 35751
rect 4065 35711 4123 35717
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 3513 35683 3571 35689
rect 3513 35649 3525 35683
rect 3559 35680 3571 35683
rect 4522 35680 4528 35692
rect 3559 35652 4528 35680
rect 3559 35649 3571 35652
rect 3513 35643 3571 35649
rect 4522 35640 4528 35652
rect 4580 35640 4586 35692
rect 4614 35640 4620 35692
rect 4672 35680 4678 35692
rect 4672 35652 4717 35680
rect 4672 35640 4678 35652
rect 1397 35615 1455 35621
rect 1397 35581 1409 35615
rect 1443 35612 1455 35615
rect 1762 35612 1768 35624
rect 1443 35584 1768 35612
rect 1443 35581 1455 35584
rect 1397 35575 1455 35581
rect 1762 35572 1768 35584
rect 1820 35572 1826 35624
rect 7837 35615 7895 35621
rect 7837 35581 7849 35615
rect 7883 35612 7895 35615
rect 8386 35612 8392 35624
rect 7883 35584 8392 35612
rect 7883 35581 7895 35584
rect 7837 35575 7895 35581
rect 8386 35572 8392 35584
rect 8444 35572 8450 35624
rect 8570 35572 8576 35624
rect 8628 35612 8634 35624
rect 8941 35615 8999 35621
rect 8941 35612 8953 35615
rect 8628 35584 8953 35612
rect 8628 35572 8634 35584
rect 8941 35581 8953 35584
rect 8987 35612 8999 35615
rect 9493 35615 9551 35621
rect 9493 35612 9505 35615
rect 8987 35584 9505 35612
rect 8987 35581 8999 35584
rect 8941 35575 8999 35581
rect 9493 35581 9505 35584
rect 9539 35581 9551 35615
rect 10045 35615 10103 35621
rect 10045 35612 10057 35615
rect 9493 35575 9551 35581
rect 9876 35584 10057 35612
rect 9876 35488 9904 35584
rect 10045 35581 10057 35584
rect 10091 35581 10103 35615
rect 11146 35612 11152 35624
rect 11107 35584 11152 35612
rect 10045 35575 10103 35581
rect 11146 35572 11152 35584
rect 11204 35572 11210 35624
rect 12437 35615 12495 35621
rect 12437 35581 12449 35615
rect 12483 35612 12495 35615
rect 12483 35584 13124 35612
rect 12483 35581 12495 35584
rect 12437 35575 12495 35581
rect 2222 35476 2228 35488
rect 2183 35448 2228 35476
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 3881 35479 3939 35485
rect 3881 35445 3893 35479
rect 3927 35476 3939 35479
rect 4525 35479 4583 35485
rect 4525 35476 4537 35479
rect 3927 35448 4537 35476
rect 3927 35445 3939 35448
rect 3881 35439 3939 35445
rect 4525 35445 4537 35448
rect 4571 35476 4583 35479
rect 4798 35476 4804 35488
rect 4571 35448 4804 35476
rect 4571 35445 4583 35448
rect 4525 35439 4583 35445
rect 4798 35436 4804 35448
rect 4856 35476 4862 35488
rect 4982 35476 4988 35488
rect 4856 35448 4988 35476
rect 4856 35436 4862 35448
rect 4982 35436 4988 35448
rect 5040 35436 5046 35488
rect 9858 35476 9864 35488
rect 9819 35448 9864 35476
rect 9858 35436 9864 35448
rect 9916 35436 9922 35488
rect 10686 35436 10692 35488
rect 10744 35476 10750 35488
rect 10781 35479 10839 35485
rect 10781 35476 10793 35479
rect 10744 35448 10793 35476
rect 10744 35436 10750 35448
rect 10781 35445 10793 35448
rect 10827 35445 10839 35479
rect 10781 35439 10839 35445
rect 11977 35479 12035 35485
rect 11977 35445 11989 35479
rect 12023 35476 12035 35479
rect 12250 35476 12256 35488
rect 12023 35448 12256 35476
rect 12023 35445 12035 35448
rect 11977 35439 12035 35445
rect 12250 35436 12256 35448
rect 12308 35436 12314 35488
rect 13096 35485 13124 35584
rect 13081 35479 13139 35485
rect 13081 35445 13093 35479
rect 13127 35476 13139 35479
rect 13262 35476 13268 35488
rect 13127 35448 13268 35476
rect 13127 35445 13139 35448
rect 13081 35439 13139 35445
rect 13262 35436 13268 35448
rect 13320 35436 13326 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 7653 35275 7711 35281
rect 7653 35241 7665 35275
rect 7699 35272 7711 35275
rect 7926 35272 7932 35284
rect 7699 35244 7932 35272
rect 7699 35241 7711 35244
rect 7653 35235 7711 35241
rect 7926 35232 7932 35244
rect 7984 35232 7990 35284
rect 9490 35232 9496 35284
rect 9548 35272 9554 35284
rect 9861 35275 9919 35281
rect 9861 35272 9873 35275
rect 9548 35244 9873 35272
rect 9548 35232 9554 35244
rect 9861 35241 9873 35244
rect 9907 35241 9919 35275
rect 9861 35235 9919 35241
rect 9950 35232 9956 35284
rect 10008 35272 10014 35284
rect 10965 35275 11023 35281
rect 10965 35272 10977 35275
rect 10008 35244 10977 35272
rect 10008 35232 10014 35244
rect 10965 35241 10977 35244
rect 11011 35241 11023 35275
rect 10965 35235 11023 35241
rect 11146 35232 11152 35284
rect 11204 35272 11210 35284
rect 11333 35275 11391 35281
rect 11333 35272 11345 35275
rect 11204 35244 11345 35272
rect 11204 35232 11210 35244
rect 11333 35241 11345 35244
rect 11379 35241 11391 35275
rect 11333 35235 11391 35241
rect 11514 35232 11520 35284
rect 11572 35272 11578 35284
rect 12069 35275 12127 35281
rect 12069 35272 12081 35275
rect 11572 35244 12081 35272
rect 11572 35232 11578 35244
rect 12069 35241 12081 35244
rect 12115 35241 12127 35275
rect 13354 35272 13360 35284
rect 13315 35244 13360 35272
rect 12069 35235 12127 35241
rect 13354 35232 13360 35244
rect 13412 35232 13418 35284
rect 2041 35207 2099 35213
rect 2041 35173 2053 35207
rect 2087 35204 2099 35207
rect 2498 35204 2504 35216
rect 2087 35176 2504 35204
rect 2087 35173 2099 35176
rect 2041 35167 2099 35173
rect 2498 35164 2504 35176
rect 2556 35204 2562 35216
rect 2685 35207 2743 35213
rect 2685 35204 2697 35207
rect 2556 35176 2697 35204
rect 2556 35164 2562 35176
rect 2685 35173 2697 35176
rect 2731 35173 2743 35207
rect 2685 35167 2743 35173
rect 5252 35207 5310 35213
rect 5252 35173 5264 35207
rect 5298 35204 5310 35207
rect 5442 35204 5448 35216
rect 5298 35176 5448 35204
rect 5298 35173 5310 35176
rect 5252 35167 5310 35173
rect 5442 35164 5448 35176
rect 5500 35164 5506 35216
rect 7469 35139 7527 35145
rect 7469 35105 7481 35139
rect 7515 35136 7527 35139
rect 7834 35136 7840 35148
rect 7515 35108 7840 35136
rect 7515 35105 7527 35108
rect 7469 35099 7527 35105
rect 7834 35096 7840 35108
rect 7892 35096 7898 35148
rect 9677 35139 9735 35145
rect 9677 35105 9689 35139
rect 9723 35136 9735 35139
rect 9766 35136 9772 35148
rect 9723 35108 9772 35136
rect 9723 35105 9735 35108
rect 9677 35099 9735 35105
rect 9766 35096 9772 35108
rect 9824 35096 9830 35148
rect 10778 35136 10784 35148
rect 10739 35108 10784 35136
rect 10778 35096 10784 35108
rect 10836 35096 10842 35148
rect 11885 35139 11943 35145
rect 11885 35105 11897 35139
rect 11931 35136 11943 35139
rect 12066 35136 12072 35148
rect 11931 35108 12072 35136
rect 11931 35105 11943 35108
rect 11885 35099 11943 35105
rect 12066 35096 12072 35108
rect 12124 35096 12130 35148
rect 13170 35136 13176 35148
rect 13131 35108 13176 35136
rect 13170 35096 13176 35108
rect 13228 35096 13234 35148
rect 2222 35028 2228 35080
rect 2280 35068 2286 35080
rect 2406 35068 2412 35080
rect 2280 35040 2412 35068
rect 2280 35028 2286 35040
rect 2406 35028 2412 35040
rect 2464 35068 2470 35080
rect 2593 35071 2651 35077
rect 2593 35068 2605 35071
rect 2464 35040 2605 35068
rect 2464 35028 2470 35040
rect 2593 35037 2605 35040
rect 2639 35037 2651 35071
rect 2593 35031 2651 35037
rect 2777 35071 2835 35077
rect 2777 35037 2789 35071
rect 2823 35068 2835 35071
rect 2958 35068 2964 35080
rect 2823 35040 2964 35068
rect 2823 35037 2835 35040
rect 2777 35031 2835 35037
rect 2958 35028 2964 35040
rect 3016 35028 3022 35080
rect 4890 35028 4896 35080
rect 4948 35068 4954 35080
rect 4985 35071 5043 35077
rect 4985 35068 4997 35071
rect 4948 35040 4997 35068
rect 4948 35028 4954 35040
rect 4985 35037 4997 35040
rect 5031 35037 5043 35071
rect 4985 35031 5043 35037
rect 1673 34935 1731 34941
rect 1673 34901 1685 34935
rect 1719 34932 1731 34935
rect 1762 34932 1768 34944
rect 1719 34904 1768 34932
rect 1719 34901 1731 34904
rect 1673 34895 1731 34901
rect 1762 34892 1768 34904
rect 1820 34892 1826 34944
rect 2222 34932 2228 34944
rect 2183 34904 2228 34932
rect 2222 34892 2228 34904
rect 2280 34892 2286 34944
rect 3234 34932 3240 34944
rect 3195 34904 3240 34932
rect 3234 34892 3240 34904
rect 3292 34892 3298 34944
rect 4341 34935 4399 34941
rect 4341 34901 4353 34935
rect 4387 34932 4399 34935
rect 4614 34932 4620 34944
rect 4387 34904 4620 34932
rect 4387 34901 4399 34904
rect 4341 34895 4399 34901
rect 4614 34892 4620 34904
rect 4672 34932 4678 34944
rect 6365 34935 6423 34941
rect 6365 34932 6377 34935
rect 4672 34904 6377 34932
rect 4672 34892 4678 34904
rect 6365 34901 6377 34904
rect 6411 34901 6423 34935
rect 7006 34932 7012 34944
rect 6967 34904 7012 34932
rect 6365 34895 6423 34901
rect 7006 34892 7012 34904
rect 7064 34892 7070 34944
rect 8481 34935 8539 34941
rect 8481 34901 8493 34935
rect 8527 34932 8539 34935
rect 8846 34932 8852 34944
rect 8527 34904 8852 34932
rect 8527 34901 8539 34904
rect 8481 34895 8539 34901
rect 8846 34892 8852 34904
rect 8904 34892 8910 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 2498 34728 2504 34740
rect 2459 34700 2504 34728
rect 2498 34688 2504 34700
rect 2556 34688 2562 34740
rect 3234 34688 3240 34740
rect 3292 34728 3298 34740
rect 4065 34731 4123 34737
rect 4065 34728 4077 34731
rect 3292 34700 4077 34728
rect 3292 34688 3298 34700
rect 4065 34697 4077 34700
rect 4111 34697 4123 34731
rect 7834 34728 7840 34740
rect 7795 34700 7840 34728
rect 4065 34691 4123 34697
rect 7834 34688 7840 34700
rect 7892 34688 7898 34740
rect 8754 34688 8760 34740
rect 8812 34728 8818 34740
rect 10137 34731 10195 34737
rect 10137 34728 10149 34731
rect 8812 34700 10149 34728
rect 8812 34688 8818 34700
rect 10137 34697 10149 34700
rect 10183 34697 10195 34731
rect 10137 34691 10195 34697
rect 10318 34688 10324 34740
rect 10376 34728 10382 34740
rect 11241 34731 11299 34737
rect 11241 34728 11253 34731
rect 10376 34700 11253 34728
rect 10376 34688 10382 34700
rect 11241 34697 11253 34700
rect 11287 34697 11299 34731
rect 13630 34728 13636 34740
rect 13591 34700 13636 34728
rect 11241 34691 11299 34697
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 5074 34660 5080 34672
rect 4448 34632 5080 34660
rect 2317 34595 2375 34601
rect 2317 34561 2329 34595
rect 2363 34592 2375 34595
rect 2961 34595 3019 34601
rect 2961 34592 2973 34595
rect 2363 34564 2973 34592
rect 2363 34561 2375 34564
rect 2317 34555 2375 34561
rect 2961 34561 2973 34564
rect 3007 34592 3019 34595
rect 3142 34592 3148 34604
rect 3007 34564 3148 34592
rect 3007 34561 3019 34564
rect 2961 34555 3019 34561
rect 3142 34552 3148 34564
rect 3200 34552 3206 34604
rect 3418 34552 3424 34604
rect 3476 34592 3482 34604
rect 4448 34601 4476 34632
rect 5074 34620 5080 34632
rect 5132 34620 5138 34672
rect 6730 34620 6736 34672
rect 6788 34660 6794 34672
rect 6917 34663 6975 34669
rect 6917 34660 6929 34663
rect 6788 34632 6929 34660
rect 6788 34620 6794 34632
rect 6917 34629 6929 34632
rect 6963 34629 6975 34663
rect 8478 34660 8484 34672
rect 8439 34632 8484 34660
rect 6917 34623 6975 34629
rect 8478 34620 8484 34632
rect 8536 34620 8542 34672
rect 3513 34595 3571 34601
rect 3513 34592 3525 34595
rect 3476 34564 3525 34592
rect 3476 34552 3482 34564
rect 3513 34561 3525 34564
rect 3559 34592 3571 34595
rect 4433 34595 4491 34601
rect 4433 34592 4445 34595
rect 3559 34564 4445 34592
rect 3559 34561 3571 34564
rect 3513 34555 3571 34561
rect 4433 34561 4445 34564
rect 4479 34561 4491 34595
rect 4433 34555 4491 34561
rect 4522 34552 4528 34604
rect 4580 34592 4586 34604
rect 5537 34595 5595 34601
rect 5537 34592 5549 34595
rect 4580 34564 5549 34592
rect 4580 34552 4586 34564
rect 5537 34561 5549 34564
rect 5583 34561 5595 34595
rect 5537 34555 5595 34561
rect 8846 34552 8852 34604
rect 8904 34592 8910 34604
rect 9033 34595 9091 34601
rect 9033 34592 9045 34595
rect 8904 34564 9045 34592
rect 8904 34552 8910 34564
rect 9033 34561 9045 34564
rect 9079 34561 9091 34595
rect 10505 34595 10563 34601
rect 10505 34592 10517 34595
rect 9033 34555 9091 34561
rect 10152 34564 10517 34592
rect 10152 34536 10180 34564
rect 10505 34561 10517 34564
rect 10551 34561 10563 34595
rect 10505 34555 10563 34561
rect 1949 34527 2007 34533
rect 1949 34493 1961 34527
rect 1995 34524 2007 34527
rect 3053 34527 3111 34533
rect 3053 34524 3065 34527
rect 1995 34496 3065 34524
rect 1995 34493 2007 34496
rect 1949 34487 2007 34493
rect 3053 34493 3065 34496
rect 3099 34524 3111 34527
rect 4338 34524 4344 34536
rect 3099 34496 4344 34524
rect 3099 34493 3111 34496
rect 3053 34487 3111 34493
rect 4338 34484 4344 34496
rect 4396 34484 4402 34536
rect 4614 34524 4620 34536
rect 4575 34496 4620 34524
rect 4614 34484 4620 34496
rect 4672 34484 4678 34536
rect 5442 34524 5448 34536
rect 5403 34496 5448 34524
rect 5442 34484 5448 34496
rect 5500 34484 5506 34536
rect 6273 34527 6331 34533
rect 6273 34493 6285 34527
rect 6319 34524 6331 34527
rect 7098 34524 7104 34536
rect 6319 34496 7104 34524
rect 6319 34493 6331 34496
rect 6273 34487 6331 34493
rect 7098 34484 7104 34496
rect 7156 34524 7162 34536
rect 7193 34527 7251 34533
rect 7193 34524 7205 34527
rect 7156 34496 7205 34524
rect 7156 34484 7162 34496
rect 7193 34493 7205 34496
rect 7239 34493 7251 34527
rect 7193 34487 7251 34493
rect 8297 34527 8355 34533
rect 8297 34493 8309 34527
rect 8343 34524 8355 34527
rect 8570 34524 8576 34536
rect 8343 34496 8576 34524
rect 8343 34493 8355 34496
rect 8297 34487 8355 34493
rect 8570 34484 8576 34496
rect 8628 34524 8634 34536
rect 8757 34527 8815 34533
rect 8757 34524 8769 34527
rect 8628 34496 8769 34524
rect 8628 34484 8634 34496
rect 8757 34493 8769 34496
rect 8803 34493 8815 34527
rect 8757 34487 8815 34493
rect 9953 34527 10011 34533
rect 9953 34493 9965 34527
rect 9999 34524 10011 34527
rect 10134 34524 10140 34536
rect 9999 34496 10140 34524
rect 9999 34493 10011 34496
rect 9953 34487 10011 34493
rect 10134 34484 10140 34496
rect 10192 34484 10198 34536
rect 11057 34527 11115 34533
rect 11057 34493 11069 34527
rect 11103 34524 11115 34527
rect 11514 34524 11520 34536
rect 11103 34496 11520 34524
rect 11103 34493 11115 34496
rect 11057 34487 11115 34493
rect 11514 34484 11520 34496
rect 11572 34524 11578 34536
rect 11609 34527 11667 34533
rect 11609 34524 11621 34527
rect 11572 34496 11621 34524
rect 11572 34484 11578 34496
rect 11609 34493 11621 34496
rect 11655 34493 11667 34527
rect 12066 34524 12072 34536
rect 12027 34496 12072 34524
rect 11609 34487 11667 34493
rect 12066 34484 12072 34496
rect 12124 34484 12130 34536
rect 13170 34524 13176 34536
rect 13131 34496 13176 34524
rect 13170 34484 13176 34496
rect 13228 34484 13234 34536
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34493 13507 34527
rect 13449 34487 13507 34493
rect 7006 34416 7012 34468
rect 7064 34456 7070 34468
rect 7282 34456 7288 34468
rect 7064 34428 7288 34456
rect 7064 34416 7070 34428
rect 7282 34416 7288 34428
rect 7340 34456 7346 34468
rect 7377 34459 7435 34465
rect 7377 34456 7389 34459
rect 7340 34428 7389 34456
rect 7340 34416 7346 34428
rect 7377 34425 7389 34428
rect 7423 34425 7435 34459
rect 7377 34419 7435 34425
rect 7469 34459 7527 34465
rect 7469 34425 7481 34459
rect 7515 34425 7527 34459
rect 7469 34419 7527 34425
rect 2961 34391 3019 34397
rect 2961 34357 2973 34391
rect 3007 34388 3019 34391
rect 3234 34388 3240 34400
rect 3007 34360 3240 34388
rect 3007 34357 3019 34360
rect 2961 34351 3019 34357
rect 3234 34348 3240 34360
rect 3292 34348 3298 34400
rect 3881 34391 3939 34397
rect 3881 34357 3893 34391
rect 3927 34388 3939 34391
rect 4525 34391 4583 34397
rect 4525 34388 4537 34391
rect 3927 34360 4537 34388
rect 3927 34357 3939 34360
rect 3881 34351 3939 34357
rect 4525 34357 4537 34360
rect 4571 34388 4583 34391
rect 4798 34388 4804 34400
rect 4571 34360 4804 34388
rect 4571 34357 4583 34360
rect 4525 34351 4583 34357
rect 4798 34348 4804 34360
rect 4856 34348 4862 34400
rect 4890 34348 4896 34400
rect 4948 34388 4954 34400
rect 5077 34391 5135 34397
rect 5077 34388 5089 34391
rect 4948 34360 5089 34388
rect 4948 34348 4954 34360
rect 5077 34357 5089 34360
rect 5123 34388 5135 34391
rect 6086 34388 6092 34400
rect 5123 34360 6092 34388
rect 5123 34357 5135 34360
rect 5077 34351 5135 34357
rect 6086 34348 6092 34360
rect 6144 34348 6150 34400
rect 6641 34391 6699 34397
rect 6641 34357 6653 34391
rect 6687 34388 6699 34391
rect 6914 34388 6920 34400
rect 6687 34360 6920 34388
rect 6687 34357 6699 34360
rect 6641 34351 6699 34357
rect 6914 34348 6920 34360
rect 6972 34388 6978 34400
rect 7484 34388 7512 34419
rect 11238 34416 11244 34468
rect 11296 34456 11302 34468
rect 13464 34456 13492 34487
rect 14001 34459 14059 34465
rect 14001 34456 14013 34459
rect 11296 34428 14013 34456
rect 11296 34416 11302 34428
rect 14001 34425 14013 34428
rect 14047 34425 14059 34459
rect 14001 34419 14059 34425
rect 6972 34360 7512 34388
rect 6972 34348 6978 34360
rect 8846 34348 8852 34400
rect 8904 34388 8910 34400
rect 8941 34391 8999 34397
rect 8941 34388 8953 34391
rect 8904 34360 8953 34388
rect 8904 34348 8910 34360
rect 8941 34357 8953 34360
rect 8987 34357 8999 34391
rect 9766 34388 9772 34400
rect 9727 34360 9772 34388
rect 8941 34351 8999 34357
rect 9766 34348 9772 34360
rect 9824 34348 9830 34400
rect 10410 34348 10416 34400
rect 10468 34388 10474 34400
rect 10778 34388 10784 34400
rect 10468 34360 10784 34388
rect 10468 34348 10474 34360
rect 10778 34348 10784 34360
rect 10836 34388 10842 34400
rect 10873 34391 10931 34397
rect 10873 34388 10885 34391
rect 10836 34360 10885 34388
rect 10836 34348 10842 34360
rect 10873 34357 10885 34360
rect 10919 34357 10931 34391
rect 10873 34351 10931 34357
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 2222 34184 2228 34196
rect 2183 34156 2228 34184
rect 2222 34144 2228 34156
rect 2280 34184 2286 34196
rect 3421 34187 3479 34193
rect 3421 34184 3433 34187
rect 2280 34156 3433 34184
rect 2280 34144 2286 34156
rect 3421 34153 3433 34156
rect 3467 34153 3479 34187
rect 3421 34147 3479 34153
rect 5442 34144 5448 34196
rect 5500 34184 5506 34196
rect 8205 34187 8263 34193
rect 8205 34184 8217 34187
rect 5500 34156 8217 34184
rect 5500 34144 5506 34156
rect 8205 34153 8217 34156
rect 8251 34153 8263 34187
rect 8205 34147 8263 34153
rect 12897 34187 12955 34193
rect 12897 34153 12909 34187
rect 12943 34184 12955 34187
rect 14182 34184 14188 34196
rect 12943 34156 14188 34184
rect 12943 34153 12955 34156
rect 12897 34147 12955 34153
rect 14182 34144 14188 34156
rect 14240 34144 14246 34196
rect 2317 34119 2375 34125
rect 2317 34085 2329 34119
rect 2363 34116 2375 34119
rect 2774 34116 2780 34128
rect 2363 34088 2780 34116
rect 2363 34085 2375 34088
rect 2317 34079 2375 34085
rect 2774 34076 2780 34088
rect 2832 34076 2838 34128
rect 4614 34125 4620 34128
rect 4608 34116 4620 34125
rect 4575 34088 4620 34116
rect 4608 34079 4620 34088
rect 4614 34076 4620 34079
rect 4672 34076 4678 34128
rect 6914 34076 6920 34128
rect 6972 34116 6978 34128
rect 7070 34119 7128 34125
rect 7070 34116 7082 34119
rect 6972 34088 7082 34116
rect 6972 34076 6978 34088
rect 7070 34085 7082 34088
rect 7116 34085 7128 34119
rect 10226 34116 10232 34128
rect 7070 34079 7128 34085
rect 9692 34088 10232 34116
rect 2038 34048 2044 34060
rect 1999 34020 2044 34048
rect 2038 34008 2044 34020
rect 2096 34008 2102 34060
rect 4154 34008 4160 34060
rect 4212 34048 4218 34060
rect 4341 34051 4399 34057
rect 4341 34048 4353 34051
rect 4212 34020 4353 34048
rect 4212 34008 4218 34020
rect 4341 34017 4353 34020
rect 4387 34048 4399 34051
rect 4890 34048 4896 34060
rect 4387 34020 4896 34048
rect 4387 34017 4399 34020
rect 4341 34011 4399 34017
rect 4890 34008 4896 34020
rect 4948 34008 4954 34060
rect 9692 34057 9720 34088
rect 10226 34076 10232 34088
rect 10284 34076 10290 34128
rect 9950 34057 9956 34060
rect 9677 34051 9735 34057
rect 9677 34017 9689 34051
rect 9723 34017 9735 34051
rect 9677 34011 9735 34017
rect 9944 34011 9956 34057
rect 10008 34048 10014 34060
rect 12710 34048 12716 34060
rect 10008 34020 10044 34048
rect 12671 34020 12716 34048
rect 9950 34008 9956 34011
rect 10008 34008 10014 34020
rect 12710 34008 12716 34020
rect 12768 34008 12774 34060
rect 2777 33983 2835 33989
rect 2777 33949 2789 33983
rect 2823 33980 2835 33983
rect 2958 33980 2964 33992
rect 2823 33952 2964 33980
rect 2823 33949 2835 33952
rect 2777 33943 2835 33949
rect 2958 33940 2964 33952
rect 3016 33980 3022 33992
rect 3053 33983 3111 33989
rect 3053 33980 3065 33983
rect 3016 33952 3065 33980
rect 3016 33940 3022 33952
rect 3053 33949 3065 33952
rect 3099 33949 3111 33983
rect 3053 33943 3111 33949
rect 6086 33940 6092 33992
rect 6144 33980 6150 33992
rect 6825 33983 6883 33989
rect 6825 33980 6837 33983
rect 6144 33952 6837 33980
rect 6144 33940 6150 33952
rect 6825 33949 6837 33952
rect 6871 33949 6883 33983
rect 6825 33943 6883 33949
rect 1762 33912 1768 33924
rect 1723 33884 1768 33912
rect 1762 33872 1768 33884
rect 1820 33872 1826 33924
rect 4338 33804 4344 33856
rect 4396 33844 4402 33856
rect 5721 33847 5779 33853
rect 5721 33844 5733 33847
rect 4396 33816 5733 33844
rect 4396 33804 4402 33816
rect 5721 33813 5733 33816
rect 5767 33813 5779 33847
rect 8846 33844 8852 33856
rect 8759 33816 8852 33844
rect 5721 33807 5779 33813
rect 8846 33804 8852 33816
rect 8904 33844 8910 33856
rect 9490 33844 9496 33856
rect 8904 33816 9496 33844
rect 8904 33804 8910 33816
rect 9490 33804 9496 33816
rect 9548 33804 9554 33856
rect 10962 33804 10968 33856
rect 11020 33844 11026 33856
rect 11057 33847 11115 33853
rect 11057 33844 11069 33847
rect 11020 33816 11069 33844
rect 11020 33804 11026 33816
rect 11057 33813 11069 33816
rect 11103 33813 11115 33847
rect 11057 33807 11115 33813
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 2774 33600 2780 33652
rect 2832 33640 2838 33652
rect 2961 33643 3019 33649
rect 2961 33640 2973 33643
rect 2832 33612 2973 33640
rect 2832 33600 2838 33612
rect 2961 33609 2973 33612
rect 3007 33609 3019 33643
rect 7098 33640 7104 33652
rect 7059 33612 7104 33640
rect 2961 33603 3019 33609
rect 7098 33600 7104 33612
rect 7156 33600 7162 33652
rect 11241 33643 11299 33649
rect 11241 33609 11253 33643
rect 11287 33640 11299 33643
rect 11974 33640 11980 33652
rect 11287 33612 11980 33640
rect 11287 33609 11299 33612
rect 11241 33603 11299 33609
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 13630 33640 13636 33652
rect 13591 33612 13636 33640
rect 13630 33600 13636 33612
rect 13688 33600 13694 33652
rect 1581 33439 1639 33445
rect 1581 33405 1593 33439
rect 1627 33436 1639 33439
rect 1670 33436 1676 33448
rect 1627 33408 1676 33436
rect 1627 33405 1639 33408
rect 1581 33399 1639 33405
rect 1670 33396 1676 33408
rect 1728 33396 1734 33448
rect 3421 33439 3479 33445
rect 3421 33405 3433 33439
rect 3467 33436 3479 33439
rect 3605 33439 3663 33445
rect 3605 33436 3617 33439
rect 3467 33408 3617 33436
rect 3467 33405 3479 33408
rect 3421 33399 3479 33405
rect 3605 33405 3617 33408
rect 3651 33436 3663 33439
rect 3973 33439 4031 33445
rect 3973 33436 3985 33439
rect 3651 33408 3985 33436
rect 3651 33405 3663 33408
rect 3605 33399 3663 33405
rect 3973 33405 3985 33408
rect 4019 33436 4031 33439
rect 4065 33439 4123 33445
rect 4065 33436 4077 33439
rect 4019 33408 4077 33436
rect 4019 33405 4031 33408
rect 3973 33399 4031 33405
rect 4065 33405 4077 33408
rect 4111 33436 4123 33439
rect 4154 33436 4160 33448
rect 4111 33408 4160 33436
rect 4111 33405 4123 33408
rect 4065 33399 4123 33405
rect 4154 33396 4160 33408
rect 4212 33396 4218 33448
rect 4338 33445 4344 33448
rect 4332 33436 4344 33445
rect 4299 33408 4344 33436
rect 4332 33399 4344 33408
rect 4338 33396 4344 33399
rect 4396 33396 4402 33448
rect 6914 33396 6920 33448
rect 6972 33436 6978 33448
rect 8021 33439 8079 33445
rect 8021 33436 8033 33439
rect 6972 33408 8033 33436
rect 6972 33396 6978 33408
rect 8021 33405 8033 33408
rect 8067 33436 8079 33439
rect 8202 33436 8208 33448
rect 8067 33408 8208 33436
rect 8067 33405 8079 33408
rect 8021 33399 8079 33405
rect 8202 33396 8208 33408
rect 8260 33396 8266 33448
rect 8478 33436 8484 33448
rect 8391 33408 8484 33436
rect 8478 33396 8484 33408
rect 8536 33436 8542 33448
rect 8573 33439 8631 33445
rect 8573 33436 8585 33439
rect 8536 33408 8585 33436
rect 8536 33396 8542 33408
rect 8573 33405 8585 33408
rect 8619 33436 8631 33439
rect 10226 33436 10232 33448
rect 8619 33408 10232 33436
rect 8619 33405 8631 33408
rect 8573 33399 8631 33405
rect 10226 33396 10232 33408
rect 10284 33396 10290 33448
rect 11057 33439 11115 33445
rect 11057 33405 11069 33439
rect 11103 33436 11115 33439
rect 13446 33436 13452 33448
rect 11103 33408 11468 33436
rect 13359 33408 13452 33436
rect 11103 33405 11115 33408
rect 11057 33399 11115 33405
rect 1848 33371 1906 33377
rect 1848 33337 1860 33371
rect 1894 33368 1906 33371
rect 2958 33368 2964 33380
rect 1894 33340 2964 33368
rect 1894 33337 1906 33340
rect 1848 33331 1906 33337
rect 2958 33328 2964 33340
rect 3016 33368 3022 33380
rect 3016 33340 4016 33368
rect 3016 33328 3022 33340
rect 1670 33260 1676 33312
rect 1728 33300 1734 33312
rect 3421 33303 3479 33309
rect 3421 33300 3433 33303
rect 1728 33272 3433 33300
rect 1728 33260 1734 33272
rect 3421 33269 3433 33272
rect 3467 33269 3479 33303
rect 3988 33300 4016 33340
rect 7098 33328 7104 33380
rect 7156 33368 7162 33380
rect 7377 33371 7435 33377
rect 7377 33368 7389 33371
rect 7156 33340 7389 33368
rect 7156 33328 7162 33340
rect 7377 33337 7389 33340
rect 7423 33337 7435 33371
rect 7558 33368 7564 33380
rect 7519 33340 7564 33368
rect 7377 33331 7435 33337
rect 7558 33328 7564 33340
rect 7616 33328 7622 33380
rect 7650 33328 7656 33380
rect 7708 33368 7714 33380
rect 8846 33377 8852 33380
rect 8840 33368 8852 33377
rect 7708 33340 7753 33368
rect 8807 33340 8852 33368
rect 7708 33328 7714 33340
rect 8840 33331 8852 33340
rect 8846 33328 8852 33331
rect 8904 33328 8910 33380
rect 5445 33303 5503 33309
rect 5445 33300 5457 33303
rect 3988 33272 5457 33300
rect 3421 33263 3479 33269
rect 5445 33269 5457 33272
rect 5491 33269 5503 33303
rect 5445 33263 5503 33269
rect 6086 33260 6092 33312
rect 6144 33300 6150 33312
rect 6181 33303 6239 33309
rect 6181 33300 6193 33303
rect 6144 33272 6193 33300
rect 6144 33260 6150 33272
rect 6181 33269 6193 33272
rect 6227 33269 6239 33303
rect 6181 33263 6239 33269
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 7576 33300 7604 33328
rect 11440 33312 11468 33408
rect 13446 33396 13452 33408
rect 13504 33436 13510 33448
rect 14001 33439 14059 33445
rect 14001 33436 14013 33439
rect 13504 33408 14013 33436
rect 13504 33396 13510 33408
rect 14001 33405 14013 33408
rect 14047 33405 14059 33439
rect 14001 33399 14059 33405
rect 6687 33272 7604 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 9674 33260 9680 33312
rect 9732 33300 9738 33312
rect 9953 33303 10011 33309
rect 9953 33300 9965 33303
rect 9732 33272 9965 33300
rect 9732 33260 9738 33272
rect 9953 33269 9965 33272
rect 9999 33269 10011 33303
rect 9953 33263 10011 33269
rect 10226 33260 10232 33312
rect 10284 33300 10290 33312
rect 10505 33303 10563 33309
rect 10505 33300 10517 33303
rect 10284 33272 10517 33300
rect 10284 33260 10290 33272
rect 10505 33269 10517 33272
rect 10551 33269 10563 33303
rect 10505 33263 10563 33269
rect 11422 33260 11428 33312
rect 11480 33300 11486 33312
rect 11609 33303 11667 33309
rect 11609 33300 11621 33303
rect 11480 33272 11621 33300
rect 11480 33260 11486 33272
rect 11609 33269 11621 33272
rect 11655 33269 11667 33303
rect 12710 33300 12716 33312
rect 12671 33272 12716 33300
rect 11609 33263 11667 33269
rect 12710 33260 12716 33272
rect 12768 33260 12774 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1670 33056 1676 33108
rect 1728 33096 1734 33108
rect 2041 33099 2099 33105
rect 2041 33096 2053 33099
rect 1728 33068 2053 33096
rect 1728 33056 1734 33068
rect 2041 33065 2053 33068
rect 2087 33065 2099 33099
rect 4614 33096 4620 33108
rect 4575 33068 4620 33096
rect 2041 33059 2099 33065
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 4706 33056 4712 33108
rect 4764 33096 4770 33108
rect 5077 33099 5135 33105
rect 5077 33096 5089 33099
rect 4764 33068 5089 33096
rect 4764 33056 4770 33068
rect 5077 33065 5089 33068
rect 5123 33065 5135 33099
rect 5077 33059 5135 33065
rect 5537 33099 5595 33105
rect 5537 33065 5549 33099
rect 5583 33096 5595 33099
rect 5718 33096 5724 33108
rect 5583 33068 5724 33096
rect 5583 33065 5595 33068
rect 5537 33059 5595 33065
rect 5718 33056 5724 33068
rect 5776 33096 5782 33108
rect 6730 33096 6736 33108
rect 5776 33068 6736 33096
rect 5776 33056 5782 33068
rect 6730 33056 6736 33068
rect 6788 33056 6794 33108
rect 7469 33099 7527 33105
rect 7469 33065 7481 33099
rect 7515 33096 7527 33099
rect 7650 33096 7656 33108
rect 7515 33068 7656 33096
rect 7515 33065 7527 33068
rect 7469 33059 7527 33065
rect 7650 33056 7656 33068
rect 7708 33096 7714 33108
rect 8665 33099 8723 33105
rect 7708 33068 8248 33096
rect 7708 33056 7714 33068
rect 1765 33031 1823 33037
rect 1765 32997 1777 33031
rect 1811 33028 1823 33031
rect 2682 33028 2688 33040
rect 1811 33000 2688 33028
rect 1811 32997 1823 33000
rect 1765 32991 1823 32997
rect 2682 32988 2688 33000
rect 2740 32988 2746 33040
rect 2774 32988 2780 33040
rect 2832 33028 2838 33040
rect 2869 33031 2927 33037
rect 2869 33028 2881 33031
rect 2832 33000 2881 33028
rect 2832 32988 2838 33000
rect 2869 32997 2881 33000
rect 2915 32997 2927 33031
rect 2869 32991 2927 32997
rect 6549 33031 6607 33037
rect 6549 32997 6561 33031
rect 6595 33028 6607 33031
rect 6638 33028 6644 33040
rect 6595 33000 6644 33028
rect 6595 32997 6607 33000
rect 6549 32991 6607 32997
rect 6638 32988 6644 33000
rect 6696 32988 6702 33040
rect 8110 33028 8116 33040
rect 8071 33000 8116 33028
rect 8110 32988 8116 33000
rect 8168 32988 8174 33040
rect 8220 33037 8248 33068
rect 8665 33065 8677 33099
rect 8711 33096 8723 33099
rect 8846 33096 8852 33108
rect 8711 33068 8852 33096
rect 8711 33065 8723 33068
rect 8665 33059 8723 33065
rect 8846 33056 8852 33068
rect 8904 33096 8910 33108
rect 9493 33099 9551 33105
rect 9493 33096 9505 33099
rect 8904 33068 9505 33096
rect 8904 33056 8910 33068
rect 9493 33065 9505 33068
rect 9539 33096 9551 33099
rect 10042 33096 10048 33108
rect 9539 33068 10048 33096
rect 9539 33065 9551 33068
rect 9493 33059 9551 33065
rect 10042 33056 10048 33068
rect 10100 33096 10106 33108
rect 10962 33096 10968 33108
rect 10100 33068 10968 33096
rect 10100 33056 10106 33068
rect 10962 33056 10968 33068
rect 11020 33056 11026 33108
rect 11517 33099 11575 33105
rect 11517 33065 11529 33099
rect 11563 33065 11575 33099
rect 11517 33059 11575 33065
rect 8205 33031 8263 33037
rect 8205 32997 8217 33031
rect 8251 33028 8263 33031
rect 8754 33028 8760 33040
rect 8251 33000 8760 33028
rect 8251 32997 8263 33000
rect 8205 32991 8263 32997
rect 8754 32988 8760 33000
rect 8812 33028 8818 33040
rect 9674 33028 9680 33040
rect 8812 33000 9680 33028
rect 8812 32988 8818 33000
rect 9674 32988 9680 33000
rect 9732 32988 9738 33040
rect 9950 33028 9956 33040
rect 9911 33000 9956 33028
rect 9950 32988 9956 33000
rect 10008 33028 10014 33040
rect 11532 33028 11560 33059
rect 10008 33000 11560 33028
rect 10008 32988 10014 33000
rect 2961 32963 3019 32969
rect 2961 32929 2973 32963
rect 3007 32960 3019 32963
rect 3142 32960 3148 32972
rect 3007 32932 3148 32960
rect 3007 32929 3019 32932
rect 2961 32923 3019 32929
rect 3142 32920 3148 32932
rect 3200 32960 3206 32972
rect 3881 32963 3939 32969
rect 3881 32960 3893 32963
rect 3200 32932 3893 32960
rect 3200 32920 3206 32932
rect 3881 32929 3893 32932
rect 3927 32960 3939 32963
rect 4338 32960 4344 32972
rect 3927 32932 4344 32960
rect 3927 32929 3939 32932
rect 3881 32923 3939 32929
rect 4338 32920 4344 32932
rect 4396 32960 4402 32972
rect 4709 32963 4767 32969
rect 4709 32960 4721 32963
rect 4396 32932 4721 32960
rect 4396 32920 4402 32932
rect 4709 32929 4721 32932
rect 4755 32929 4767 32963
rect 4709 32923 4767 32929
rect 6178 32920 6184 32972
rect 6236 32960 6242 32972
rect 6914 32960 6920 32972
rect 6236 32932 6920 32960
rect 6236 32920 6242 32932
rect 2869 32895 2927 32901
rect 2869 32861 2881 32895
rect 2915 32892 2927 32895
rect 3234 32892 3240 32904
rect 2915 32864 3240 32892
rect 2915 32861 2927 32864
rect 2869 32855 2927 32861
rect 3234 32852 3240 32864
rect 3292 32852 3298 32904
rect 4617 32895 4675 32901
rect 4617 32861 4629 32895
rect 4663 32892 4675 32895
rect 4890 32892 4896 32904
rect 4663 32864 4896 32892
rect 4663 32861 4675 32864
rect 4617 32855 4675 32861
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 6656 32901 6684 32932
rect 6914 32920 6920 32932
rect 6972 32920 6978 32972
rect 10137 32963 10195 32969
rect 10137 32929 10149 32963
rect 10183 32960 10195 32963
rect 10226 32960 10232 32972
rect 10183 32932 10232 32960
rect 10183 32929 10195 32932
rect 10137 32923 10195 32929
rect 10226 32920 10232 32932
rect 10284 32920 10290 32972
rect 10404 32963 10462 32969
rect 10404 32929 10416 32963
rect 10450 32960 10462 32963
rect 10778 32960 10784 32972
rect 10450 32932 10784 32960
rect 10450 32929 10462 32932
rect 10404 32923 10462 32929
rect 10778 32920 10784 32932
rect 10836 32920 10842 32972
rect 6549 32895 6607 32901
rect 6549 32861 6561 32895
rect 6595 32861 6607 32895
rect 6549 32855 6607 32861
rect 6641 32895 6699 32901
rect 6641 32861 6653 32895
rect 6687 32861 6699 32895
rect 8110 32892 8116 32904
rect 8071 32864 8116 32892
rect 6641 32855 6699 32861
rect 2406 32824 2412 32836
rect 2367 32796 2412 32824
rect 2406 32784 2412 32796
rect 2464 32784 2470 32836
rect 3421 32827 3479 32833
rect 3421 32793 3433 32827
rect 3467 32824 3479 32827
rect 3510 32824 3516 32836
rect 3467 32796 3516 32824
rect 3467 32793 3479 32796
rect 3421 32787 3479 32793
rect 3510 32784 3516 32796
rect 3568 32824 3574 32836
rect 4157 32827 4215 32833
rect 4157 32824 4169 32827
rect 3568 32796 4169 32824
rect 3568 32784 3574 32796
rect 4157 32793 4169 32796
rect 4203 32793 4215 32827
rect 4157 32787 4215 32793
rect 5905 32827 5963 32833
rect 5905 32793 5917 32827
rect 5951 32824 5963 32827
rect 6564 32824 6592 32855
rect 8110 32852 8116 32864
rect 8168 32852 8174 32904
rect 6730 32824 6736 32836
rect 5951 32796 6736 32824
rect 5951 32793 5963 32796
rect 5905 32787 5963 32793
rect 6730 32784 6736 32796
rect 6788 32784 6794 32836
rect 7282 32784 7288 32836
rect 7340 32824 7346 32836
rect 7653 32827 7711 32833
rect 7653 32824 7665 32827
rect 7340 32796 7665 32824
rect 7340 32784 7346 32796
rect 7653 32793 7665 32796
rect 7699 32793 7711 32827
rect 7653 32787 7711 32793
rect 6086 32756 6092 32768
rect 6047 32728 6092 32756
rect 6086 32716 6092 32728
rect 6144 32716 6150 32768
rect 7098 32756 7104 32768
rect 7059 32728 7104 32756
rect 7098 32716 7104 32728
rect 7156 32716 7162 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 2038 32512 2044 32564
rect 2096 32552 2102 32564
rect 3145 32555 3203 32561
rect 3145 32552 3157 32555
rect 2096 32524 3157 32552
rect 2096 32512 2102 32524
rect 3145 32521 3157 32524
rect 3191 32521 3203 32555
rect 3145 32515 3203 32521
rect 4338 32512 4344 32564
rect 4396 32552 4402 32564
rect 4525 32555 4583 32561
rect 4525 32552 4537 32555
rect 4396 32524 4537 32552
rect 4396 32512 4402 32524
rect 4525 32521 4537 32524
rect 4571 32552 4583 32555
rect 4614 32552 4620 32564
rect 4571 32524 4620 32552
rect 4571 32521 4583 32524
rect 4525 32515 4583 32521
rect 4614 32512 4620 32524
rect 4672 32512 4678 32564
rect 8294 32552 8300 32564
rect 8255 32524 8300 32552
rect 8294 32512 8300 32524
rect 8352 32512 8358 32564
rect 8386 32512 8392 32564
rect 8444 32552 8450 32564
rect 8662 32552 8668 32564
rect 8444 32524 8668 32552
rect 8444 32512 8450 32524
rect 8662 32512 8668 32524
rect 8720 32552 8726 32564
rect 9217 32555 9275 32561
rect 9217 32552 9229 32555
rect 8720 32524 9229 32552
rect 8720 32512 8726 32524
rect 9217 32521 9229 32524
rect 9263 32521 9275 32555
rect 9490 32552 9496 32564
rect 9451 32524 9496 32552
rect 9217 32515 9275 32521
rect 2409 32487 2467 32493
rect 2409 32453 2421 32487
rect 2455 32484 2467 32487
rect 3234 32484 3240 32496
rect 2455 32456 3240 32484
rect 2455 32453 2467 32456
rect 2409 32447 2467 32453
rect 3234 32444 3240 32456
rect 3292 32444 3298 32496
rect 4157 32487 4215 32493
rect 4157 32453 4169 32487
rect 4203 32484 4215 32487
rect 4890 32484 4896 32496
rect 4203 32456 4896 32484
rect 4203 32453 4215 32456
rect 4157 32447 4215 32453
rect 4890 32444 4896 32456
rect 4948 32444 4954 32496
rect 5258 32484 5264 32496
rect 5219 32456 5264 32484
rect 5258 32444 5264 32456
rect 5316 32444 5322 32496
rect 8754 32444 8760 32496
rect 8812 32484 8818 32496
rect 8849 32487 8907 32493
rect 8849 32484 8861 32487
rect 8812 32456 8861 32484
rect 8812 32444 8818 32456
rect 8849 32453 8861 32456
rect 8895 32453 8907 32487
rect 8849 32447 8907 32453
rect 1578 32416 1584 32428
rect 1539 32388 1584 32416
rect 1578 32376 1584 32388
rect 1636 32376 1642 32428
rect 3605 32419 3663 32425
rect 3605 32385 3617 32419
rect 3651 32416 3663 32419
rect 3970 32416 3976 32428
rect 3651 32388 3976 32416
rect 3651 32385 3663 32388
rect 3605 32379 3663 32385
rect 3970 32376 3976 32388
rect 4028 32376 4034 32428
rect 5718 32416 5724 32428
rect 5679 32388 5724 32416
rect 5718 32376 5724 32388
rect 5776 32376 5782 32428
rect 6273 32419 6331 32425
rect 6273 32385 6285 32419
rect 6319 32416 6331 32419
rect 6319 32388 7052 32416
rect 6319 32385 6331 32388
rect 6273 32379 6331 32385
rect 1394 32348 1400 32360
rect 1355 32320 1400 32348
rect 1394 32308 1400 32320
rect 1452 32308 1458 32360
rect 2774 32308 2780 32360
rect 2832 32348 2838 32360
rect 4154 32348 4160 32360
rect 2832 32320 4160 32348
rect 2832 32308 2838 32320
rect 4154 32308 4160 32320
rect 4212 32308 4218 32360
rect 5077 32351 5135 32357
rect 5077 32317 5089 32351
rect 5123 32348 5135 32351
rect 5442 32348 5448 32360
rect 5123 32320 5448 32348
rect 5123 32317 5135 32320
rect 5077 32311 5135 32317
rect 5442 32308 5448 32320
rect 5500 32348 5506 32360
rect 5813 32351 5871 32357
rect 5813 32348 5825 32351
rect 5500 32320 5825 32348
rect 5500 32308 5506 32320
rect 5813 32317 5825 32320
rect 5859 32317 5871 32351
rect 5813 32311 5871 32317
rect 5994 32308 6000 32360
rect 6052 32348 6058 32360
rect 6641 32351 6699 32357
rect 6641 32348 6653 32351
rect 6052 32320 6653 32348
rect 6052 32308 6058 32320
rect 6641 32317 6653 32320
rect 6687 32348 6699 32351
rect 6917 32351 6975 32357
rect 6917 32348 6929 32351
rect 6687 32320 6929 32348
rect 6687 32317 6699 32320
rect 6641 32311 6699 32317
rect 6917 32317 6929 32320
rect 6963 32317 6975 32351
rect 7024 32348 7052 32388
rect 7184 32351 7242 32357
rect 7184 32348 7196 32351
rect 7024 32320 7196 32348
rect 6917 32311 6975 32317
rect 7184 32317 7196 32320
rect 7230 32348 7242 32351
rect 7650 32348 7656 32360
rect 7230 32320 7656 32348
rect 7230 32317 7242 32320
rect 7184 32311 7242 32317
rect 3510 32240 3516 32292
rect 3568 32280 3574 32292
rect 3605 32283 3663 32289
rect 3605 32280 3617 32283
rect 3568 32252 3617 32280
rect 3568 32240 3574 32252
rect 3605 32249 3617 32252
rect 3651 32249 3663 32283
rect 3605 32243 3663 32249
rect 3697 32283 3755 32289
rect 3697 32249 3709 32283
rect 3743 32249 3755 32283
rect 6932 32280 6960 32311
rect 7650 32308 7656 32320
rect 7708 32308 7714 32360
rect 9232 32348 9260 32515
rect 9490 32512 9496 32524
rect 9548 32512 9554 32564
rect 10226 32512 10232 32564
rect 10284 32552 10290 32564
rect 10413 32555 10471 32561
rect 10413 32552 10425 32555
rect 10284 32524 10425 32552
rect 10284 32512 10290 32524
rect 10413 32521 10425 32524
rect 10459 32521 10471 32555
rect 10778 32552 10784 32564
rect 10739 32524 10784 32552
rect 10413 32515 10471 32521
rect 10778 32512 10784 32524
rect 10836 32512 10842 32564
rect 11149 32555 11207 32561
rect 11149 32521 11161 32555
rect 11195 32552 11207 32555
rect 12158 32552 12164 32564
rect 11195 32524 12164 32552
rect 11195 32521 11207 32524
rect 11149 32515 11207 32521
rect 12158 32512 12164 32524
rect 12216 32512 12222 32564
rect 10042 32416 10048 32428
rect 10003 32388 10048 32416
rect 10042 32376 10048 32388
rect 10100 32376 10106 32428
rect 10962 32348 10968 32360
rect 9232 32320 9996 32348
rect 10875 32320 10968 32348
rect 8478 32280 8484 32292
rect 6932 32252 8484 32280
rect 3697 32243 3755 32249
rect 2958 32172 2964 32224
rect 3016 32212 3022 32224
rect 3712 32212 3740 32243
rect 8478 32240 8484 32252
rect 8536 32240 8542 32292
rect 9398 32240 9404 32292
rect 9456 32280 9462 32292
rect 9968 32289 9996 32320
rect 10962 32308 10968 32320
rect 11020 32348 11026 32360
rect 11517 32351 11575 32357
rect 11517 32348 11529 32351
rect 11020 32320 11529 32348
rect 11020 32308 11026 32320
rect 11517 32317 11529 32320
rect 11563 32317 11575 32351
rect 11517 32311 11575 32317
rect 9769 32283 9827 32289
rect 9769 32280 9781 32283
rect 9456 32252 9781 32280
rect 9456 32240 9462 32252
rect 9769 32249 9781 32252
rect 9815 32249 9827 32283
rect 9769 32243 9827 32249
rect 9953 32283 10011 32289
rect 9953 32249 9965 32283
rect 9999 32249 10011 32283
rect 9953 32243 10011 32249
rect 3016 32184 3740 32212
rect 3016 32172 3022 32184
rect 5258 32172 5264 32224
rect 5316 32212 5322 32224
rect 5721 32215 5779 32221
rect 5721 32212 5733 32215
rect 5316 32184 5733 32212
rect 5316 32172 5322 32184
rect 5721 32181 5733 32184
rect 5767 32212 5779 32215
rect 6086 32212 6092 32224
rect 5767 32184 6092 32212
rect 5767 32181 5779 32184
rect 5721 32175 5779 32181
rect 6086 32172 6092 32184
rect 6144 32172 6150 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 1394 31968 1400 32020
rect 1452 32008 1458 32020
rect 1581 32011 1639 32017
rect 1581 32008 1593 32011
rect 1452 31980 1593 32008
rect 1452 31968 1458 31980
rect 1581 31977 1593 31980
rect 1627 31977 1639 32011
rect 2038 32008 2044 32020
rect 1999 31980 2044 32008
rect 1581 31971 1639 31977
rect 2038 31968 2044 31980
rect 2096 31968 2102 32020
rect 2409 32011 2467 32017
rect 2409 31977 2421 32011
rect 2455 32008 2467 32011
rect 2455 31980 2912 32008
rect 2455 31977 2467 31980
rect 2409 31971 2467 31977
rect 2884 31940 2912 31980
rect 2958 31968 2964 32020
rect 3016 32008 3022 32020
rect 3053 32011 3111 32017
rect 3053 32008 3065 32011
rect 3016 31980 3065 32008
rect 3016 31968 3022 31980
rect 3053 31977 3065 31980
rect 3099 31977 3111 32011
rect 3053 31971 3111 31977
rect 3513 32011 3571 32017
rect 3513 31977 3525 32011
rect 3559 32008 3571 32011
rect 3970 32008 3976 32020
rect 3559 31980 3976 32008
rect 3559 31977 3571 31980
rect 3513 31971 3571 31977
rect 3970 31968 3976 31980
rect 4028 31968 4034 32020
rect 5258 32008 5264 32020
rect 5219 31980 5264 32008
rect 5258 31968 5264 31980
rect 5316 31968 5322 32020
rect 6089 32011 6147 32017
rect 6089 31977 6101 32011
rect 6135 32008 6147 32011
rect 6178 32008 6184 32020
rect 6135 31980 6184 32008
rect 6135 31977 6147 31980
rect 6089 31971 6147 31977
rect 6178 31968 6184 31980
rect 6236 31968 6242 32020
rect 6457 32011 6515 32017
rect 6457 31977 6469 32011
rect 6503 32008 6515 32011
rect 6638 32008 6644 32020
rect 6503 31980 6644 32008
rect 6503 31977 6515 31980
rect 6457 31971 6515 31977
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 6730 31968 6736 32020
rect 6788 32008 6794 32020
rect 6899 32011 6957 32017
rect 6899 32008 6911 32011
rect 6788 31980 6911 32008
rect 6788 31968 6794 31980
rect 6899 31977 6911 31980
rect 6945 31977 6957 32011
rect 6899 31971 6957 31977
rect 7098 31968 7104 32020
rect 7156 32008 7162 32020
rect 8389 32011 8447 32017
rect 8389 32008 8401 32011
rect 7156 31980 8401 32008
rect 7156 31968 7162 31980
rect 8389 31977 8401 31980
rect 8435 31977 8447 32011
rect 9398 32008 9404 32020
rect 9359 31980 9404 32008
rect 8389 31971 8447 31977
rect 9398 31968 9404 31980
rect 9456 31968 9462 32020
rect 10781 32011 10839 32017
rect 10781 31977 10793 32011
rect 10827 32008 10839 32011
rect 11057 32011 11115 32017
rect 11057 32008 11069 32011
rect 10827 31980 11069 32008
rect 10827 31977 10839 31980
rect 10781 31971 10839 31977
rect 11057 31977 11069 31980
rect 11103 32008 11115 32011
rect 11103 31980 11928 32008
rect 11103 31977 11115 31980
rect 11057 31971 11115 31977
rect 11900 31952 11928 31980
rect 3142 31940 3148 31952
rect 2884 31912 3148 31940
rect 3142 31900 3148 31912
rect 3200 31940 3206 31952
rect 4249 31943 4307 31949
rect 4249 31940 4261 31943
rect 3200 31912 4261 31940
rect 3200 31900 3206 31912
rect 4249 31909 4261 31912
rect 4295 31909 4307 31943
rect 7190 31940 7196 31952
rect 7151 31912 7196 31940
rect 4249 31903 4307 31909
rect 7190 31900 7196 31912
rect 7248 31900 7254 31952
rect 7374 31940 7380 31952
rect 7335 31912 7380 31940
rect 7374 31900 7380 31912
rect 7432 31900 7438 31952
rect 7469 31943 7527 31949
rect 7469 31909 7481 31943
rect 7515 31940 7527 31943
rect 7650 31940 7656 31952
rect 7515 31912 7656 31940
rect 7515 31909 7527 31912
rect 7469 31903 7527 31909
rect 2866 31764 2872 31816
rect 2924 31804 2930 31816
rect 3142 31804 3148 31816
rect 2924 31776 3148 31804
rect 2924 31764 2930 31776
rect 3142 31764 3148 31776
rect 3200 31764 3206 31816
rect 6638 31764 6644 31816
rect 6696 31804 6702 31816
rect 7484 31804 7512 31903
rect 7650 31900 7656 31912
rect 7708 31900 7714 31952
rect 7929 31943 7987 31949
rect 7929 31909 7941 31943
rect 7975 31940 7987 31943
rect 8110 31940 8116 31952
rect 7975 31912 8116 31940
rect 7975 31909 7987 31912
rect 7929 31903 7987 31909
rect 8110 31900 8116 31912
rect 8168 31900 8174 31952
rect 9950 31900 9956 31952
rect 10008 31940 10014 31952
rect 10229 31943 10287 31949
rect 10229 31940 10241 31943
rect 10008 31912 10241 31940
rect 10008 31900 10014 31912
rect 10229 31909 10241 31912
rect 10275 31909 10287 31943
rect 10229 31903 10287 31909
rect 11146 31900 11152 31952
rect 11204 31940 11210 31952
rect 11790 31940 11796 31952
rect 11204 31912 11796 31940
rect 11204 31900 11210 31912
rect 11790 31900 11796 31912
rect 11848 31900 11854 31952
rect 11882 31900 11888 31952
rect 11940 31940 11946 31952
rect 11940 31912 11985 31940
rect 11940 31900 11946 31912
rect 8018 31832 8024 31884
rect 8076 31872 8082 31884
rect 8205 31875 8263 31881
rect 8205 31872 8217 31875
rect 8076 31844 8217 31872
rect 8076 31832 8082 31844
rect 8205 31841 8217 31844
rect 8251 31872 8263 31875
rect 8846 31872 8852 31884
rect 8251 31844 8852 31872
rect 8251 31841 8263 31844
rect 8205 31835 8263 31841
rect 8846 31832 8852 31844
rect 8904 31832 8910 31884
rect 10042 31832 10048 31884
rect 10100 31872 10106 31884
rect 10321 31875 10379 31881
rect 10321 31872 10333 31875
rect 10100 31844 10333 31872
rect 10100 31832 10106 31844
rect 10321 31841 10333 31844
rect 10367 31841 10379 31875
rect 10321 31835 10379 31841
rect 11315 31875 11373 31881
rect 11315 31841 11327 31875
rect 11361 31872 11373 31875
rect 12434 31872 12440 31884
rect 11361 31844 12440 31872
rect 11361 31841 11373 31844
rect 11315 31835 11373 31841
rect 12434 31832 12440 31844
rect 12492 31832 12498 31884
rect 9858 31804 9864 31816
rect 6696 31776 7512 31804
rect 9692 31776 9864 31804
rect 6696 31764 6702 31776
rect 9692 31748 9720 31776
rect 9858 31764 9864 31776
rect 9916 31764 9922 31816
rect 10226 31804 10232 31816
rect 10187 31776 10232 31804
rect 10226 31764 10232 31776
rect 10284 31764 10290 31816
rect 11793 31807 11851 31813
rect 11793 31773 11805 31807
rect 11839 31804 11851 31807
rect 11839 31776 11873 31804
rect 11839 31773 11851 31776
rect 11793 31767 11851 31773
rect 9674 31696 9680 31748
rect 9732 31696 9738 31748
rect 11808 31736 11836 31767
rect 12158 31736 12164 31748
rect 11808 31708 12164 31736
rect 12158 31696 12164 31708
rect 12216 31696 12222 31748
rect 8754 31628 8760 31680
rect 8812 31668 8818 31680
rect 9306 31668 9312 31680
rect 8812 31640 9312 31668
rect 8812 31628 8818 31640
rect 9306 31628 9312 31640
rect 9364 31628 9370 31680
rect 9766 31668 9772 31680
rect 9727 31640 9772 31668
rect 9766 31628 9772 31640
rect 9824 31628 9830 31680
rect 12529 31671 12587 31677
rect 12529 31637 12541 31671
rect 12575 31668 12587 31671
rect 12618 31668 12624 31680
rect 12575 31640 12624 31668
rect 12575 31637 12587 31640
rect 12529 31631 12587 31637
rect 12618 31628 12624 31640
rect 12676 31628 12682 31680
rect 12894 31668 12900 31680
rect 12855 31640 12900 31668
rect 12894 31628 12900 31640
rect 12952 31628 12958 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 6638 31464 6644 31476
rect 6599 31436 6644 31464
rect 6638 31424 6644 31436
rect 6696 31424 6702 31476
rect 7101 31467 7159 31473
rect 7101 31433 7113 31467
rect 7147 31464 7159 31467
rect 7190 31464 7196 31476
rect 7147 31436 7196 31464
rect 7147 31433 7159 31436
rect 7101 31427 7159 31433
rect 7190 31424 7196 31436
rect 7248 31424 7254 31476
rect 10042 31424 10048 31476
rect 10100 31464 10106 31476
rect 10229 31467 10287 31473
rect 10229 31464 10241 31467
rect 10100 31436 10241 31464
rect 10100 31424 10106 31436
rect 10229 31433 10241 31436
rect 10275 31433 10287 31467
rect 10229 31427 10287 31433
rect 10318 31424 10324 31476
rect 10376 31464 10382 31476
rect 10502 31464 10508 31476
rect 10376 31436 10508 31464
rect 10376 31424 10382 31436
rect 10502 31424 10508 31436
rect 10560 31424 10566 31476
rect 12618 31424 12624 31476
rect 12676 31424 12682 31476
rect 7374 31396 7380 31408
rect 7335 31368 7380 31396
rect 7374 31356 7380 31368
rect 7432 31396 7438 31408
rect 8018 31396 8024 31408
rect 7432 31368 8024 31396
rect 7432 31356 7438 31368
rect 8018 31356 8024 31368
rect 8076 31356 8082 31408
rect 9309 31399 9367 31405
rect 9309 31365 9321 31399
rect 9355 31396 9367 31399
rect 9950 31396 9956 31408
rect 9355 31368 9956 31396
rect 9355 31365 9367 31368
rect 9309 31359 9367 31365
rect 9950 31356 9956 31368
rect 10008 31356 10014 31408
rect 10873 31399 10931 31405
rect 10873 31365 10885 31399
rect 10919 31396 10931 31399
rect 12069 31399 12127 31405
rect 12069 31396 12081 31399
rect 10919 31368 12081 31396
rect 10919 31365 10931 31368
rect 10873 31359 10931 31365
rect 12069 31365 12081 31368
rect 12115 31365 12127 31399
rect 12526 31396 12532 31408
rect 12487 31368 12532 31396
rect 12069 31359 12127 31365
rect 12526 31356 12532 31368
rect 12584 31356 12590 31408
rect 8757 31331 8815 31337
rect 8757 31297 8769 31331
rect 8803 31328 8815 31331
rect 9769 31331 9827 31337
rect 9769 31328 9781 31331
rect 8803 31300 9781 31328
rect 8803 31297 8815 31300
rect 8757 31291 8815 31297
rect 9769 31297 9781 31300
rect 9815 31328 9827 31331
rect 10042 31328 10048 31340
rect 9815 31300 10048 31328
rect 9815 31297 9827 31300
rect 9769 31291 9827 31297
rect 10042 31288 10048 31300
rect 10100 31288 10106 31340
rect 11425 31331 11483 31337
rect 11425 31297 11437 31331
rect 11471 31328 11483 31331
rect 11882 31328 11888 31340
rect 11471 31300 11888 31328
rect 11471 31297 11483 31300
rect 11425 31291 11483 31297
rect 11882 31288 11888 31300
rect 11940 31328 11946 31340
rect 12342 31328 12348 31340
rect 11940 31300 12348 31328
rect 11940 31288 11946 31300
rect 12342 31288 12348 31300
rect 12400 31288 12406 31340
rect 12636 31328 12664 31424
rect 12897 31331 12955 31337
rect 12897 31328 12909 31331
rect 12636 31300 12909 31328
rect 12897 31297 12909 31300
rect 12943 31328 12955 31331
rect 13449 31331 13507 31337
rect 13449 31328 13461 31331
rect 12943 31300 13461 31328
rect 12943 31297 12955 31300
rect 12897 31291 12955 31297
rect 13449 31297 13461 31300
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 9125 31263 9183 31269
rect 9125 31229 9137 31263
rect 9171 31260 9183 31263
rect 9861 31263 9919 31269
rect 9861 31260 9873 31263
rect 9171 31232 9873 31260
rect 9171 31229 9183 31232
rect 9125 31223 9183 31229
rect 9861 31229 9873 31232
rect 9907 31260 9919 31263
rect 10778 31260 10784 31272
rect 9907 31232 10784 31260
rect 9907 31229 9919 31232
rect 9861 31223 9919 31229
rect 10778 31220 10784 31232
rect 10836 31220 10842 31272
rect 10870 31220 10876 31272
rect 10928 31260 10934 31272
rect 11054 31260 11060 31272
rect 10928 31232 11060 31260
rect 10928 31220 10934 31232
rect 11054 31220 11060 31232
rect 11112 31220 11118 31272
rect 11149 31263 11207 31269
rect 11149 31229 11161 31263
rect 11195 31260 11207 31263
rect 11238 31260 11244 31272
rect 11195 31232 11244 31260
rect 11195 31229 11207 31232
rect 11149 31223 11207 31229
rect 11164 31192 11192 31223
rect 11238 31220 11244 31232
rect 11296 31220 11302 31272
rect 11330 31220 11336 31272
rect 11388 31260 11394 31272
rect 11790 31260 11796 31272
rect 11388 31232 11796 31260
rect 11388 31220 11394 31232
rect 11790 31220 11796 31232
rect 11848 31220 11854 31272
rect 12434 31220 12440 31272
rect 12492 31260 12498 31272
rect 13081 31263 13139 31269
rect 13081 31260 13093 31263
rect 12492 31232 13093 31260
rect 12492 31220 12498 31232
rect 13081 31229 13093 31232
rect 13127 31229 13139 31263
rect 13081 31223 13139 31229
rect 10612 31164 11192 31192
rect 12069 31195 12127 31201
rect 9306 31084 9312 31136
rect 9364 31124 9370 31136
rect 9769 31127 9827 31133
rect 9769 31124 9781 31127
rect 9364 31096 9781 31124
rect 9364 31084 9370 31096
rect 9769 31093 9781 31096
rect 9815 31093 9827 31127
rect 9769 31087 9827 31093
rect 9858 31084 9864 31136
rect 9916 31124 9922 31136
rect 10612 31133 10640 31164
rect 12069 31161 12081 31195
rect 12115 31192 12127 31195
rect 12894 31192 12900 31204
rect 12115 31164 12900 31192
rect 12115 31161 12127 31164
rect 12069 31155 12127 31161
rect 12894 31152 12900 31164
rect 12952 31192 12958 31204
rect 12989 31195 13047 31201
rect 12989 31192 13001 31195
rect 12952 31164 13001 31192
rect 12952 31152 12958 31164
rect 12989 31161 13001 31164
rect 13035 31161 13047 31195
rect 12989 31155 13047 31161
rect 10597 31127 10655 31133
rect 10597 31124 10609 31127
rect 9916 31096 10609 31124
rect 9916 31084 9922 31096
rect 10597 31093 10609 31096
rect 10643 31093 10655 31127
rect 10597 31087 10655 31093
rect 11238 31084 11244 31136
rect 11296 31124 11302 31136
rect 11333 31127 11391 31133
rect 11333 31124 11345 31127
rect 11296 31096 11345 31124
rect 11296 31084 11302 31096
rect 11333 31093 11345 31096
rect 11379 31093 11391 31127
rect 12158 31124 12164 31136
rect 12119 31096 12164 31124
rect 11333 31087 11391 31093
rect 12158 31084 12164 31096
rect 12216 31084 12222 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 9950 30920 9956 30932
rect 9911 30892 9956 30920
rect 9950 30880 9956 30892
rect 10008 30880 10014 30932
rect 10226 30920 10232 30932
rect 10187 30892 10232 30920
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 12492 30892 12537 30920
rect 12492 30880 12498 30892
rect 1670 30852 1676 30864
rect 1631 30824 1676 30852
rect 1670 30812 1676 30824
rect 1728 30812 1734 30864
rect 10778 30852 10784 30864
rect 10739 30824 10784 30852
rect 10778 30812 10784 30824
rect 10836 30852 10842 30864
rect 11238 30852 11244 30864
rect 10836 30824 11244 30852
rect 10836 30812 10842 30824
rect 11238 30812 11244 30824
rect 11296 30812 11302 30864
rect 1397 30787 1455 30793
rect 1397 30753 1409 30787
rect 1443 30753 1455 30787
rect 1397 30747 1455 30753
rect 11324 30787 11382 30793
rect 11324 30753 11336 30787
rect 11370 30784 11382 30787
rect 12342 30784 12348 30796
rect 11370 30756 12348 30784
rect 11370 30753 11382 30756
rect 11324 30747 11382 30753
rect 1412 30716 1440 30747
rect 12342 30744 12348 30756
rect 12400 30744 12406 30796
rect 1670 30716 1676 30728
rect 1412 30688 1676 30716
rect 1670 30676 1676 30688
rect 1728 30676 1734 30728
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30685 11115 30719
rect 11057 30679 11115 30685
rect 6917 30583 6975 30589
rect 6917 30549 6929 30583
rect 6963 30580 6975 30583
rect 7374 30580 7380 30592
rect 6963 30552 7380 30580
rect 6963 30549 6975 30552
rect 6917 30543 6975 30549
rect 7374 30540 7380 30552
rect 7432 30540 7438 30592
rect 9306 30580 9312 30592
rect 9267 30552 9312 30580
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 11072 30580 11100 30679
rect 11238 30580 11244 30592
rect 11072 30552 11244 30580
rect 11238 30540 11244 30552
rect 11296 30540 11302 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 1670 30376 1676 30388
rect 1631 30348 1676 30376
rect 1670 30336 1676 30348
rect 1728 30336 1734 30388
rect 9306 30336 9312 30388
rect 9364 30376 9370 30388
rect 9861 30379 9919 30385
rect 9861 30376 9873 30379
rect 9364 30348 9873 30376
rect 9364 30336 9370 30348
rect 9861 30345 9873 30348
rect 9907 30345 9919 30379
rect 9861 30339 9919 30345
rect 6917 30311 6975 30317
rect 6917 30277 6929 30311
rect 6963 30308 6975 30311
rect 7006 30308 7012 30320
rect 6963 30280 7012 30308
rect 6963 30277 6975 30280
rect 6917 30271 6975 30277
rect 7006 30268 7012 30280
rect 7064 30268 7070 30320
rect 10134 30200 10140 30252
rect 10192 30240 10198 30252
rect 10410 30240 10416 30252
rect 10192 30212 10416 30240
rect 10192 30200 10198 30212
rect 10410 30200 10416 30212
rect 10468 30200 10474 30252
rect 11333 30243 11391 30249
rect 11333 30209 11345 30243
rect 11379 30240 11391 30243
rect 12158 30240 12164 30252
rect 11379 30212 12164 30240
rect 11379 30209 11391 30212
rect 11333 30203 11391 30209
rect 12158 30200 12164 30212
rect 12216 30200 12222 30252
rect 3329 30175 3387 30181
rect 3329 30141 3341 30175
rect 3375 30172 3387 30175
rect 3421 30175 3479 30181
rect 3421 30172 3433 30175
rect 3375 30144 3433 30172
rect 3375 30141 3387 30144
rect 3329 30135 3387 30141
rect 3421 30141 3433 30144
rect 3467 30172 3479 30175
rect 4246 30172 4252 30184
rect 3467 30144 4252 30172
rect 3467 30141 3479 30144
rect 3421 30135 3479 30141
rect 4246 30132 4252 30144
rect 4304 30132 4310 30184
rect 6641 30175 6699 30181
rect 6641 30141 6653 30175
rect 6687 30172 6699 30175
rect 7469 30175 7527 30181
rect 7469 30172 7481 30175
rect 6687 30144 7481 30172
rect 6687 30141 6699 30144
rect 6641 30135 6699 30141
rect 7469 30141 7481 30144
rect 7515 30172 7527 30175
rect 8202 30172 8208 30184
rect 7515 30144 8208 30172
rect 7515 30141 7527 30144
rect 7469 30135 7527 30141
rect 8202 30132 8208 30144
rect 8260 30132 8266 30184
rect 9677 30175 9735 30181
rect 9677 30141 9689 30175
rect 9723 30172 9735 30175
rect 11149 30175 11207 30181
rect 9723 30144 10456 30172
rect 9723 30141 9735 30144
rect 9677 30135 9735 30141
rect 3666 30107 3724 30113
rect 3666 30104 3678 30107
rect 3436 30076 3678 30104
rect 3436 30048 3464 30076
rect 3666 30073 3678 30076
rect 3712 30073 3724 30107
rect 3666 30067 3724 30073
rect 6273 30107 6331 30113
rect 6273 30073 6285 30107
rect 6319 30104 6331 30107
rect 7190 30104 7196 30116
rect 6319 30076 7196 30104
rect 6319 30073 6331 30076
rect 6273 30067 6331 30073
rect 7190 30064 7196 30076
rect 7248 30064 7254 30116
rect 7374 30104 7380 30116
rect 7335 30076 7380 30104
rect 7374 30064 7380 30076
rect 7432 30064 7438 30116
rect 9309 30107 9367 30113
rect 9309 30073 9321 30107
rect 9355 30104 9367 30107
rect 9766 30104 9772 30116
rect 9355 30076 9772 30104
rect 9355 30073 9367 30076
rect 9309 30067 9367 30073
rect 9766 30064 9772 30076
rect 9824 30064 9830 30116
rect 10134 30104 10140 30116
rect 10095 30076 10140 30104
rect 10134 30064 10140 30076
rect 10192 30064 10198 30116
rect 10428 30113 10456 30144
rect 11149 30141 11161 30175
rect 11195 30172 11207 30175
rect 11238 30172 11244 30184
rect 11195 30144 11244 30172
rect 11195 30141 11207 30144
rect 11149 30135 11207 30141
rect 11238 30132 11244 30144
rect 11296 30172 11302 30184
rect 11296 30144 12204 30172
rect 11296 30132 11302 30144
rect 12176 30116 12204 30144
rect 10413 30107 10471 30113
rect 10413 30073 10425 30107
rect 10459 30073 10471 30107
rect 10413 30067 10471 30073
rect 3418 29996 3424 30048
rect 3476 29996 3482 30048
rect 4430 29996 4436 30048
rect 4488 30036 4494 30048
rect 4801 30039 4859 30045
rect 4801 30036 4813 30039
rect 4488 30008 4813 30036
rect 4488 29996 4494 30008
rect 4801 30005 4813 30008
rect 4847 30005 4859 30039
rect 9784 30036 9812 30064
rect 10321 30039 10379 30045
rect 10321 30036 10333 30039
rect 9784 30008 10333 30036
rect 4801 29999 4859 30005
rect 10321 30005 10333 30008
rect 10367 30005 10379 30039
rect 10428 30036 10456 30067
rect 12158 30064 12164 30116
rect 12216 30064 12222 30116
rect 11885 30039 11943 30045
rect 11885 30036 11897 30039
rect 10428 30008 11897 30036
rect 10321 29999 10379 30005
rect 11885 30005 11897 30008
rect 11931 30036 11943 30039
rect 12342 30036 12348 30048
rect 11931 30008 12348 30036
rect 11931 30005 11943 30008
rect 11885 29999 11943 30005
rect 12342 29996 12348 30008
rect 12400 29996 12406 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 10311 29835 10369 29841
rect 10311 29801 10323 29835
rect 10357 29832 10369 29835
rect 12345 29835 12403 29841
rect 12345 29832 12357 29835
rect 10357 29804 12357 29832
rect 10357 29801 10369 29804
rect 10311 29795 10369 29801
rect 12345 29801 12357 29804
rect 12391 29832 12403 29835
rect 12618 29832 12624 29844
rect 12391 29804 12624 29832
rect 12391 29801 12403 29804
rect 12345 29795 12403 29801
rect 12618 29792 12624 29804
rect 12676 29792 12682 29844
rect 5436 29767 5494 29773
rect 5436 29733 5448 29767
rect 5482 29764 5494 29767
rect 5626 29764 5632 29776
rect 5482 29736 5632 29764
rect 5482 29733 5494 29736
rect 5436 29727 5494 29733
rect 5626 29724 5632 29736
rect 5684 29724 5690 29776
rect 6086 29724 6092 29776
rect 6144 29724 6150 29776
rect 6638 29724 6644 29776
rect 6696 29764 6702 29776
rect 8110 29764 8116 29776
rect 6696 29736 8116 29764
rect 6696 29724 6702 29736
rect 8110 29724 8116 29736
rect 8168 29764 8174 29776
rect 8205 29767 8263 29773
rect 8205 29764 8217 29767
rect 8168 29736 8217 29764
rect 8168 29724 8174 29736
rect 8205 29733 8217 29736
rect 8251 29733 8263 29767
rect 10594 29764 10600 29776
rect 10555 29736 10600 29764
rect 8205 29727 8263 29733
rect 10594 29724 10600 29736
rect 10652 29724 10658 29776
rect 10781 29767 10839 29773
rect 10781 29733 10793 29767
rect 10827 29764 10839 29767
rect 10870 29764 10876 29776
rect 10827 29736 10876 29764
rect 10827 29733 10839 29736
rect 10781 29727 10839 29733
rect 10870 29724 10876 29736
rect 10928 29724 10934 29776
rect 4246 29656 4252 29708
rect 4304 29696 4310 29708
rect 5169 29699 5227 29705
rect 5169 29696 5181 29699
rect 4304 29668 5181 29696
rect 4304 29656 4310 29668
rect 5169 29665 5181 29668
rect 5215 29696 5227 29699
rect 6104 29696 6132 29724
rect 6270 29696 6276 29708
rect 5215 29668 6276 29696
rect 5215 29665 5227 29668
rect 5169 29659 5227 29665
rect 6270 29656 6276 29668
rect 6328 29656 6334 29708
rect 7282 29656 7288 29708
rect 7340 29696 7346 29708
rect 8297 29699 8355 29705
rect 8297 29696 8309 29699
rect 7340 29668 8309 29696
rect 7340 29656 7346 29668
rect 8297 29665 8309 29668
rect 8343 29665 8355 29699
rect 8297 29659 8355 29665
rect 11974 29656 11980 29708
rect 12032 29696 12038 29708
rect 12161 29699 12219 29705
rect 12161 29696 12173 29699
rect 12032 29668 12173 29696
rect 12032 29656 12038 29668
rect 12161 29665 12173 29668
rect 12207 29696 12219 29699
rect 12250 29696 12256 29708
rect 12207 29668 12256 29696
rect 12207 29665 12219 29668
rect 12161 29659 12219 29665
rect 12250 29656 12256 29668
rect 12308 29656 12314 29708
rect 8113 29631 8171 29637
rect 8113 29597 8125 29631
rect 8159 29597 8171 29631
rect 10870 29628 10876 29640
rect 10831 29600 10876 29628
rect 8113 29591 8171 29597
rect 7190 29520 7196 29572
rect 7248 29560 7254 29572
rect 7745 29563 7803 29569
rect 7745 29560 7757 29563
rect 7248 29532 7757 29560
rect 7248 29520 7254 29532
rect 7745 29529 7757 29532
rect 7791 29529 7803 29563
rect 7745 29523 7803 29529
rect 3418 29492 3424 29504
rect 3379 29464 3424 29492
rect 3418 29452 3424 29464
rect 3476 29452 3482 29504
rect 5810 29452 5816 29504
rect 5868 29492 5874 29504
rect 6549 29495 6607 29501
rect 6549 29492 6561 29495
rect 5868 29464 6561 29492
rect 5868 29452 5874 29464
rect 6549 29461 6561 29464
rect 6595 29461 6607 29495
rect 6549 29455 6607 29461
rect 7101 29495 7159 29501
rect 7101 29461 7113 29495
rect 7147 29492 7159 29495
rect 7282 29492 7288 29504
rect 7147 29464 7288 29492
rect 7147 29461 7159 29464
rect 7101 29455 7159 29461
rect 7282 29452 7288 29464
rect 7340 29452 7346 29504
rect 7466 29492 7472 29504
rect 7427 29464 7472 29492
rect 7466 29452 7472 29464
rect 7524 29492 7530 29504
rect 8128 29492 8156 29591
rect 10870 29588 10876 29600
rect 10928 29588 10934 29640
rect 12342 29588 12348 29640
rect 12400 29628 12406 29640
rect 12437 29631 12495 29637
rect 12437 29628 12449 29631
rect 12400 29600 12449 29628
rect 12400 29588 12406 29600
rect 12437 29597 12449 29600
rect 12483 29597 12495 29631
rect 12437 29591 12495 29597
rect 10042 29520 10048 29572
rect 10100 29560 10106 29572
rect 11885 29563 11943 29569
rect 11885 29560 11897 29563
rect 10100 29532 11897 29560
rect 10100 29520 10106 29532
rect 11885 29529 11897 29532
rect 11931 29529 11943 29563
rect 11885 29523 11943 29529
rect 7524 29464 8156 29492
rect 7524 29452 7530 29464
rect 8478 29452 8484 29504
rect 8536 29492 8542 29504
rect 8665 29495 8723 29501
rect 8665 29492 8677 29495
rect 8536 29464 8677 29492
rect 8536 29452 8542 29464
rect 8665 29461 8677 29464
rect 8711 29461 8723 29495
rect 8665 29455 8723 29461
rect 9953 29495 10011 29501
rect 9953 29461 9965 29495
rect 9999 29492 10011 29495
rect 10134 29492 10140 29504
rect 9999 29464 10140 29492
rect 9999 29461 10011 29464
rect 9953 29455 10011 29461
rect 10134 29452 10140 29464
rect 10192 29492 10198 29504
rect 10686 29492 10692 29504
rect 10192 29464 10692 29492
rect 10192 29452 10198 29464
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 6917 29291 6975 29297
rect 6917 29257 6929 29291
rect 6963 29288 6975 29291
rect 7374 29288 7380 29300
rect 6963 29260 7380 29288
rect 6963 29257 6975 29260
rect 6917 29251 6975 29257
rect 7374 29248 7380 29260
rect 7432 29248 7438 29300
rect 9953 29291 10011 29297
rect 9953 29257 9965 29291
rect 9999 29288 10011 29291
rect 10226 29288 10232 29300
rect 9999 29260 10232 29288
rect 9999 29257 10011 29260
rect 9953 29251 10011 29257
rect 10226 29248 10232 29260
rect 10284 29288 10290 29300
rect 10870 29288 10876 29300
rect 10284 29260 10876 29288
rect 10284 29248 10290 29260
rect 10870 29248 10876 29260
rect 10928 29248 10934 29300
rect 12618 29288 12624 29300
rect 12579 29260 12624 29288
rect 12618 29248 12624 29260
rect 12676 29248 12682 29300
rect 10134 29180 10140 29232
rect 10192 29220 10198 29232
rect 10597 29223 10655 29229
rect 10597 29220 10609 29223
rect 10192 29192 10609 29220
rect 10192 29180 10198 29192
rect 10597 29189 10609 29192
rect 10643 29220 10655 29223
rect 10778 29220 10784 29232
rect 10643 29192 10784 29220
rect 10643 29189 10655 29192
rect 10597 29183 10655 29189
rect 10778 29180 10784 29192
rect 10836 29180 10842 29232
rect 4157 29155 4215 29161
rect 4157 29121 4169 29155
rect 4203 29152 4215 29155
rect 4246 29152 4252 29164
rect 4203 29124 4252 29152
rect 4203 29121 4215 29124
rect 4157 29115 4215 29121
rect 4246 29112 4252 29124
rect 4304 29112 4310 29164
rect 6641 29155 6699 29161
rect 6641 29121 6653 29155
rect 6687 29152 6699 29155
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 6687 29124 7389 29152
rect 6687 29121 6699 29124
rect 6641 29115 6699 29121
rect 7377 29121 7389 29124
rect 7423 29152 7435 29155
rect 7558 29152 7564 29164
rect 7423 29124 7564 29152
rect 7423 29121 7435 29124
rect 7377 29115 7435 29121
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 9950 29112 9956 29164
rect 10008 29152 10014 29164
rect 10873 29155 10931 29161
rect 10873 29152 10885 29155
rect 10008 29124 10885 29152
rect 10008 29112 10014 29124
rect 10873 29121 10885 29124
rect 10919 29121 10931 29155
rect 10873 29115 10931 29121
rect 8389 29087 8447 29093
rect 8389 29053 8401 29087
rect 8435 29084 8447 29087
rect 8573 29087 8631 29093
rect 8573 29084 8585 29087
rect 8435 29056 8585 29084
rect 8435 29053 8447 29056
rect 8389 29047 8447 29053
rect 8573 29053 8585 29056
rect 8619 29084 8631 29087
rect 8619 29056 9628 29084
rect 8619 29053 8631 29056
rect 8573 29047 8631 29053
rect 4430 28976 4436 29028
rect 4488 29025 4494 29028
rect 4488 29019 4552 29025
rect 4488 28985 4506 29019
rect 4540 28985 4552 29019
rect 4488 28979 4552 28985
rect 4488 28976 4494 28979
rect 4614 28976 4620 29028
rect 4672 29016 4678 29028
rect 4982 29016 4988 29028
rect 4672 28988 4988 29016
rect 4672 28976 4678 28988
rect 4982 28976 4988 28988
rect 5040 28976 5046 29028
rect 5534 28976 5540 29028
rect 5592 29016 5598 29028
rect 5994 29016 6000 29028
rect 5592 28988 6000 29016
rect 5592 28976 5598 28988
rect 5994 28976 6000 28988
rect 6052 28976 6058 29028
rect 6270 29016 6276 29028
rect 6183 28988 6276 29016
rect 6270 28976 6276 28988
rect 6328 29016 6334 29028
rect 6328 28988 6868 29016
rect 6328 28976 6334 28988
rect 5626 28948 5632 28960
rect 5587 28920 5632 28948
rect 5626 28908 5632 28920
rect 5684 28908 5690 28960
rect 6840 28948 6868 28988
rect 7282 28976 7288 29028
rect 7340 29016 7346 29028
rect 7469 29019 7527 29025
rect 7469 29016 7481 29019
rect 7340 28988 7481 29016
rect 7340 28976 7346 28988
rect 7469 28985 7481 28988
rect 7515 29016 7527 29019
rect 7742 29016 7748 29028
rect 7515 28988 7748 29016
rect 7515 28985 7527 28988
rect 7469 28979 7527 28985
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 7929 29019 7987 29025
rect 7929 28985 7941 29019
rect 7975 29016 7987 29019
rect 8110 29016 8116 29028
rect 7975 28988 8116 29016
rect 7975 28985 7987 28988
rect 7929 28979 7987 28985
rect 8110 28976 8116 28988
rect 8168 28976 8174 29028
rect 8404 29016 8432 29047
rect 8312 28988 8432 29016
rect 7098 28948 7104 28960
rect 6840 28920 7104 28948
rect 7098 28908 7104 28920
rect 7156 28908 7162 28960
rect 7374 28948 7380 28960
rect 7335 28920 7380 28948
rect 7374 28908 7380 28920
rect 7432 28908 7438 28960
rect 7834 28908 7840 28960
rect 7892 28948 7898 28960
rect 8312 28948 8340 28988
rect 8478 28976 8484 29028
rect 8536 29016 8542 29028
rect 8818 29019 8876 29025
rect 8818 29016 8830 29019
rect 8536 28988 8830 29016
rect 8536 28976 8542 28988
rect 8818 28985 8830 28988
rect 8864 28985 8876 29019
rect 8818 28979 8876 28985
rect 7892 28920 8340 28948
rect 9600 28948 9628 29056
rect 11885 29019 11943 29025
rect 11885 28985 11897 29019
rect 11931 29016 11943 29019
rect 11974 29016 11980 29028
rect 11931 28988 11980 29016
rect 11931 28985 11943 28988
rect 11885 28979 11943 28985
rect 11974 28976 11980 28988
rect 12032 28976 12038 29028
rect 11054 28948 11060 28960
rect 9600 28920 11060 28948
rect 7892 28908 7898 28920
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 12253 28951 12311 28957
rect 12253 28917 12265 28951
rect 12299 28948 12311 28951
rect 12342 28948 12348 28960
rect 12299 28920 12348 28948
rect 12299 28917 12311 28920
rect 12253 28911 12311 28917
rect 12342 28908 12348 28920
rect 12400 28908 12406 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 6917 28747 6975 28753
rect 6917 28713 6929 28747
rect 6963 28744 6975 28747
rect 7374 28744 7380 28756
rect 6963 28716 7380 28744
rect 6963 28713 6975 28716
rect 6917 28707 6975 28713
rect 7374 28704 7380 28716
rect 7432 28704 7438 28756
rect 8294 28704 8300 28756
rect 8352 28744 8358 28756
rect 8481 28747 8539 28753
rect 8481 28744 8493 28747
rect 8352 28716 8493 28744
rect 8352 28704 8358 28716
rect 8481 28713 8493 28716
rect 8527 28713 8539 28747
rect 10226 28744 10232 28756
rect 10187 28716 10232 28744
rect 8481 28707 8539 28713
rect 10226 28704 10232 28716
rect 10284 28704 10290 28756
rect 12342 28744 12348 28756
rect 12303 28716 12348 28744
rect 12342 28704 12348 28716
rect 12400 28704 12406 28756
rect 1670 28676 1676 28688
rect 1631 28648 1676 28676
rect 1670 28636 1676 28648
rect 1728 28636 1734 28688
rect 4062 28636 4068 28688
rect 4120 28676 4126 28688
rect 4522 28676 4528 28688
rect 4120 28648 4528 28676
rect 4120 28636 4126 28648
rect 4522 28636 4528 28648
rect 4580 28636 4586 28688
rect 4798 28636 4804 28688
rect 4856 28676 4862 28688
rect 5166 28676 5172 28688
rect 4856 28648 5172 28676
rect 4856 28636 4862 28648
rect 5166 28636 5172 28648
rect 5224 28676 5230 28688
rect 5353 28679 5411 28685
rect 5353 28676 5365 28679
rect 5224 28648 5365 28676
rect 5224 28636 5230 28648
rect 5353 28645 5365 28648
rect 5399 28645 5411 28679
rect 10244 28676 10272 28704
rect 11238 28685 11244 28688
rect 11210 28679 11244 28685
rect 11210 28676 11222 28679
rect 10244 28648 11222 28676
rect 5353 28639 5411 28645
rect 11210 28645 11222 28648
rect 11296 28676 11302 28688
rect 11296 28648 11358 28676
rect 11210 28639 11244 28645
rect 11238 28636 11244 28639
rect 11296 28636 11302 28648
rect 1397 28611 1455 28617
rect 1397 28577 1409 28611
rect 1443 28577 1455 28611
rect 1397 28571 1455 28577
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28608 4399 28611
rect 4430 28608 4436 28620
rect 4387 28580 4436 28608
rect 4387 28577 4399 28580
rect 4341 28571 4399 28577
rect 1412 28540 1440 28571
rect 4430 28568 4436 28580
rect 4488 28608 4494 28620
rect 6549 28611 6607 28617
rect 4488 28580 5488 28608
rect 4488 28568 4494 28580
rect 1670 28540 1676 28552
rect 1412 28512 1676 28540
rect 1670 28500 1676 28512
rect 1728 28500 1734 28552
rect 4522 28500 4528 28552
rect 4580 28540 4586 28552
rect 5074 28540 5080 28552
rect 4580 28512 5080 28540
rect 4580 28500 4586 28512
rect 5074 28500 5080 28512
rect 5132 28540 5138 28552
rect 5460 28549 5488 28580
rect 6549 28577 6561 28611
rect 6595 28608 6607 28611
rect 7368 28611 7426 28617
rect 7368 28608 7380 28611
rect 6595 28580 7380 28608
rect 6595 28577 6607 28580
rect 6549 28571 6607 28577
rect 7368 28577 7380 28580
rect 7414 28608 7426 28611
rect 7742 28608 7748 28620
rect 7414 28580 7748 28608
rect 7414 28577 7426 28580
rect 7368 28571 7426 28577
rect 7742 28568 7748 28580
rect 7800 28568 7806 28620
rect 10965 28611 11023 28617
rect 10965 28577 10977 28611
rect 11011 28608 11023 28611
rect 11054 28608 11060 28620
rect 11011 28580 11060 28608
rect 11011 28577 11023 28580
rect 10965 28571 11023 28577
rect 11054 28568 11060 28580
rect 11112 28568 11118 28620
rect 5261 28543 5319 28549
rect 5261 28540 5273 28543
rect 5132 28512 5273 28540
rect 5132 28500 5138 28512
rect 5261 28509 5273 28512
rect 5307 28509 5319 28543
rect 5261 28503 5319 28509
rect 5445 28543 5503 28549
rect 5445 28509 5457 28543
rect 5491 28540 5503 28543
rect 5902 28540 5908 28552
rect 5491 28512 5908 28540
rect 5491 28509 5503 28512
rect 5445 28503 5503 28509
rect 5902 28500 5908 28512
rect 5960 28500 5966 28552
rect 7098 28540 7104 28552
rect 7011 28512 7104 28540
rect 7098 28500 7104 28512
rect 7156 28500 7162 28552
rect 4709 28407 4767 28413
rect 4709 28373 4721 28407
rect 4755 28404 4767 28407
rect 4893 28407 4951 28413
rect 4893 28404 4905 28407
rect 4755 28376 4905 28404
rect 4755 28373 4767 28376
rect 4709 28367 4767 28373
rect 4893 28373 4905 28376
rect 4939 28404 4951 28407
rect 5442 28404 5448 28416
rect 4939 28376 5448 28404
rect 4939 28373 4951 28376
rect 4893 28367 4951 28373
rect 5442 28364 5448 28376
rect 5500 28364 5506 28416
rect 5626 28364 5632 28416
rect 5684 28404 5690 28416
rect 5813 28407 5871 28413
rect 5813 28404 5825 28407
rect 5684 28376 5825 28404
rect 5684 28364 5690 28376
rect 5813 28373 5825 28376
rect 5859 28373 5871 28407
rect 7116 28404 7144 28500
rect 7834 28404 7840 28416
rect 7116 28376 7840 28404
rect 5813 28367 5871 28373
rect 7834 28364 7840 28376
rect 7892 28364 7898 28416
rect 9858 28364 9864 28416
rect 9916 28404 9922 28416
rect 10597 28407 10655 28413
rect 10597 28404 10609 28407
rect 9916 28376 10609 28404
rect 9916 28364 9922 28376
rect 10597 28373 10609 28376
rect 10643 28373 10655 28407
rect 10597 28367 10655 28373
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 5902 28200 5908 28212
rect 5863 28172 5908 28200
rect 5902 28160 5908 28172
rect 5960 28160 5966 28212
rect 7653 28203 7711 28209
rect 7653 28169 7665 28203
rect 7699 28200 7711 28203
rect 7834 28200 7840 28212
rect 7699 28172 7840 28200
rect 7699 28169 7711 28172
rect 7653 28163 7711 28169
rect 7834 28160 7840 28172
rect 7892 28200 7898 28212
rect 7929 28203 7987 28209
rect 7929 28200 7941 28203
rect 7892 28172 7941 28200
rect 7892 28160 7898 28172
rect 7929 28169 7941 28172
rect 7975 28169 7987 28203
rect 7929 28163 7987 28169
rect 10137 28203 10195 28209
rect 10137 28169 10149 28203
rect 10183 28200 10195 28203
rect 10226 28200 10232 28212
rect 10183 28172 10232 28200
rect 10183 28169 10195 28172
rect 10137 28163 10195 28169
rect 4890 28092 4896 28144
rect 4948 28132 4954 28144
rect 4985 28135 5043 28141
rect 4985 28132 4997 28135
rect 4948 28104 4997 28132
rect 4948 28092 4954 28104
rect 4985 28101 4997 28104
rect 5031 28101 5043 28135
rect 4985 28095 5043 28101
rect 7101 28067 7159 28073
rect 7101 28033 7113 28067
rect 7147 28064 7159 28067
rect 7466 28064 7472 28076
rect 7147 28036 7472 28064
rect 7147 28033 7159 28036
rect 7101 28027 7159 28033
rect 7466 28024 7472 28036
rect 7524 28024 7530 28076
rect 7944 28064 7972 28163
rect 10226 28160 10232 28172
rect 10284 28160 10290 28212
rect 10410 28200 10416 28212
rect 10371 28172 10416 28200
rect 10410 28160 10416 28172
rect 10468 28160 10474 28212
rect 10686 28200 10692 28212
rect 10647 28172 10692 28200
rect 10686 28160 10692 28172
rect 10744 28160 10750 28212
rect 10778 28160 10784 28212
rect 10836 28200 10842 28212
rect 11054 28200 11060 28212
rect 10836 28172 11060 28200
rect 10836 28160 10842 28172
rect 11054 28160 11060 28172
rect 11112 28200 11118 28212
rect 11609 28203 11667 28209
rect 11609 28200 11621 28203
rect 11112 28172 11621 28200
rect 11112 28160 11118 28172
rect 11609 28169 11621 28172
rect 11655 28169 11667 28203
rect 11609 28163 11667 28169
rect 8113 28067 8171 28073
rect 8113 28064 8125 28067
rect 7944 28036 8125 28064
rect 8113 28033 8125 28036
rect 8159 28033 8171 28067
rect 11238 28064 11244 28076
rect 11199 28036 11244 28064
rect 8113 28027 8171 28033
rect 11238 28024 11244 28036
rect 11296 28024 11302 28076
rect 2409 27999 2467 28005
rect 2409 27965 2421 27999
rect 2455 27965 2467 27999
rect 2409 27959 2467 27965
rect 2424 27872 2452 27959
rect 2498 27888 2504 27940
rect 2556 27928 2562 27940
rect 2654 27931 2712 27937
rect 2654 27928 2666 27931
rect 2556 27900 2666 27928
rect 2556 27888 2562 27900
rect 2654 27897 2666 27900
rect 2700 27897 2712 27931
rect 2654 27891 2712 27897
rect 4433 27931 4491 27937
rect 4433 27897 4445 27931
rect 4479 27928 4491 27931
rect 5258 27928 5264 27940
rect 4479 27900 5264 27928
rect 4479 27897 4491 27900
rect 4433 27891 4491 27897
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 5442 27928 5448 27940
rect 5403 27900 5448 27928
rect 5442 27888 5448 27900
rect 5500 27888 5506 27940
rect 5537 27931 5595 27937
rect 5537 27897 5549 27931
rect 5583 27928 5595 27931
rect 5626 27928 5632 27940
rect 5583 27900 5632 27928
rect 5583 27897 5595 27900
rect 5537 27891 5595 27897
rect 5626 27888 5632 27900
rect 5684 27928 5690 27940
rect 6273 27931 6331 27937
rect 6273 27928 6285 27931
rect 5684 27900 6285 27928
rect 5684 27888 5690 27900
rect 6273 27897 6285 27900
rect 6319 27897 6331 27931
rect 6273 27891 6331 27897
rect 8294 27888 8300 27940
rect 8352 27937 8358 27940
rect 8352 27931 8416 27937
rect 8352 27897 8370 27931
rect 8404 27897 8416 27931
rect 8352 27891 8416 27897
rect 8352 27888 8358 27891
rect 9858 27888 9864 27940
rect 9916 27928 9922 27940
rect 10965 27931 11023 27937
rect 10965 27928 10977 27931
rect 9916 27900 10977 27928
rect 9916 27888 9922 27900
rect 10965 27897 10977 27900
rect 11011 27897 11023 27931
rect 10965 27891 11023 27897
rect 1670 27860 1676 27872
rect 1631 27832 1676 27860
rect 1670 27820 1676 27832
rect 1728 27820 1734 27872
rect 2317 27863 2375 27869
rect 2317 27829 2329 27863
rect 2363 27860 2375 27863
rect 2406 27860 2412 27872
rect 2363 27832 2412 27860
rect 2363 27829 2375 27832
rect 2317 27823 2375 27829
rect 2406 27820 2412 27832
rect 2464 27820 2470 27872
rect 2774 27820 2780 27872
rect 2832 27860 2838 27872
rect 3418 27860 3424 27872
rect 2832 27832 3424 27860
rect 2832 27820 2838 27832
rect 3418 27820 3424 27832
rect 3476 27860 3482 27872
rect 3789 27863 3847 27869
rect 3789 27860 3801 27863
rect 3476 27832 3801 27860
rect 3476 27820 3482 27832
rect 3789 27829 3801 27832
rect 3835 27829 3847 27863
rect 3789 27823 3847 27829
rect 4801 27863 4859 27869
rect 4801 27829 4813 27863
rect 4847 27860 4859 27863
rect 5166 27860 5172 27872
rect 4847 27832 5172 27860
rect 4847 27829 4859 27832
rect 4801 27823 4859 27829
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 8478 27820 8484 27872
rect 8536 27860 8542 27872
rect 9493 27863 9551 27869
rect 9493 27860 9505 27863
rect 8536 27832 9505 27860
rect 8536 27820 8542 27832
rect 9493 27829 9505 27832
rect 9539 27829 9551 27863
rect 9493 27823 9551 27829
rect 10410 27820 10416 27872
rect 10468 27860 10474 27872
rect 11149 27863 11207 27869
rect 11149 27860 11161 27863
rect 10468 27832 11161 27860
rect 10468 27820 10474 27832
rect 11149 27829 11161 27832
rect 11195 27829 11207 27863
rect 11149 27823 11207 27829
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 10410 27656 10416 27668
rect 10323 27628 10416 27656
rect 4154 27548 4160 27600
rect 4212 27588 4218 27600
rect 5537 27591 5595 27597
rect 5537 27588 5549 27591
rect 4212 27560 5549 27588
rect 4212 27548 4218 27560
rect 5537 27557 5549 27560
rect 5583 27588 5595 27591
rect 6730 27588 6736 27600
rect 5583 27560 6736 27588
rect 5583 27557 5595 27560
rect 5537 27551 5595 27557
rect 6730 27548 6736 27560
rect 6788 27548 6794 27600
rect 6914 27548 6920 27600
rect 6972 27588 6978 27600
rect 7101 27591 7159 27597
rect 7101 27588 7113 27591
rect 6972 27560 7113 27588
rect 6972 27548 6978 27560
rect 7101 27557 7113 27560
rect 7147 27557 7159 27591
rect 8202 27588 8208 27600
rect 8163 27560 8208 27588
rect 7101 27551 7159 27557
rect 8202 27548 8208 27560
rect 8260 27548 8266 27600
rect 10134 27588 10140 27600
rect 9968 27560 10140 27588
rect 5350 27520 5356 27532
rect 5311 27492 5356 27520
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 8294 27480 8300 27532
rect 8352 27520 8358 27532
rect 9968 27520 9996 27560
rect 10134 27548 10140 27560
rect 10192 27548 10198 27600
rect 10336 27597 10364 27628
rect 10410 27616 10416 27628
rect 10468 27656 10474 27668
rect 11057 27659 11115 27665
rect 11057 27656 11069 27659
rect 10468 27628 11069 27656
rect 10468 27616 10474 27628
rect 11057 27625 11069 27628
rect 11103 27656 11115 27659
rect 11238 27656 11244 27668
rect 11103 27628 11244 27656
rect 11103 27625 11115 27628
rect 11057 27619 11115 27625
rect 11238 27616 11244 27628
rect 11296 27616 11302 27668
rect 10229 27591 10287 27597
rect 10229 27557 10241 27591
rect 10275 27557 10287 27591
rect 10229 27551 10287 27557
rect 10321 27591 10379 27597
rect 10321 27557 10333 27591
rect 10367 27588 10379 27591
rect 10367 27560 10401 27588
rect 10367 27557 10379 27560
rect 10321 27551 10379 27557
rect 8352 27492 9996 27520
rect 8352 27480 8358 27492
rect 10244 27464 10272 27551
rect 5626 27452 5632 27464
rect 5587 27424 5632 27452
rect 5626 27412 5632 27424
rect 5684 27412 5690 27464
rect 6457 27455 6515 27461
rect 6457 27421 6469 27455
rect 6503 27452 6515 27455
rect 7006 27452 7012 27464
rect 6503 27424 7012 27452
rect 6503 27421 6515 27424
rect 6457 27415 6515 27421
rect 7006 27412 7012 27424
rect 7064 27412 7070 27464
rect 7190 27452 7196 27464
rect 7151 27424 7196 27452
rect 7190 27412 7196 27424
rect 7248 27452 7254 27464
rect 8478 27452 8484 27464
rect 7248 27424 8484 27452
rect 7248 27412 7254 27424
rect 8478 27412 8484 27424
rect 8536 27412 8542 27464
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27421 10195 27455
rect 10137 27415 10195 27421
rect 5534 27344 5540 27396
rect 5592 27384 5598 27396
rect 6641 27387 6699 27393
rect 6641 27384 6653 27387
rect 5592 27356 6653 27384
rect 5592 27344 5598 27356
rect 6641 27353 6653 27356
rect 6687 27353 6699 27387
rect 9766 27384 9772 27396
rect 9727 27356 9772 27384
rect 6641 27347 6699 27353
rect 9766 27344 9772 27356
rect 9824 27344 9830 27396
rect 10152 27384 10180 27415
rect 10226 27412 10232 27464
rect 10284 27412 10290 27464
rect 10060 27356 10180 27384
rect 10060 27328 10088 27356
rect 2498 27316 2504 27328
rect 2459 27288 2504 27316
rect 2498 27276 2504 27288
rect 2556 27276 2562 27328
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 4801 27319 4859 27325
rect 4801 27316 4813 27319
rect 4580 27288 4813 27316
rect 4580 27276 4586 27288
rect 4801 27285 4813 27288
rect 4847 27285 4859 27319
rect 5074 27316 5080 27328
rect 5035 27288 5080 27316
rect 4801 27279 4859 27285
rect 5074 27276 5080 27288
rect 5132 27276 5138 27328
rect 7653 27319 7711 27325
rect 7653 27285 7665 27319
rect 7699 27316 7711 27319
rect 7742 27316 7748 27328
rect 7699 27288 7748 27316
rect 7699 27285 7711 27288
rect 7653 27279 7711 27285
rect 7742 27276 7748 27288
rect 7800 27276 7806 27328
rect 10042 27276 10048 27328
rect 10100 27276 10106 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 4341 27115 4399 27121
rect 4341 27112 4353 27115
rect 4212 27084 4353 27112
rect 4212 27072 4218 27084
rect 4341 27081 4353 27084
rect 4387 27081 4399 27115
rect 4341 27075 4399 27081
rect 6641 27115 6699 27121
rect 6641 27081 6653 27115
rect 6687 27112 6699 27115
rect 7190 27112 7196 27124
rect 6687 27084 7196 27112
rect 6687 27081 6699 27084
rect 6641 27075 6699 27081
rect 7190 27072 7196 27084
rect 7248 27072 7254 27124
rect 9769 27115 9827 27121
rect 9769 27081 9781 27115
rect 9815 27112 9827 27115
rect 10226 27112 10232 27124
rect 9815 27084 10232 27112
rect 9815 27081 9827 27084
rect 9769 27075 9827 27081
rect 10226 27072 10232 27084
rect 10284 27072 10290 27124
rect 10410 27112 10416 27124
rect 10371 27084 10416 27112
rect 10410 27072 10416 27084
rect 10468 27072 10474 27124
rect 4614 27044 4620 27056
rect 4575 27016 4620 27044
rect 4614 27004 4620 27016
rect 4672 27004 4678 27056
rect 6914 27044 6920 27056
rect 6875 27016 6920 27044
rect 6914 27004 6920 27016
rect 6972 27004 6978 27056
rect 10042 27044 10048 27056
rect 10003 27016 10048 27044
rect 10042 27004 10048 27016
rect 10100 27004 10106 27056
rect 5074 26976 5080 26988
rect 5035 26948 5080 26976
rect 5074 26936 5080 26948
rect 5132 26976 5138 26988
rect 5905 26979 5963 26985
rect 5905 26976 5917 26979
rect 5132 26948 5917 26976
rect 5132 26936 5138 26948
rect 5905 26945 5917 26948
rect 5951 26945 5963 26979
rect 5905 26939 5963 26945
rect 6638 26936 6644 26988
rect 6696 26976 6702 26988
rect 7006 26976 7012 26988
rect 6696 26948 7012 26976
rect 6696 26936 6702 26948
rect 7006 26936 7012 26948
rect 7064 26936 7070 26988
rect 7098 26936 7104 26988
rect 7156 26976 7162 26988
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 7156 26948 7389 26976
rect 7156 26936 7162 26948
rect 7377 26945 7389 26948
rect 7423 26976 7435 26979
rect 8205 26979 8263 26985
rect 8205 26976 8217 26979
rect 7423 26948 8217 26976
rect 7423 26945 7435 26948
rect 7377 26939 7435 26945
rect 8205 26945 8217 26948
rect 8251 26945 8263 26979
rect 8205 26939 8263 26945
rect 4065 26911 4123 26917
rect 4065 26877 4077 26911
rect 4111 26908 4123 26911
rect 5169 26911 5227 26917
rect 5169 26908 5181 26911
rect 4111 26880 5181 26908
rect 4111 26877 4123 26880
rect 4065 26871 4123 26877
rect 5169 26877 5181 26880
rect 5215 26908 5227 26911
rect 5258 26908 5264 26920
rect 5215 26880 5264 26908
rect 5215 26877 5227 26880
rect 5169 26871 5227 26877
rect 5258 26868 5264 26880
rect 5316 26908 5322 26920
rect 5810 26908 5816 26920
rect 5316 26880 5816 26908
rect 5316 26868 5322 26880
rect 5810 26868 5816 26880
rect 5868 26868 5874 26920
rect 11330 26868 11336 26920
rect 11388 26908 11394 26920
rect 11514 26908 11520 26920
rect 11388 26880 11520 26908
rect 11388 26868 11394 26880
rect 11514 26868 11520 26880
rect 11572 26868 11578 26920
rect 13814 26868 13820 26920
rect 13872 26908 13878 26920
rect 15746 26908 15752 26920
rect 13872 26880 15752 26908
rect 13872 26868 13878 26880
rect 15746 26868 15752 26880
rect 15804 26868 15810 26920
rect 3697 26843 3755 26849
rect 3697 26809 3709 26843
rect 3743 26840 3755 26843
rect 4890 26840 4896 26852
rect 3743 26812 4896 26840
rect 3743 26809 3755 26812
rect 3697 26803 3755 26809
rect 4890 26800 4896 26812
rect 4948 26840 4954 26852
rect 5077 26843 5135 26849
rect 5077 26840 5089 26843
rect 4948 26812 5089 26840
rect 4948 26800 4954 26812
rect 5077 26809 5089 26812
rect 5123 26809 5135 26843
rect 5077 26803 5135 26809
rect 7006 26800 7012 26852
rect 7064 26840 7070 26852
rect 7469 26843 7527 26849
rect 7469 26840 7481 26843
rect 7064 26812 7481 26840
rect 7064 26800 7070 26812
rect 7469 26809 7481 26812
rect 7515 26840 7527 26843
rect 8202 26840 8208 26852
rect 7515 26812 8208 26840
rect 7515 26809 7527 26812
rect 7469 26803 7527 26809
rect 8202 26800 8208 26812
rect 8260 26800 8266 26852
rect 5350 26732 5356 26784
rect 5408 26772 5414 26784
rect 5534 26772 5540 26784
rect 5408 26744 5540 26772
rect 5408 26732 5414 26744
rect 5534 26732 5540 26744
rect 5592 26732 5598 26784
rect 7374 26772 7380 26784
rect 7287 26744 7380 26772
rect 7374 26732 7380 26744
rect 7432 26772 7438 26784
rect 7837 26775 7895 26781
rect 7837 26772 7849 26775
rect 7432 26744 7849 26772
rect 7432 26732 7438 26744
rect 7837 26741 7849 26744
rect 7883 26741 7895 26775
rect 7837 26735 7895 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 6549 26571 6607 26577
rect 6549 26537 6561 26571
rect 6595 26568 6607 26571
rect 6914 26568 6920 26580
rect 6595 26540 6920 26568
rect 6595 26537 6607 26540
rect 6549 26531 6607 26537
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 4614 26460 4620 26512
rect 4672 26500 4678 26512
rect 4801 26503 4859 26509
rect 4801 26500 4813 26503
rect 4672 26472 4813 26500
rect 4672 26460 4678 26472
rect 4801 26469 4813 26472
rect 4847 26500 4859 26503
rect 4982 26500 4988 26512
rect 4847 26472 4988 26500
rect 4847 26469 4859 26472
rect 4801 26463 4859 26469
rect 4982 26460 4988 26472
rect 5040 26460 5046 26512
rect 7558 26500 7564 26512
rect 7519 26472 7564 26500
rect 7558 26460 7564 26472
rect 7616 26460 7622 26512
rect 9306 26460 9312 26512
rect 9364 26500 9370 26512
rect 10229 26503 10287 26509
rect 10229 26500 10241 26503
rect 9364 26472 10241 26500
rect 9364 26460 9370 26472
rect 10229 26469 10241 26472
rect 10275 26469 10287 26503
rect 10229 26463 10287 26469
rect 6917 26435 6975 26441
rect 6917 26401 6929 26435
rect 6963 26432 6975 26435
rect 7006 26432 7012 26444
rect 6963 26404 7012 26432
rect 6963 26401 6975 26404
rect 6917 26395 6975 26401
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 9674 26392 9680 26444
rect 9732 26432 9738 26444
rect 10321 26435 10379 26441
rect 10321 26432 10333 26435
rect 9732 26404 10333 26432
rect 9732 26392 9738 26404
rect 10321 26401 10333 26404
rect 10367 26401 10379 26435
rect 10321 26395 10379 26401
rect 4798 26364 4804 26376
rect 4759 26336 4804 26364
rect 4798 26324 4804 26336
rect 4856 26324 4862 26376
rect 4890 26324 4896 26376
rect 4948 26364 4954 26376
rect 7466 26364 7472 26376
rect 4948 26336 4993 26364
rect 7427 26336 7472 26364
rect 4948 26324 4954 26336
rect 7466 26324 7472 26336
rect 7524 26324 7530 26376
rect 7653 26367 7711 26373
rect 7653 26333 7665 26367
rect 7699 26364 7711 26367
rect 7742 26364 7748 26376
rect 7699 26336 7748 26364
rect 7699 26333 7711 26336
rect 7653 26327 7711 26333
rect 7742 26324 7748 26336
rect 7800 26324 7806 26376
rect 10134 26364 10140 26376
rect 10095 26336 10140 26364
rect 10134 26324 10140 26336
rect 10192 26324 10198 26376
rect 4338 26296 4344 26308
rect 4299 26268 4344 26296
rect 4338 26256 4344 26268
rect 4396 26256 4402 26308
rect 5353 26299 5411 26305
rect 5353 26265 5365 26299
rect 5399 26296 5411 26299
rect 5626 26296 5632 26308
rect 5399 26268 5632 26296
rect 5399 26265 5411 26268
rect 5353 26259 5411 26265
rect 5626 26256 5632 26268
rect 5684 26296 5690 26308
rect 6086 26296 6092 26308
rect 5684 26268 6092 26296
rect 5684 26256 5690 26268
rect 6086 26256 6092 26268
rect 6144 26256 6150 26308
rect 7098 26296 7104 26308
rect 7059 26268 7104 26296
rect 7098 26256 7104 26268
rect 7156 26256 7162 26308
rect 9490 26256 9496 26308
rect 9548 26296 9554 26308
rect 9769 26299 9827 26305
rect 9769 26296 9781 26299
rect 9548 26268 9781 26296
rect 9548 26256 9554 26268
rect 9769 26265 9781 26268
rect 9815 26265 9827 26299
rect 9769 26259 9827 26265
rect 2777 26231 2835 26237
rect 2777 26197 2789 26231
rect 2823 26228 2835 26231
rect 3050 26228 3056 26240
rect 2823 26200 3056 26228
rect 2823 26197 2835 26200
rect 2777 26191 2835 26197
rect 3050 26188 3056 26200
rect 3108 26188 3114 26240
rect 7834 26188 7840 26240
rect 7892 26228 7898 26240
rect 8021 26231 8079 26237
rect 8021 26228 8033 26231
rect 7892 26200 8033 26228
rect 7892 26188 7898 26200
rect 8021 26197 8033 26200
rect 8067 26197 8079 26231
rect 8021 26191 8079 26197
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 2222 26024 2228 26036
rect 2183 25996 2228 26024
rect 2222 25984 2228 25996
rect 2280 25984 2286 26036
rect 2498 25984 2504 26036
rect 2556 26024 2562 26036
rect 3326 26024 3332 26036
rect 2556 25996 3332 26024
rect 2556 25984 2562 25996
rect 3326 25984 3332 25996
rect 3384 26024 3390 26036
rect 4065 26027 4123 26033
rect 4065 26024 4077 26027
rect 3384 25996 4077 26024
rect 3384 25984 3390 25996
rect 4065 25993 4077 25996
rect 4111 25993 4123 26027
rect 4982 26024 4988 26036
rect 4943 25996 4988 26024
rect 4065 25987 4123 25993
rect 4982 25984 4988 25996
rect 5040 25984 5046 26036
rect 7374 26024 7380 26036
rect 7335 25996 7380 26024
rect 7374 25984 7380 25996
rect 7432 25984 7438 26036
rect 4709 25959 4767 25965
rect 4709 25925 4721 25959
rect 4755 25956 4767 25959
rect 4890 25956 4896 25968
rect 4755 25928 4896 25956
rect 4755 25925 4767 25928
rect 4709 25919 4767 25925
rect 4890 25916 4896 25928
rect 4948 25916 4954 25968
rect 6730 25916 6736 25968
rect 6788 25956 6794 25968
rect 7101 25959 7159 25965
rect 7101 25956 7113 25959
rect 6788 25928 7113 25956
rect 6788 25916 6794 25928
rect 7101 25925 7113 25928
rect 7147 25956 7159 25959
rect 7466 25956 7472 25968
rect 7147 25928 7472 25956
rect 7147 25925 7159 25928
rect 7101 25919 7159 25925
rect 7466 25916 7472 25928
rect 7524 25916 7530 25968
rect 9122 25916 9128 25968
rect 9180 25956 9186 25968
rect 9677 25959 9735 25965
rect 9677 25956 9689 25959
rect 9180 25928 9689 25956
rect 9180 25916 9186 25928
rect 9677 25925 9689 25928
rect 9723 25925 9735 25959
rect 9950 25956 9956 25968
rect 9911 25928 9956 25956
rect 9677 25919 9735 25925
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 6273 25891 6331 25897
rect 6273 25857 6285 25891
rect 6319 25888 6331 25891
rect 7837 25891 7895 25897
rect 7837 25888 7849 25891
rect 6319 25860 7849 25888
rect 6319 25857 6331 25860
rect 6273 25851 6331 25857
rect 7837 25857 7849 25860
rect 7883 25888 7895 25891
rect 7926 25888 7932 25900
rect 7883 25860 7932 25888
rect 7883 25857 7895 25860
rect 7837 25851 7895 25857
rect 7926 25848 7932 25860
rect 7984 25848 7990 25900
rect 9692 25888 9720 25919
rect 9950 25916 9956 25928
rect 10008 25916 10014 25968
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 9692 25860 10333 25888
rect 10321 25857 10333 25860
rect 10367 25888 10379 25891
rect 10594 25888 10600 25900
rect 10367 25860 10600 25888
rect 10367 25857 10379 25860
rect 10321 25851 10379 25857
rect 10594 25848 10600 25860
rect 10652 25848 10658 25900
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25820 1455 25823
rect 2222 25820 2228 25832
rect 1443 25792 2228 25820
rect 1443 25789 1455 25792
rect 1397 25783 1455 25789
rect 2222 25780 2228 25792
rect 2280 25780 2286 25832
rect 2406 25780 2412 25832
rect 2464 25820 2470 25832
rect 2685 25823 2743 25829
rect 2685 25820 2697 25823
rect 2464 25792 2697 25820
rect 2464 25780 2470 25792
rect 2608 25696 2636 25792
rect 2685 25789 2697 25792
rect 2731 25789 2743 25823
rect 2685 25783 2743 25789
rect 9033 25823 9091 25829
rect 9033 25789 9045 25823
rect 9079 25820 9091 25823
rect 9306 25820 9312 25832
rect 9079 25792 9312 25820
rect 9079 25789 9091 25792
rect 9033 25783 9091 25789
rect 9306 25780 9312 25792
rect 9364 25820 9370 25832
rect 9674 25820 9680 25832
rect 9364 25792 9680 25820
rect 9364 25780 9370 25792
rect 9674 25780 9680 25792
rect 9732 25780 9738 25832
rect 2952 25755 3010 25761
rect 2952 25721 2964 25755
rect 2998 25752 3010 25755
rect 3050 25752 3056 25764
rect 2998 25724 3056 25752
rect 2998 25721 3010 25724
rect 2952 25715 3010 25721
rect 3050 25712 3056 25724
rect 3108 25712 3114 25764
rect 6641 25755 6699 25761
rect 6641 25721 6653 25755
rect 6687 25752 6699 25755
rect 7834 25752 7840 25764
rect 6687 25724 7604 25752
rect 7795 25724 7840 25752
rect 6687 25721 6699 25724
rect 6641 25715 6699 25721
rect 2590 25684 2596 25696
rect 2551 25656 2596 25684
rect 2590 25644 2596 25656
rect 2648 25644 2654 25696
rect 4798 25644 4804 25696
rect 4856 25684 4862 25696
rect 5353 25687 5411 25693
rect 5353 25684 5365 25687
rect 4856 25656 5365 25684
rect 4856 25644 4862 25656
rect 5353 25653 5365 25656
rect 5399 25653 5411 25687
rect 7576 25684 7604 25724
rect 7834 25712 7840 25724
rect 7892 25712 7898 25764
rect 7929 25755 7987 25761
rect 7929 25721 7941 25755
rect 7975 25721 7987 25755
rect 7929 25715 7987 25721
rect 10505 25755 10563 25761
rect 10505 25721 10517 25755
rect 10551 25752 10563 25755
rect 11054 25752 11060 25764
rect 10551 25724 11060 25752
rect 10551 25721 10563 25724
rect 10505 25715 10563 25721
rect 7742 25684 7748 25696
rect 7576 25656 7748 25684
rect 5353 25647 5411 25653
rect 7742 25644 7748 25656
rect 7800 25684 7806 25696
rect 7944 25684 7972 25715
rect 11054 25712 11060 25724
rect 11112 25712 11118 25764
rect 8389 25687 8447 25693
rect 8389 25684 8401 25687
rect 7800 25656 8401 25684
rect 7800 25644 7806 25656
rect 8389 25653 8401 25656
rect 8435 25684 8447 25687
rect 8478 25684 8484 25696
rect 8435 25656 8484 25684
rect 8435 25653 8447 25656
rect 8389 25647 8447 25653
rect 8478 25644 8484 25656
rect 8536 25644 8542 25696
rect 8570 25644 8576 25696
rect 8628 25684 8634 25696
rect 9214 25684 9220 25696
rect 8628 25656 9220 25684
rect 8628 25644 8634 25656
rect 9214 25644 9220 25656
rect 9272 25684 9278 25696
rect 9309 25687 9367 25693
rect 9309 25684 9321 25687
rect 9272 25656 9321 25684
rect 9272 25644 9278 25656
rect 9309 25653 9321 25656
rect 9355 25653 9367 25687
rect 9309 25647 9367 25653
rect 10413 25687 10471 25693
rect 10413 25653 10425 25687
rect 10459 25684 10471 25687
rect 10962 25684 10968 25696
rect 10459 25656 10968 25684
rect 10459 25653 10471 25656
rect 10413 25647 10471 25653
rect 10962 25644 10968 25656
rect 11020 25644 11026 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 2958 25480 2964 25492
rect 2919 25452 2964 25480
rect 2958 25440 2964 25452
rect 3016 25440 3022 25492
rect 5169 25483 5227 25489
rect 5169 25449 5181 25483
rect 5215 25480 5227 25483
rect 5258 25480 5264 25492
rect 5215 25452 5264 25480
rect 5215 25449 5227 25452
rect 5169 25443 5227 25449
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 8018 25480 8024 25492
rect 7979 25452 8024 25480
rect 8018 25440 8024 25452
rect 8076 25440 8082 25492
rect 9953 25483 10011 25489
rect 9953 25449 9965 25483
rect 9999 25480 10011 25483
rect 10134 25480 10140 25492
rect 9999 25452 10140 25480
rect 9999 25449 10011 25452
rect 9953 25443 10011 25449
rect 4154 25372 4160 25424
rect 4212 25412 4218 25424
rect 4617 25415 4675 25421
rect 4617 25412 4629 25415
rect 4212 25384 4629 25412
rect 4212 25372 4218 25384
rect 4617 25381 4629 25384
rect 4663 25381 4675 25415
rect 4617 25375 4675 25381
rect 4890 25372 4896 25424
rect 4948 25412 4954 25424
rect 5626 25412 5632 25424
rect 4948 25384 5632 25412
rect 4948 25372 4954 25384
rect 5626 25372 5632 25384
rect 5684 25412 5690 25424
rect 6058 25415 6116 25421
rect 6058 25412 6070 25415
rect 5684 25384 6070 25412
rect 5684 25372 5690 25384
rect 6058 25381 6070 25384
rect 6104 25381 6116 25415
rect 6058 25375 6116 25381
rect 9398 25372 9404 25424
rect 9456 25412 9462 25424
rect 9968 25412 9996 25443
rect 10134 25440 10140 25452
rect 10192 25440 10198 25492
rect 9456 25384 9996 25412
rect 9456 25372 9462 25384
rect 4706 25344 4712 25356
rect 3068 25316 4712 25344
rect 3068 25288 3096 25316
rect 4706 25304 4712 25316
rect 4764 25304 4770 25356
rect 5813 25347 5871 25353
rect 5813 25313 5825 25347
rect 5859 25344 5871 25347
rect 6638 25344 6644 25356
rect 5859 25316 6644 25344
rect 5859 25313 5871 25316
rect 5813 25307 5871 25313
rect 6638 25304 6644 25316
rect 6696 25304 6702 25356
rect 10778 25344 10784 25356
rect 10739 25316 10784 25344
rect 10778 25304 10784 25316
rect 10836 25304 10842 25356
rect 11054 25353 11060 25356
rect 11048 25344 11060 25353
rect 11015 25316 11060 25344
rect 11048 25307 11060 25316
rect 11054 25304 11060 25307
rect 11112 25304 11118 25356
rect 2958 25276 2964 25288
rect 2919 25248 2964 25276
rect 2958 25236 2964 25248
rect 3016 25236 3022 25288
rect 3050 25236 3056 25288
rect 3108 25276 3114 25288
rect 4614 25276 4620 25288
rect 3108 25248 3153 25276
rect 4575 25248 4620 25276
rect 3108 25236 3114 25248
rect 4614 25236 4620 25248
rect 4672 25236 4678 25288
rect 1949 25211 2007 25217
rect 1949 25177 1961 25211
rect 1995 25208 2007 25211
rect 2501 25211 2559 25217
rect 2501 25208 2513 25211
rect 1995 25180 2513 25208
rect 1995 25177 2007 25180
rect 1949 25171 2007 25177
rect 2501 25177 2513 25180
rect 2547 25208 2559 25211
rect 2774 25208 2780 25220
rect 2547 25180 2780 25208
rect 2547 25177 2559 25180
rect 2501 25171 2559 25177
rect 2774 25168 2780 25180
rect 2832 25168 2838 25220
rect 2317 25143 2375 25149
rect 2317 25109 2329 25143
rect 2363 25140 2375 25143
rect 3050 25140 3056 25152
rect 2363 25112 3056 25140
rect 2363 25109 2375 25112
rect 2317 25103 2375 25109
rect 3050 25100 3056 25112
rect 3108 25100 3114 25152
rect 3234 25100 3240 25152
rect 3292 25140 3298 25152
rect 3513 25143 3571 25149
rect 3513 25140 3525 25143
rect 3292 25112 3525 25140
rect 3292 25100 3298 25112
rect 3513 25109 3525 25112
rect 3559 25140 3571 25143
rect 4157 25143 4215 25149
rect 4157 25140 4169 25143
rect 3559 25112 4169 25140
rect 3559 25109 3571 25112
rect 3513 25103 3571 25109
rect 4157 25109 4169 25112
rect 4203 25109 4215 25143
rect 7190 25140 7196 25152
rect 7151 25112 7196 25140
rect 4157 25103 4215 25109
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 10321 25143 10379 25149
rect 10321 25109 10333 25143
rect 10367 25140 10379 25143
rect 11054 25140 11060 25152
rect 10367 25112 11060 25140
rect 10367 25109 10379 25112
rect 10321 25103 10379 25109
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 12158 25140 12164 25152
rect 12119 25112 12164 25140
rect 12158 25100 12164 25112
rect 12216 25100 12222 25152
rect 12805 25143 12863 25149
rect 12805 25109 12817 25143
rect 12851 25140 12863 25143
rect 13078 25140 13084 25152
rect 12851 25112 13084 25140
rect 12851 25109 12863 25112
rect 12805 25103 12863 25109
rect 13078 25100 13084 25112
rect 13136 25100 13142 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 2501 24939 2559 24945
rect 2501 24905 2513 24939
rect 2547 24936 2559 24939
rect 2866 24936 2872 24948
rect 2547 24908 2872 24936
rect 2547 24905 2559 24908
rect 2501 24899 2559 24905
rect 2866 24896 2872 24908
rect 2924 24896 2930 24948
rect 4157 24939 4215 24945
rect 4157 24905 4169 24939
rect 4203 24936 4215 24939
rect 4246 24936 4252 24948
rect 4203 24908 4252 24936
rect 4203 24905 4215 24908
rect 4157 24899 4215 24905
rect 4246 24896 4252 24908
rect 4304 24936 4310 24948
rect 4614 24936 4620 24948
rect 4304 24908 4620 24936
rect 4304 24896 4310 24908
rect 4614 24896 4620 24908
rect 4672 24896 4678 24948
rect 5626 24936 5632 24948
rect 5587 24908 5632 24936
rect 5626 24896 5632 24908
rect 5684 24936 5690 24948
rect 6549 24939 6607 24945
rect 6549 24936 6561 24939
rect 5684 24908 6561 24936
rect 5684 24896 5690 24908
rect 6549 24905 6561 24908
rect 6595 24905 6607 24939
rect 6549 24899 6607 24905
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 7377 24939 7435 24945
rect 7377 24936 7389 24939
rect 7248 24908 7389 24936
rect 7248 24896 7254 24908
rect 7377 24905 7389 24908
rect 7423 24905 7435 24939
rect 7377 24899 7435 24905
rect 7834 24896 7840 24948
rect 7892 24936 7898 24948
rect 8021 24939 8079 24945
rect 8021 24936 8033 24939
rect 7892 24908 8033 24936
rect 7892 24896 7898 24908
rect 8021 24905 8033 24908
rect 8067 24905 8079 24939
rect 10778 24936 10784 24948
rect 10739 24908 10784 24936
rect 8021 24899 8079 24905
rect 10778 24896 10784 24908
rect 10836 24936 10842 24948
rect 11146 24936 11152 24948
rect 10836 24908 11152 24936
rect 10836 24896 10842 24908
rect 11146 24896 11152 24908
rect 11204 24896 11210 24948
rect 12526 24936 12532 24948
rect 12487 24908 12532 24936
rect 12526 24896 12532 24908
rect 12584 24896 12590 24948
rect 2777 24871 2835 24877
rect 2777 24837 2789 24871
rect 2823 24837 2835 24871
rect 2777 24831 2835 24837
rect 6273 24871 6331 24877
rect 6273 24837 6285 24871
rect 6319 24868 6331 24871
rect 6638 24868 6644 24880
rect 6319 24840 6644 24868
rect 6319 24837 6331 24840
rect 6273 24831 6331 24837
rect 2314 24760 2320 24812
rect 2372 24800 2378 24812
rect 2792 24800 2820 24831
rect 3326 24800 3332 24812
rect 2372 24772 2820 24800
rect 3287 24772 3332 24800
rect 2372 24760 2378 24772
rect 3326 24760 3332 24772
rect 3384 24760 3390 24812
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1578 24732 1584 24744
rect 1443 24704 1584 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1578 24692 1584 24704
rect 1636 24692 1642 24744
rect 2774 24692 2780 24744
rect 2832 24732 2838 24744
rect 3053 24735 3111 24741
rect 3053 24732 3065 24735
rect 2832 24704 3065 24732
rect 2832 24692 2838 24704
rect 3053 24701 3065 24704
rect 3099 24701 3111 24735
rect 3053 24695 3111 24701
rect 3142 24692 3148 24744
rect 3200 24732 3206 24744
rect 3697 24735 3755 24741
rect 3697 24732 3709 24735
rect 3200 24704 3709 24732
rect 3200 24692 3206 24704
rect 3697 24701 3709 24704
rect 3743 24732 3755 24735
rect 4154 24732 4160 24744
rect 3743 24704 4160 24732
rect 3743 24701 3755 24704
rect 3697 24695 3755 24701
rect 4154 24692 4160 24704
rect 4212 24692 4218 24744
rect 4249 24735 4307 24741
rect 4249 24701 4261 24735
rect 4295 24701 4307 24735
rect 4249 24695 4307 24701
rect 4516 24735 4574 24741
rect 4516 24701 4528 24735
rect 4562 24732 4574 24735
rect 5258 24732 5264 24744
rect 4562 24704 5264 24732
rect 4562 24701 4574 24704
rect 4516 24695 4574 24701
rect 1670 24664 1676 24676
rect 1631 24636 1676 24664
rect 1670 24624 1676 24636
rect 1728 24624 1734 24676
rect 3234 24664 3240 24676
rect 3195 24636 3240 24664
rect 3234 24624 3240 24636
rect 3292 24624 3298 24676
rect 4264 24664 4292 24695
rect 5258 24692 5264 24704
rect 5316 24692 5322 24744
rect 4338 24664 4344 24676
rect 4251 24636 4344 24664
rect 4338 24624 4344 24636
rect 4396 24664 4402 24676
rect 4614 24664 4620 24676
rect 4396 24636 4620 24664
rect 4396 24624 4402 24636
rect 4614 24624 4620 24636
rect 4672 24664 4678 24676
rect 6288 24664 6316 24831
rect 6638 24828 6644 24840
rect 6696 24828 6702 24880
rect 9585 24871 9643 24877
rect 9585 24837 9597 24871
rect 9631 24837 9643 24871
rect 9585 24831 9643 24837
rect 7101 24803 7159 24809
rect 7101 24769 7113 24803
rect 7147 24800 7159 24803
rect 7558 24800 7564 24812
rect 7147 24772 7564 24800
rect 7147 24769 7159 24772
rect 7101 24763 7159 24769
rect 7558 24760 7564 24772
rect 7616 24800 7622 24812
rect 9600 24800 9628 24831
rect 7616 24772 9628 24800
rect 7616 24760 7622 24772
rect 12066 24760 12072 24812
rect 12124 24800 12130 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 12124 24772 12173 24800
rect 12124 24760 12130 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 8294 24732 8300 24744
rect 8255 24704 8300 24732
rect 8294 24692 8300 24704
rect 8352 24692 8358 24744
rect 8386 24692 8392 24744
rect 8444 24732 8450 24744
rect 8941 24735 8999 24741
rect 8941 24732 8953 24735
rect 8444 24704 8953 24732
rect 8444 24692 8450 24704
rect 8941 24701 8953 24704
rect 8987 24732 8999 24735
rect 9861 24735 9919 24741
rect 9861 24732 9873 24735
rect 8987 24704 9873 24732
rect 8987 24701 8999 24704
rect 8941 24695 8999 24701
rect 9861 24701 9873 24704
rect 9907 24701 9919 24735
rect 11790 24732 11796 24744
rect 11751 24704 11796 24732
rect 9861 24695 9919 24701
rect 11790 24692 11796 24704
rect 11848 24692 11854 24744
rect 8570 24664 8576 24676
rect 4672 24636 6316 24664
rect 8531 24636 8576 24664
rect 4672 24624 4678 24636
rect 8570 24624 8576 24636
rect 8628 24624 8634 24676
rect 10134 24664 10140 24676
rect 10095 24636 10140 24664
rect 10134 24624 10140 24636
rect 10192 24624 10198 24676
rect 7834 24596 7840 24608
rect 7747 24568 7840 24596
rect 7834 24556 7840 24568
rect 7892 24596 7898 24608
rect 8481 24599 8539 24605
rect 8481 24596 8493 24599
rect 7892 24568 8493 24596
rect 7892 24556 7898 24568
rect 8481 24565 8493 24568
rect 8527 24596 8539 24599
rect 8662 24596 8668 24608
rect 8527 24568 8668 24596
rect 8527 24565 8539 24568
rect 8481 24559 8539 24565
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 9401 24599 9459 24605
rect 9401 24565 9413 24599
rect 9447 24596 9459 24599
rect 9858 24596 9864 24608
rect 9447 24568 9864 24596
rect 9447 24565 9459 24568
rect 9401 24559 9459 24565
rect 9858 24556 9864 24568
rect 9916 24596 9922 24608
rect 10045 24599 10103 24605
rect 10045 24596 10057 24599
rect 9916 24568 10057 24596
rect 9916 24556 9922 24568
rect 10045 24565 10057 24568
rect 10091 24565 10103 24599
rect 10045 24559 10103 24565
rect 11054 24556 11060 24608
rect 11112 24596 11118 24608
rect 11149 24599 11207 24605
rect 11149 24596 11161 24599
rect 11112 24568 11161 24596
rect 11112 24556 11118 24568
rect 11149 24565 11161 24568
rect 11195 24565 11207 24599
rect 12176 24596 12204 24763
rect 12250 24692 12256 24744
rect 12308 24732 12314 24744
rect 13078 24732 13084 24744
rect 12308 24704 13084 24732
rect 12308 24692 12314 24704
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 12342 24624 12348 24676
rect 12400 24664 12406 24676
rect 12805 24667 12863 24673
rect 12805 24664 12817 24667
rect 12400 24636 12817 24664
rect 12400 24624 12406 24636
rect 12805 24633 12817 24636
rect 12851 24633 12863 24667
rect 12805 24627 12863 24633
rect 12989 24599 13047 24605
rect 12989 24596 13001 24599
rect 12176 24568 13001 24596
rect 11149 24559 11207 24565
rect 12989 24565 13001 24568
rect 13035 24565 13047 24599
rect 12989 24559 13047 24565
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24392 1642 24404
rect 2023 24395 2081 24401
rect 2023 24392 2035 24395
rect 1636 24364 2035 24392
rect 1636 24352 1642 24364
rect 2023 24361 2035 24364
rect 2069 24361 2081 24395
rect 2958 24392 2964 24404
rect 2919 24364 2964 24392
rect 2023 24355 2081 24361
rect 2958 24352 2964 24364
rect 3016 24392 3022 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 3016 24364 4077 24392
rect 3016 24352 3022 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4614 24392 4620 24404
rect 4575 24364 4620 24392
rect 4065 24355 4123 24361
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 4706 24352 4712 24404
rect 4764 24392 4770 24404
rect 4893 24395 4951 24401
rect 4893 24392 4905 24395
rect 4764 24364 4905 24392
rect 4764 24352 4770 24364
rect 4893 24361 4905 24364
rect 4939 24361 4951 24395
rect 4893 24355 4951 24361
rect 5718 24352 5724 24404
rect 5776 24392 5782 24404
rect 5905 24395 5963 24401
rect 5905 24392 5917 24395
rect 5776 24364 5917 24392
rect 5776 24352 5782 24364
rect 5905 24361 5917 24364
rect 5951 24361 5963 24395
rect 8478 24392 8484 24404
rect 8439 24364 8484 24392
rect 5905 24355 5963 24361
rect 8478 24352 8484 24364
rect 8536 24352 8542 24404
rect 11054 24352 11060 24404
rect 11112 24392 11118 24404
rect 12529 24395 12587 24401
rect 12529 24392 12541 24395
rect 11112 24364 12541 24392
rect 11112 24352 11118 24364
rect 12529 24361 12541 24364
rect 12575 24392 12587 24395
rect 13078 24392 13084 24404
rect 12575 24364 13084 24392
rect 12575 24361 12587 24364
rect 12529 24355 12587 24361
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 2498 24324 2504 24336
rect 2459 24296 2504 24324
rect 2498 24284 2504 24296
rect 2556 24284 2562 24336
rect 2593 24327 2651 24333
rect 2593 24293 2605 24327
rect 2639 24324 2651 24327
rect 2682 24324 2688 24336
rect 2639 24296 2688 24324
rect 2639 24293 2651 24296
rect 2593 24287 2651 24293
rect 2682 24284 2688 24296
rect 2740 24284 2746 24336
rect 3326 24324 3332 24336
rect 3287 24296 3332 24324
rect 3326 24284 3332 24296
rect 3384 24284 3390 24336
rect 7190 24284 7196 24336
rect 7248 24324 7254 24336
rect 7346 24327 7404 24333
rect 7346 24324 7358 24327
rect 7248 24296 7358 24324
rect 7248 24284 7254 24296
rect 7346 24293 7358 24296
rect 7392 24293 7404 24327
rect 11790 24324 11796 24336
rect 7346 24287 7404 24293
rect 11164 24296 11796 24324
rect 11164 24268 11192 24296
rect 11790 24284 11796 24296
rect 11848 24284 11854 24336
rect 2314 24256 2320 24268
rect 2275 24228 2320 24256
rect 2314 24216 2320 24228
rect 2372 24216 2378 24268
rect 6638 24216 6644 24268
rect 6696 24256 6702 24268
rect 7101 24259 7159 24265
rect 7101 24256 7113 24259
rect 6696 24228 7113 24256
rect 6696 24216 6702 24228
rect 7101 24225 7113 24228
rect 7147 24225 7159 24259
rect 7101 24219 7159 24225
rect 10226 24216 10232 24268
rect 10284 24256 10290 24268
rect 11146 24256 11152 24268
rect 10284 24228 11152 24256
rect 10284 24216 10290 24228
rect 11146 24216 11152 24228
rect 11204 24216 11210 24268
rect 11416 24259 11474 24265
rect 11416 24225 11428 24259
rect 11462 24256 11474 24259
rect 11974 24256 11980 24268
rect 11462 24228 11980 24256
rect 11462 24225 11474 24228
rect 11416 24219 11474 24225
rect 11974 24216 11980 24228
rect 12032 24256 12038 24268
rect 12250 24256 12256 24268
rect 12032 24228 12256 24256
rect 12032 24216 12038 24228
rect 12250 24216 12256 24228
rect 12308 24216 12314 24268
rect 5902 24188 5908 24200
rect 5863 24160 5908 24188
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24188 6055 24191
rect 6086 24188 6092 24200
rect 6043 24160 6092 24188
rect 6043 24157 6055 24160
rect 5997 24151 6055 24157
rect 6086 24148 6092 24160
rect 6144 24148 6150 24200
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 8628 24160 9873 24188
rect 8628 24148 8634 24160
rect 9861 24157 9873 24160
rect 9907 24188 9919 24191
rect 10134 24188 10140 24200
rect 9907 24160 10140 24188
rect 9907 24157 9919 24160
rect 9861 24151 9919 24157
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 5258 24012 5264 24064
rect 5316 24052 5322 24064
rect 5445 24055 5503 24061
rect 5445 24052 5457 24055
rect 5316 24024 5457 24052
rect 5316 24012 5322 24024
rect 5445 24021 5457 24024
rect 5491 24021 5503 24055
rect 5445 24015 5503 24021
rect 10873 24055 10931 24061
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11146 24052 11152 24064
rect 10919 24024 11152 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 2498 23848 2504 23860
rect 2363 23820 2504 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 2498 23808 2504 23820
rect 2556 23848 2562 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 2556 23820 3617 23848
rect 2556 23808 2562 23820
rect 3605 23817 3617 23820
rect 3651 23817 3663 23851
rect 4798 23848 4804 23860
rect 4759 23820 4804 23848
rect 3605 23811 3663 23817
rect 4798 23808 4804 23820
rect 4856 23808 4862 23860
rect 5813 23851 5871 23857
rect 5813 23817 5825 23851
rect 5859 23848 5871 23851
rect 5902 23848 5908 23860
rect 5859 23820 5908 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 6638 23808 6644 23860
rect 6696 23848 6702 23860
rect 7006 23848 7012 23860
rect 6696 23820 7012 23848
rect 6696 23808 6702 23820
rect 7006 23808 7012 23820
rect 7064 23848 7070 23860
rect 7285 23851 7343 23857
rect 7285 23848 7297 23851
rect 7064 23820 7297 23848
rect 7064 23808 7070 23820
rect 7285 23817 7297 23820
rect 7331 23817 7343 23851
rect 7926 23848 7932 23860
rect 7887 23820 7932 23848
rect 7285 23811 7343 23817
rect 7926 23808 7932 23820
rect 7984 23808 7990 23860
rect 11790 23848 11796 23860
rect 11751 23820 11796 23848
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 2041 23783 2099 23789
rect 2041 23749 2053 23783
rect 2087 23780 2099 23783
rect 2682 23780 2688 23792
rect 2087 23752 2688 23780
rect 2087 23749 2099 23752
rect 2041 23743 2099 23749
rect 2682 23740 2688 23752
rect 2740 23740 2746 23792
rect 4617 23783 4675 23789
rect 4617 23749 4629 23783
rect 4663 23780 4675 23783
rect 6086 23780 6092 23792
rect 4663 23752 6092 23780
rect 4663 23749 4675 23752
rect 4617 23743 4675 23749
rect 6086 23740 6092 23752
rect 6144 23740 6150 23792
rect 7558 23740 7564 23792
rect 7616 23780 7622 23792
rect 7653 23783 7711 23789
rect 7653 23780 7665 23783
rect 7616 23752 7665 23780
rect 7616 23740 7622 23752
rect 7653 23749 7665 23752
rect 7699 23749 7711 23783
rect 10594 23780 10600 23792
rect 10555 23752 10600 23780
rect 7653 23743 7711 23749
rect 10594 23740 10600 23752
rect 10652 23740 10658 23792
rect 10873 23783 10931 23789
rect 10873 23749 10885 23783
rect 10919 23780 10931 23783
rect 10962 23780 10968 23792
rect 10919 23752 10968 23780
rect 10919 23749 10931 23752
rect 10873 23743 10931 23749
rect 10962 23740 10968 23752
rect 11020 23740 11026 23792
rect 12250 23740 12256 23792
rect 12308 23780 12314 23792
rect 12529 23783 12587 23789
rect 12529 23780 12541 23783
rect 12308 23752 12541 23780
rect 12308 23740 12314 23752
rect 12529 23749 12541 23752
rect 12575 23749 12587 23783
rect 12529 23743 12587 23749
rect 2498 23672 2504 23724
rect 2556 23712 2562 23724
rect 2777 23715 2835 23721
rect 2777 23712 2789 23715
rect 2556 23684 2789 23712
rect 2556 23672 2562 23684
rect 2777 23681 2789 23684
rect 2823 23712 2835 23715
rect 3237 23715 3295 23721
rect 3237 23712 3249 23715
rect 2823 23684 3249 23712
rect 2823 23681 2835 23684
rect 2777 23675 2835 23681
rect 3237 23681 3249 23684
rect 3283 23681 3295 23715
rect 5350 23712 5356 23724
rect 5311 23684 5356 23712
rect 3237 23675 3295 23681
rect 5350 23672 5356 23684
rect 5408 23672 5414 23724
rect 7190 23672 7196 23724
rect 7248 23712 7254 23724
rect 8481 23715 8539 23721
rect 8481 23712 8493 23715
rect 7248 23684 8493 23712
rect 7248 23672 7254 23684
rect 8481 23681 8493 23684
rect 8527 23712 8539 23715
rect 8570 23712 8576 23724
rect 8527 23684 8576 23712
rect 8527 23681 8539 23684
rect 8481 23675 8539 23681
rect 8570 23672 8576 23684
rect 8628 23712 8634 23724
rect 8849 23715 8907 23721
rect 8849 23712 8861 23715
rect 8628 23684 8861 23712
rect 8628 23672 8634 23684
rect 8849 23681 8861 23684
rect 8895 23681 8907 23715
rect 13078 23712 13084 23724
rect 13039 23684 13084 23712
rect 8849 23675 8907 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 2682 23604 2688 23656
rect 2740 23644 2746 23656
rect 2869 23647 2927 23653
rect 2869 23644 2881 23647
rect 2740 23616 2881 23644
rect 2740 23604 2746 23616
rect 2869 23613 2881 23616
rect 2915 23644 2927 23647
rect 3326 23644 3332 23656
rect 2915 23616 3332 23644
rect 2915 23613 2927 23616
rect 2869 23607 2927 23613
rect 3326 23604 3332 23616
rect 3384 23604 3390 23656
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 4295 23616 5304 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 5276 23588 5304 23616
rect 5718 23604 5724 23656
rect 5776 23644 5782 23656
rect 6089 23647 6147 23653
rect 6089 23644 6101 23647
rect 5776 23616 6101 23644
rect 5776 23604 5782 23616
rect 6089 23613 6101 23616
rect 6135 23613 6147 23647
rect 6089 23607 6147 23613
rect 7926 23604 7932 23656
rect 7984 23644 7990 23656
rect 8205 23647 8263 23653
rect 8205 23644 8217 23647
rect 7984 23616 8217 23644
rect 7984 23604 7990 23616
rect 8205 23613 8217 23616
rect 8251 23644 8263 23647
rect 9398 23644 9404 23656
rect 8251 23616 9404 23644
rect 8251 23613 8263 23616
rect 8205 23607 8263 23613
rect 9398 23604 9404 23616
rect 9456 23604 9462 23656
rect 11146 23644 11152 23656
rect 11107 23616 11152 23644
rect 11146 23604 11152 23616
rect 11204 23604 11210 23656
rect 12253 23647 12311 23653
rect 12253 23613 12265 23647
rect 12299 23644 12311 23647
rect 12342 23644 12348 23656
rect 12299 23616 12348 23644
rect 12299 23613 12311 23616
rect 12253 23607 12311 23613
rect 12342 23604 12348 23616
rect 12400 23644 12406 23656
rect 12802 23644 12808 23656
rect 12400 23616 12808 23644
rect 12400 23604 12406 23616
rect 12802 23604 12808 23616
rect 12860 23604 12866 23656
rect 1673 23579 1731 23585
rect 1673 23545 1685 23579
rect 1719 23576 1731 23579
rect 2406 23576 2412 23588
rect 1719 23548 2412 23576
rect 1719 23545 1731 23548
rect 1673 23539 1731 23545
rect 2406 23536 2412 23548
rect 2464 23576 2470 23588
rect 2777 23579 2835 23585
rect 2777 23576 2789 23579
rect 2464 23548 2789 23576
rect 2464 23536 2470 23548
rect 2777 23545 2789 23548
rect 2823 23545 2835 23579
rect 2777 23539 2835 23545
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 4522 23576 4528 23588
rect 4120 23548 4528 23576
rect 4120 23536 4126 23548
rect 4522 23536 4528 23548
rect 4580 23536 4586 23588
rect 5074 23576 5080 23588
rect 5035 23548 5080 23576
rect 5074 23536 5080 23548
rect 5132 23536 5138 23588
rect 5258 23576 5264 23588
rect 5219 23548 5264 23576
rect 5258 23536 5264 23548
rect 5316 23536 5322 23588
rect 4982 23468 4988 23520
rect 5040 23508 5046 23520
rect 5736 23508 5764 23604
rect 5902 23536 5908 23588
rect 5960 23576 5966 23588
rect 6825 23579 6883 23585
rect 6825 23576 6837 23579
rect 5960 23548 6837 23576
rect 5960 23536 5966 23548
rect 6825 23545 6837 23548
rect 6871 23545 6883 23579
rect 11054 23576 11060 23588
rect 6825 23539 6883 23545
rect 10244 23548 11060 23576
rect 5040 23480 5764 23508
rect 5040 23468 5046 23480
rect 7558 23468 7564 23520
rect 7616 23508 7622 23520
rect 8110 23508 8116 23520
rect 7616 23480 8116 23508
rect 7616 23468 7622 23480
rect 8110 23468 8116 23480
rect 8168 23508 8174 23520
rect 8389 23511 8447 23517
rect 8389 23508 8401 23511
rect 8168 23480 8401 23508
rect 8168 23468 8174 23480
rect 8389 23477 8401 23480
rect 8435 23477 8447 23511
rect 8389 23471 8447 23477
rect 9398 23468 9404 23520
rect 9456 23508 9462 23520
rect 10244 23517 10272 23548
rect 11054 23536 11060 23548
rect 11112 23576 11118 23588
rect 11425 23579 11483 23585
rect 11425 23576 11437 23579
rect 11112 23548 11437 23576
rect 11112 23536 11118 23548
rect 11425 23545 11437 23548
rect 11471 23545 11483 23579
rect 11425 23539 11483 23545
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 9456 23480 10241 23508
rect 9456 23468 9462 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 10229 23471 10287 23477
rect 10594 23468 10600 23520
rect 10652 23508 10658 23520
rect 11333 23511 11391 23517
rect 11333 23508 11345 23511
rect 10652 23480 11345 23508
rect 10652 23468 10658 23480
rect 11333 23477 11345 23480
rect 11379 23477 11391 23511
rect 11333 23471 11391 23477
rect 12526 23468 12532 23520
rect 12584 23508 12590 23520
rect 12989 23511 13047 23517
rect 12989 23508 13001 23511
rect 12584 23480 13001 23508
rect 12584 23468 12590 23480
rect 12989 23477 13001 23480
rect 13035 23477 13047 23511
rect 12989 23471 13047 23477
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1949 23307 2007 23313
rect 1949 23273 1961 23307
rect 1995 23304 2007 23307
rect 2314 23304 2320 23316
rect 1995 23276 2320 23304
rect 1995 23273 2007 23276
rect 1949 23267 2007 23273
rect 2314 23264 2320 23276
rect 2372 23264 2378 23316
rect 5074 23304 5080 23316
rect 5035 23276 5080 23304
rect 5074 23264 5080 23276
rect 5132 23304 5138 23316
rect 5427 23307 5485 23313
rect 5427 23304 5439 23307
rect 5132 23276 5439 23304
rect 5132 23264 5138 23276
rect 5427 23273 5439 23276
rect 5473 23273 5485 23307
rect 5427 23267 5485 23273
rect 5905 23307 5963 23313
rect 5905 23273 5917 23307
rect 5951 23304 5963 23307
rect 5994 23304 6000 23316
rect 5951 23276 6000 23304
rect 5951 23273 5963 23276
rect 5905 23267 5963 23273
rect 5994 23264 6000 23276
rect 6052 23264 6058 23316
rect 7190 23304 7196 23316
rect 7151 23276 7196 23304
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 7926 23304 7932 23316
rect 7887 23276 7932 23304
rect 7926 23264 7932 23276
rect 7984 23264 7990 23316
rect 9950 23304 9956 23316
rect 9911 23276 9956 23304
rect 9950 23264 9956 23276
rect 10008 23264 10014 23316
rect 11146 23264 11152 23316
rect 11204 23304 11210 23316
rect 12069 23307 12127 23313
rect 12069 23304 12081 23307
rect 11204 23276 12081 23304
rect 11204 23264 11210 23276
rect 12069 23273 12081 23276
rect 12115 23273 12127 23307
rect 12069 23267 12127 23273
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12529 23307 12587 23313
rect 12529 23304 12541 23307
rect 12492 23276 12541 23304
rect 12492 23264 12498 23276
rect 12529 23273 12541 23276
rect 12575 23273 12587 23307
rect 12529 23267 12587 23273
rect 12989 23307 13047 23313
rect 12989 23273 13001 23307
rect 13035 23304 13047 23307
rect 13078 23304 13084 23316
rect 13035 23276 13084 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 2958 23236 2964 23248
rect 2919 23208 2964 23236
rect 2958 23196 2964 23208
rect 3016 23196 3022 23248
rect 6822 23236 6828 23248
rect 3988 23208 6828 23236
rect 2317 23171 2375 23177
rect 2317 23137 2329 23171
rect 2363 23168 2375 23171
rect 2682 23168 2688 23180
rect 2363 23140 2688 23168
rect 2363 23137 2375 23140
rect 2317 23131 2375 23137
rect 2682 23128 2688 23140
rect 2740 23128 2746 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 3234 23168 3240 23180
rect 2832 23140 3240 23168
rect 2832 23128 2838 23140
rect 3234 23128 3240 23140
rect 3292 23168 3298 23180
rect 3988 23168 4016 23208
rect 6822 23196 6828 23208
rect 6880 23196 6886 23248
rect 8570 23236 8576 23248
rect 8531 23208 8576 23236
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 11057 23239 11115 23245
rect 11057 23205 11069 23239
rect 11103 23236 11115 23239
rect 11606 23236 11612 23248
rect 11103 23208 11612 23236
rect 11103 23205 11115 23208
rect 11057 23199 11115 23205
rect 11606 23196 11612 23208
rect 11664 23236 11670 23248
rect 12250 23236 12256 23248
rect 11664 23208 12256 23236
rect 11664 23196 11670 23208
rect 12250 23196 12256 23208
rect 12308 23196 12314 23248
rect 3292 23140 4016 23168
rect 4801 23171 4859 23177
rect 3292 23128 3298 23140
rect 4801 23137 4813 23171
rect 4847 23168 4859 23171
rect 5350 23168 5356 23180
rect 4847 23140 5356 23168
rect 4847 23137 4859 23140
rect 4801 23131 4859 23137
rect 5350 23128 5356 23140
rect 5408 23128 5414 23180
rect 8389 23171 8447 23177
rect 8389 23137 8401 23171
rect 8435 23168 8447 23171
rect 8754 23168 8760 23180
rect 8435 23140 8760 23168
rect 8435 23137 8447 23140
rect 8389 23131 8447 23137
rect 8754 23128 8760 23140
rect 8812 23168 8818 23180
rect 9490 23168 9496 23180
rect 8812 23140 9496 23168
rect 8812 23128 8818 23140
rect 9490 23128 9496 23140
rect 9548 23128 9554 23180
rect 10686 23128 10692 23180
rect 10744 23168 10750 23180
rect 11149 23171 11207 23177
rect 11149 23168 11161 23171
rect 10744 23140 11161 23168
rect 10744 23128 10750 23140
rect 11149 23137 11161 23140
rect 11195 23168 11207 23171
rect 12158 23168 12164 23180
rect 11195 23140 12164 23168
rect 11195 23137 11207 23140
rect 11149 23131 11207 23137
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 3050 23100 3056 23112
rect 3011 23072 3056 23100
rect 3050 23060 3056 23072
rect 3108 23060 3114 23112
rect 5902 23100 5908 23112
rect 5863 23072 5908 23100
rect 5902 23060 5908 23072
rect 5960 23060 5966 23112
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23100 6055 23103
rect 6086 23100 6092 23112
rect 6043 23072 6092 23100
rect 6043 23069 6055 23072
rect 5997 23063 6055 23069
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 7190 23060 7196 23112
rect 7248 23100 7254 23112
rect 8665 23103 8723 23109
rect 8665 23100 8677 23103
rect 7248 23072 8677 23100
rect 7248 23060 7254 23072
rect 8665 23069 8677 23072
rect 8711 23100 8723 23103
rect 9398 23100 9404 23112
rect 8711 23072 9404 23100
rect 8711 23069 8723 23072
rect 8665 23063 8723 23069
rect 9398 23060 9404 23072
rect 9456 23060 9462 23112
rect 11054 23100 11060 23112
rect 11015 23072 11060 23100
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 2498 23032 2504 23044
rect 2459 23004 2504 23032
rect 2498 22992 2504 23004
rect 2556 22992 2562 23044
rect 8478 22992 8484 23044
rect 8536 23032 8542 23044
rect 9306 23032 9312 23044
rect 8536 23004 9312 23032
rect 8536 22992 8542 23004
rect 9306 22992 9312 23004
rect 9364 23032 9370 23044
rect 11517 23035 11575 23041
rect 11517 23032 11529 23035
rect 9364 23004 11529 23032
rect 9364 22992 9370 23004
rect 11517 23001 11529 23004
rect 11563 23032 11575 23035
rect 11974 23032 11980 23044
rect 11563 23004 11980 23032
rect 11563 23001 11575 23004
rect 11517 22995 11575 23001
rect 11974 22992 11980 23004
rect 12032 22992 12038 23044
rect 8110 22964 8116 22976
rect 8071 22936 8116 22964
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 10594 22964 10600 22976
rect 10555 22936 10600 22964
rect 10594 22924 10600 22936
rect 10652 22924 10658 22976
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2501 22763 2559 22769
rect 2501 22729 2513 22763
rect 2547 22760 2559 22763
rect 2774 22760 2780 22772
rect 2547 22732 2780 22760
rect 2547 22729 2559 22732
rect 2501 22723 2559 22729
rect 2774 22720 2780 22732
rect 2832 22720 2838 22772
rect 2869 22763 2927 22769
rect 2869 22729 2881 22763
rect 2915 22760 2927 22763
rect 2958 22760 2964 22772
rect 2915 22732 2964 22760
rect 2915 22729 2927 22732
rect 2869 22723 2927 22729
rect 2958 22720 2964 22732
rect 3016 22720 3022 22772
rect 5813 22763 5871 22769
rect 5813 22729 5825 22763
rect 5859 22760 5871 22763
rect 5902 22760 5908 22772
rect 5859 22732 5908 22760
rect 5859 22729 5871 22732
rect 5813 22723 5871 22729
rect 5902 22720 5908 22732
rect 5960 22720 5966 22772
rect 6086 22760 6092 22772
rect 6047 22732 6092 22760
rect 6086 22720 6092 22732
rect 6144 22720 6150 22772
rect 7190 22760 7196 22772
rect 7151 22732 7196 22760
rect 7190 22720 7196 22732
rect 7248 22720 7254 22772
rect 7834 22760 7840 22772
rect 7795 22732 7840 22760
rect 7834 22720 7840 22732
rect 7892 22720 7898 22772
rect 8113 22763 8171 22769
rect 8113 22729 8125 22763
rect 8159 22760 8171 22763
rect 8570 22760 8576 22772
rect 8159 22732 8576 22760
rect 8159 22729 8171 22732
rect 8113 22723 8171 22729
rect 8570 22720 8576 22732
rect 8628 22760 8634 22772
rect 9033 22763 9091 22769
rect 9033 22760 9045 22763
rect 8628 22732 9045 22760
rect 8628 22720 8634 22732
rect 9033 22729 9045 22732
rect 9079 22729 9091 22763
rect 9033 22723 9091 22729
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10318 22760 10324 22772
rect 9916 22732 10324 22760
rect 9916 22720 9922 22732
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 10686 22760 10692 22772
rect 10647 22732 10692 22760
rect 10686 22720 10692 22732
rect 10744 22720 10750 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 11333 22763 11391 22769
rect 11333 22760 11345 22763
rect 11112 22732 11345 22760
rect 11112 22720 11118 22732
rect 11333 22729 11345 22732
rect 11379 22729 11391 22763
rect 11333 22723 11391 22729
rect 5445 22695 5503 22701
rect 5445 22661 5457 22695
rect 5491 22692 5503 22695
rect 5626 22692 5632 22704
rect 5491 22664 5632 22692
rect 5491 22661 5503 22664
rect 5445 22655 5503 22661
rect 5626 22652 5632 22664
rect 5684 22692 5690 22704
rect 5994 22692 6000 22704
rect 5684 22664 6000 22692
rect 5684 22652 5690 22664
rect 5994 22652 6000 22664
rect 6052 22652 6058 22704
rect 9674 22692 9680 22704
rect 9635 22664 9680 22692
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22624 9551 22627
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 9539 22596 10241 22624
rect 9539 22593 9551 22596
rect 9493 22587 9551 22593
rect 10229 22593 10241 22596
rect 10275 22624 10287 22627
rect 10704 22624 10732 22720
rect 10275 22596 10732 22624
rect 11057 22627 11115 22633
rect 10275 22593 10287 22596
rect 10229 22587 10287 22593
rect 11057 22593 11069 22627
rect 11103 22624 11115 22627
rect 11606 22624 11612 22636
rect 11103 22596 11612 22624
rect 11103 22593 11115 22596
rect 11057 22587 11115 22593
rect 11606 22584 11612 22596
rect 11664 22584 11670 22636
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 7561 22559 7619 22565
rect 7561 22556 7573 22559
rect 6972 22528 7573 22556
rect 6972 22516 6978 22528
rect 7561 22525 7573 22528
rect 7607 22556 7619 22559
rect 8294 22556 8300 22568
rect 7607 22528 8300 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 8294 22516 8300 22528
rect 8352 22556 8358 22568
rect 8389 22559 8447 22565
rect 8389 22556 8401 22559
rect 8352 22528 8401 22556
rect 8352 22516 8358 22528
rect 8389 22525 8401 22528
rect 8435 22525 8447 22559
rect 9950 22556 9956 22568
rect 9911 22528 9956 22556
rect 8389 22519 8447 22525
rect 9950 22516 9956 22528
rect 10008 22516 10014 22568
rect 8478 22448 8484 22500
rect 8536 22488 8542 22500
rect 8665 22491 8723 22497
rect 8665 22488 8677 22491
rect 8536 22460 8677 22488
rect 8536 22448 8542 22460
rect 8665 22457 8677 22460
rect 8711 22457 8723 22491
rect 10134 22488 10140 22500
rect 10095 22460 10140 22488
rect 8665 22451 8723 22457
rect 10134 22448 10140 22460
rect 10192 22448 10198 22500
rect 10778 22448 10784 22500
rect 10836 22488 10842 22500
rect 11054 22488 11060 22500
rect 10836 22460 11060 22488
rect 10836 22448 10842 22460
rect 11054 22448 11060 22460
rect 11112 22448 11118 22500
rect 3050 22380 3056 22432
rect 3108 22420 3114 22432
rect 3145 22423 3203 22429
rect 3145 22420 3157 22423
rect 3108 22392 3157 22420
rect 3108 22380 3114 22392
rect 3145 22389 3157 22392
rect 3191 22389 3203 22423
rect 3145 22383 3203 22389
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 7892 22392 8585 22420
rect 7892 22380 7898 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 8573 22383 8631 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 4614 22216 4620 22228
rect 4120 22188 4620 22216
rect 4120 22176 4126 22188
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 8018 22176 8024 22228
rect 8076 22176 8082 22228
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8478 22216 8484 22228
rect 8343 22188 8484 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8478 22176 8484 22188
rect 8536 22176 8542 22228
rect 8665 22219 8723 22225
rect 8665 22185 8677 22219
rect 8711 22216 8723 22219
rect 8754 22216 8760 22228
rect 8711 22188 8760 22216
rect 8711 22185 8723 22188
rect 8665 22179 8723 22185
rect 8754 22176 8760 22188
rect 8812 22176 8818 22228
rect 9953 22219 10011 22225
rect 9953 22185 9965 22219
rect 9999 22216 10011 22219
rect 10134 22216 10140 22228
rect 9999 22188 10140 22216
rect 9999 22185 10011 22188
rect 9953 22179 10011 22185
rect 10134 22176 10140 22188
rect 10192 22176 10198 22228
rect 10321 22219 10379 22225
rect 10321 22185 10333 22219
rect 10367 22216 10379 22219
rect 10594 22216 10600 22228
rect 10367 22188 10600 22216
rect 10367 22185 10379 22188
rect 10321 22179 10379 22185
rect 10594 22176 10600 22188
rect 10652 22176 10658 22228
rect 2774 22108 2780 22160
rect 2832 22148 2838 22160
rect 2961 22151 3019 22157
rect 2961 22148 2973 22151
rect 2832 22120 2973 22148
rect 2832 22108 2838 22120
rect 2961 22117 2973 22120
rect 3007 22148 3019 22151
rect 6178 22148 6184 22160
rect 3007 22120 4108 22148
rect 6139 22120 6184 22148
rect 3007 22117 3019 22120
rect 2961 22111 3019 22117
rect 1486 22040 1492 22092
rect 1544 22080 1550 22092
rect 2130 22080 2136 22092
rect 1544 22052 2136 22080
rect 1544 22040 1550 22052
rect 2130 22040 2136 22052
rect 2188 22040 2194 22092
rect 3142 22080 3148 22092
rect 2976 22052 3148 22080
rect 2976 22021 3004 22052
rect 3142 22040 3148 22052
rect 3200 22040 3206 22092
rect 4080 22080 4108 22120
rect 6178 22108 6184 22120
rect 6236 22108 6242 22160
rect 7282 22108 7288 22160
rect 7340 22148 7346 22160
rect 7745 22151 7803 22157
rect 7745 22148 7757 22151
rect 7340 22120 7757 22148
rect 7340 22108 7346 22120
rect 7745 22117 7757 22120
rect 7791 22148 7803 22151
rect 8036 22148 8064 22176
rect 7791 22120 8064 22148
rect 7791 22117 7803 22120
rect 7745 22111 7803 22117
rect 10226 22108 10232 22160
rect 10284 22108 10290 22160
rect 10686 22108 10692 22160
rect 10744 22148 10750 22160
rect 11146 22157 11152 22160
rect 11118 22151 11152 22157
rect 11118 22148 11130 22151
rect 10744 22120 11130 22148
rect 10744 22108 10750 22120
rect 11118 22117 11130 22120
rect 11204 22148 11210 22160
rect 11204 22120 11266 22148
rect 11118 22111 11152 22117
rect 11146 22108 11152 22111
rect 11204 22108 11210 22120
rect 7558 22080 7564 22092
rect 4080 22052 4200 22080
rect 7519 22052 7564 22080
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 21981 3019 22015
rect 2961 21975 3019 21981
rect 3050 21972 3056 22024
rect 3108 22012 3114 22024
rect 3108 21984 3153 22012
rect 3108 21972 3114 21984
rect 2406 21904 2412 21956
rect 2464 21944 2470 21956
rect 4172 21953 4200 22052
rect 7558 22040 7564 22052
rect 7616 22040 7622 22092
rect 10244 22080 10272 22108
rect 10873 22083 10931 22089
rect 10873 22080 10885 22083
rect 10244 22052 10885 22080
rect 10873 22049 10885 22052
rect 10919 22080 10931 22083
rect 10962 22080 10968 22092
rect 10919 22052 10968 22080
rect 10919 22049 10931 22052
rect 10873 22043 10931 22049
rect 10962 22040 10968 22052
rect 11020 22040 11026 22092
rect 4525 22015 4583 22021
rect 4525 21981 4537 22015
rect 4571 21981 4583 22015
rect 4706 22012 4712 22024
rect 4667 21984 4712 22012
rect 4525 21975 4583 21981
rect 2501 21947 2559 21953
rect 2501 21944 2513 21947
rect 2464 21916 2513 21944
rect 2464 21904 2470 21916
rect 2501 21913 2513 21916
rect 2547 21913 2559 21947
rect 2501 21907 2559 21913
rect 4157 21947 4215 21953
rect 4157 21913 4169 21947
rect 4203 21913 4215 21947
rect 4540 21944 4568 21975
rect 4706 21972 4712 21984
rect 4764 21972 4770 22024
rect 6086 22012 6092 22024
rect 6047 21984 6092 22012
rect 6086 21972 6092 21984
rect 6144 21972 6150 22024
rect 6270 22012 6276 22024
rect 6231 21984 6276 22012
rect 6270 21972 6276 21984
rect 6328 21972 6334 22024
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 7374 22012 7380 22024
rect 7064 21984 7380 22012
rect 7064 21972 7070 21984
rect 7374 21972 7380 21984
rect 7432 21972 7438 22024
rect 7834 22012 7840 22024
rect 7795 21984 7840 22012
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 5534 21944 5540 21956
rect 4540 21916 5540 21944
rect 4157 21907 4215 21913
rect 5534 21904 5540 21916
rect 5592 21904 5598 21956
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4706 21876 4712 21888
rect 3927 21848 4712 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5718 21876 5724 21888
rect 5679 21848 5724 21876
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7285 21879 7343 21885
rect 7285 21876 7297 21879
rect 7064 21848 7297 21876
rect 7064 21836 7070 21848
rect 7285 21845 7297 21848
rect 7331 21845 7343 21879
rect 7285 21839 7343 21845
rect 10318 21836 10324 21888
rect 10376 21876 10382 21888
rect 12253 21879 12311 21885
rect 12253 21876 12265 21879
rect 10376 21848 12265 21876
rect 10376 21836 10382 21848
rect 12253 21845 12265 21848
rect 12299 21845 12311 21879
rect 12253 21839 12311 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 2133 21675 2191 21681
rect 2133 21641 2145 21675
rect 2179 21672 2191 21675
rect 3050 21672 3056 21684
rect 2179 21644 3056 21672
rect 2179 21641 2191 21644
rect 2133 21635 2191 21641
rect 3050 21632 3056 21644
rect 3108 21672 3114 21684
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 3108 21644 4905 21672
rect 3108 21632 3114 21644
rect 4893 21641 4905 21644
rect 4939 21641 4951 21675
rect 6178 21672 6184 21684
rect 6139 21644 6184 21672
rect 4893 21635 4951 21641
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 6638 21672 6644 21684
rect 6551 21644 6644 21672
rect 6638 21632 6644 21644
rect 6696 21672 6702 21684
rect 7834 21672 7840 21684
rect 6696 21644 7840 21672
rect 6696 21632 6702 21644
rect 7834 21632 7840 21644
rect 7892 21632 7898 21684
rect 10962 21672 10968 21684
rect 10923 21644 10968 21672
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11241 21675 11299 21681
rect 11241 21672 11253 21675
rect 11204 21644 11253 21672
rect 11204 21632 11210 21644
rect 11241 21641 11253 21644
rect 11287 21641 11299 21675
rect 11241 21635 11299 21641
rect 2406 21564 2412 21616
rect 2464 21604 2470 21616
rect 3142 21604 3148 21616
rect 2464 21576 3148 21604
rect 2464 21564 2470 21576
rect 3142 21564 3148 21576
rect 3200 21564 3206 21616
rect 5902 21604 5908 21616
rect 5815 21576 5908 21604
rect 5902 21564 5908 21576
rect 5960 21604 5966 21616
rect 6270 21604 6276 21616
rect 5960 21576 6276 21604
rect 5960 21564 5966 21576
rect 6270 21564 6276 21576
rect 6328 21564 6334 21616
rect 7742 21564 7748 21616
rect 7800 21604 7806 21616
rect 8205 21607 8263 21613
rect 8205 21604 8217 21607
rect 7800 21576 8217 21604
rect 7800 21564 7806 21576
rect 8205 21573 8217 21576
rect 8251 21573 8263 21607
rect 9766 21604 9772 21616
rect 9727 21576 9772 21604
rect 8205 21567 8263 21573
rect 9766 21564 9772 21576
rect 9824 21564 9830 21616
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 3099 21508 3648 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 3510 21468 3516 21480
rect 3471 21440 3516 21468
rect 3510 21428 3516 21440
rect 3568 21428 3574 21480
rect 3620 21468 3648 21508
rect 5166 21496 5172 21548
rect 5224 21536 5230 21548
rect 5534 21536 5540 21548
rect 5224 21508 5540 21536
rect 5224 21496 5230 21508
rect 5534 21496 5540 21508
rect 5592 21536 5598 21548
rect 6822 21536 6828 21548
rect 5592 21508 6828 21536
rect 5592 21496 5598 21508
rect 6822 21496 6828 21508
rect 6880 21496 6886 21548
rect 7650 21496 7656 21548
rect 7708 21536 7714 21548
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7708 21508 7941 21536
rect 7708 21496 7714 21508
rect 7929 21505 7941 21508
rect 7975 21536 7987 21539
rect 8018 21536 8024 21548
rect 7975 21508 8024 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 8018 21496 8024 21508
rect 8076 21536 8082 21548
rect 10229 21539 10287 21545
rect 8076 21508 8616 21536
rect 8076 21496 8082 21508
rect 3780 21471 3838 21477
rect 3780 21468 3792 21471
rect 3620 21440 3792 21468
rect 3780 21437 3792 21440
rect 3826 21468 3838 21471
rect 4706 21468 4712 21480
rect 3826 21440 4712 21468
rect 3826 21437 3838 21440
rect 3780 21431 3838 21437
rect 4706 21428 4712 21440
rect 4764 21428 4770 21480
rect 7098 21428 7104 21480
rect 7156 21468 7162 21480
rect 7156 21440 8340 21468
rect 7156 21428 7162 21440
rect 8312 21412 8340 21440
rect 8294 21360 8300 21412
rect 8352 21400 8358 21412
rect 8481 21403 8539 21409
rect 8481 21400 8493 21403
rect 8352 21372 8493 21400
rect 8352 21360 8358 21372
rect 8481 21369 8493 21372
rect 8527 21369 8539 21403
rect 8481 21363 8539 21369
rect 2406 21332 2412 21344
rect 2367 21304 2412 21332
rect 2406 21292 2412 21304
rect 2464 21292 2470 21344
rect 3142 21292 3148 21344
rect 3200 21332 3206 21344
rect 3329 21335 3387 21341
rect 3329 21332 3341 21335
rect 3200 21304 3341 21332
rect 3200 21292 3206 21304
rect 3329 21301 3341 21304
rect 3375 21332 3387 21335
rect 4062 21332 4068 21344
rect 3375 21304 4068 21332
rect 3375 21301 3387 21304
rect 3329 21295 3387 21301
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 7282 21332 7288 21344
rect 7243 21304 7288 21332
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7558 21332 7564 21344
rect 7519 21304 7564 21332
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 8588 21332 8616 21508
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 10594 21536 10600 21548
rect 10275 21508 10600 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 9585 21471 9643 21477
rect 9585 21437 9597 21471
rect 9631 21468 9643 21471
rect 10318 21468 10324 21480
rect 9631 21440 10324 21468
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 8754 21400 8760 21412
rect 8715 21372 8760 21400
rect 8754 21360 8760 21372
rect 8812 21360 8818 21412
rect 9217 21403 9275 21409
rect 9217 21369 9229 21403
rect 9263 21400 9275 21403
rect 9674 21400 9680 21412
rect 9263 21372 9680 21400
rect 9263 21369 9275 21372
rect 9217 21363 9275 21369
rect 9674 21360 9680 21372
rect 9732 21400 9738 21412
rect 10229 21403 10287 21409
rect 10229 21400 10241 21403
rect 9732 21372 10241 21400
rect 9732 21360 9738 21372
rect 10229 21369 10241 21372
rect 10275 21369 10287 21403
rect 10229 21363 10287 21369
rect 8665 21335 8723 21341
rect 8665 21332 8677 21335
rect 8588 21304 8677 21332
rect 8665 21301 8677 21304
rect 8711 21301 8723 21335
rect 8665 21295 8723 21301
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 2501 21131 2559 21137
rect 2501 21097 2513 21131
rect 2547 21128 2559 21131
rect 2682 21128 2688 21140
rect 2547 21100 2688 21128
rect 2547 21097 2559 21100
rect 2501 21091 2559 21097
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 4706 21088 4712 21140
rect 4764 21128 4770 21140
rect 5445 21131 5503 21137
rect 5445 21128 5457 21131
rect 4764 21100 5457 21128
rect 4764 21088 4770 21100
rect 5445 21097 5457 21100
rect 5491 21097 5503 21131
rect 5445 21091 5503 21097
rect 7282 21088 7288 21140
rect 7340 21128 7346 21140
rect 7650 21128 7656 21140
rect 7340 21100 7656 21128
rect 7340 21088 7346 21100
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 1670 21060 1676 21072
rect 1631 21032 1676 21060
rect 1670 21020 1676 21032
rect 1728 21020 1734 21072
rect 7101 21063 7159 21069
rect 7101 21029 7113 21063
rect 7147 21060 7159 21063
rect 7466 21060 7472 21072
rect 7147 21032 7472 21060
rect 7147 21029 7159 21032
rect 7101 21023 7159 21029
rect 7466 21020 7472 21032
rect 7524 21020 7530 21072
rect 9944 21063 10002 21069
rect 9944 21029 9956 21063
rect 9990 21060 10002 21063
rect 10318 21060 10324 21072
rect 9990 21032 10324 21060
rect 9990 21029 10002 21032
rect 9944 21023 10002 21029
rect 10318 21020 10324 21032
rect 10376 21020 10382 21072
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 4338 21001 4344 21004
rect 4332 20992 4344 21001
rect 4299 20964 4344 20992
rect 4332 20955 4344 20964
rect 4338 20952 4344 20955
rect 4396 20952 4402 21004
rect 6086 20952 6092 21004
rect 6144 20952 6150 21004
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 6972 20964 7205 20992
rect 6972 20952 6978 20964
rect 7193 20961 7205 20964
rect 7239 20961 7251 20995
rect 7193 20955 7251 20961
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 10962 20992 10968 21004
rect 9723 20964 10968 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 3510 20884 3516 20936
rect 3568 20924 3574 20936
rect 3605 20927 3663 20933
rect 3605 20924 3617 20927
rect 3568 20896 3617 20924
rect 3568 20884 3574 20896
rect 3605 20893 3617 20896
rect 3651 20924 3663 20927
rect 4062 20924 4068 20936
rect 3651 20896 4068 20924
rect 3651 20893 3663 20896
rect 3605 20887 3663 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6104 20924 6132 20952
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 5592 20896 6377 20924
rect 5592 20884 5598 20896
rect 6365 20893 6377 20896
rect 6411 20893 6423 20927
rect 7098 20924 7104 20936
rect 7059 20896 7104 20924
rect 6365 20887 6423 20893
rect 7098 20884 7104 20896
rect 7156 20884 7162 20936
rect 6178 20816 6184 20868
rect 6236 20856 6242 20868
rect 6641 20859 6699 20865
rect 6641 20856 6653 20859
rect 6236 20828 6653 20856
rect 6236 20816 6242 20828
rect 6641 20825 6653 20828
rect 6687 20825 6699 20859
rect 6641 20819 6699 20825
rect 5994 20788 6000 20800
rect 5955 20760 6000 20788
rect 5994 20748 6000 20760
rect 6052 20748 6058 20800
rect 8205 20791 8263 20797
rect 8205 20757 8217 20791
rect 8251 20788 8263 20791
rect 8294 20788 8300 20800
rect 8251 20760 8300 20788
rect 8251 20757 8263 20760
rect 8205 20751 8263 20757
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 8573 20791 8631 20797
rect 8573 20788 8585 20791
rect 8536 20760 8585 20788
rect 8536 20748 8542 20760
rect 8573 20757 8585 20760
rect 8619 20788 8631 20791
rect 8754 20788 8760 20800
rect 8619 20760 8760 20788
rect 8619 20757 8631 20760
rect 8573 20751 8631 20757
rect 8754 20748 8760 20760
rect 8812 20788 8818 20800
rect 9398 20788 9404 20800
rect 8812 20760 9404 20788
rect 8812 20748 8818 20760
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 11054 20788 11060 20800
rect 11015 20760 11060 20788
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5534 20584 5540 20596
rect 5307 20556 5540 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 7374 20544 7380 20596
rect 7432 20584 7438 20596
rect 8021 20587 8079 20593
rect 8021 20584 8033 20587
rect 7432 20556 8033 20584
rect 7432 20544 7438 20556
rect 8021 20553 8033 20556
rect 8067 20553 8079 20587
rect 8021 20547 8079 20553
rect 3697 20519 3755 20525
rect 3697 20485 3709 20519
rect 3743 20485 3755 20519
rect 7006 20516 7012 20528
rect 3697 20479 3755 20485
rect 5736 20488 7012 20516
rect 2222 20448 2228 20460
rect 1412 20420 2228 20448
rect 1412 20389 1440 20420
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20349 1455 20383
rect 3712 20380 3740 20479
rect 4062 20408 4068 20460
rect 4120 20448 4126 20460
rect 4614 20448 4620 20460
rect 4120 20420 4620 20448
rect 4120 20408 4126 20420
rect 4614 20408 4620 20420
rect 4672 20408 4678 20460
rect 4706 20408 4712 20460
rect 4764 20448 4770 20460
rect 5736 20457 5764 20488
rect 7006 20476 7012 20488
rect 7064 20476 7070 20528
rect 5721 20451 5779 20457
rect 5721 20448 5733 20451
rect 4764 20420 5733 20448
rect 4764 20408 4770 20420
rect 5721 20417 5733 20420
rect 5767 20417 5779 20451
rect 5721 20411 5779 20417
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20448 6883 20451
rect 7558 20448 7564 20460
rect 6871 20420 7564 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 7558 20408 7564 20420
rect 7616 20408 7622 20460
rect 8036 20448 8064 20547
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 10505 20587 10563 20593
rect 10505 20584 10517 20587
rect 10376 20556 10517 20584
rect 10376 20544 10382 20556
rect 10505 20553 10517 20556
rect 10551 20553 10563 20587
rect 10505 20547 10563 20553
rect 10229 20519 10287 20525
rect 10229 20485 10241 20519
rect 10275 20516 10287 20519
rect 10594 20516 10600 20528
rect 10275 20488 10600 20516
rect 10275 20485 10287 20488
rect 10229 20479 10287 20485
rect 10594 20476 10600 20488
rect 10652 20516 10658 20528
rect 10962 20516 10968 20528
rect 10652 20488 10968 20516
rect 10652 20476 10658 20488
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 8205 20451 8263 20457
rect 8205 20448 8217 20451
rect 8036 20420 8217 20448
rect 8205 20417 8217 20420
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 5994 20380 6000 20392
rect 3712 20352 6000 20380
rect 1397 20343 1455 20349
rect 1670 20312 1676 20324
rect 1631 20284 1676 20312
rect 1670 20272 1676 20284
rect 1728 20272 1734 20324
rect 3513 20315 3571 20321
rect 3513 20281 3525 20315
rect 3559 20312 3571 20315
rect 3878 20312 3884 20324
rect 3559 20284 3884 20312
rect 3559 20281 3571 20284
rect 3513 20275 3571 20281
rect 3878 20272 3884 20284
rect 3936 20312 3942 20324
rect 3973 20315 4031 20321
rect 3973 20312 3985 20315
rect 3936 20284 3985 20312
rect 3936 20272 3942 20284
rect 3973 20281 3985 20284
rect 4019 20281 4031 20315
rect 3973 20275 4031 20281
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 4157 20315 4215 20321
rect 4157 20312 4169 20315
rect 4120 20284 4169 20312
rect 4120 20272 4126 20284
rect 4157 20281 4169 20284
rect 4203 20281 4215 20315
rect 4157 20275 4215 20281
rect 4249 20315 4307 20321
rect 4249 20281 4261 20315
rect 4295 20312 4307 20315
rect 5442 20312 5448 20324
rect 4295 20284 5448 20312
rect 4295 20281 4307 20284
rect 4249 20275 4307 20281
rect 3145 20247 3203 20253
rect 3145 20213 3157 20247
rect 3191 20244 3203 20247
rect 4347 20244 4375 20284
rect 5442 20272 5448 20284
rect 5500 20272 5506 20324
rect 5736 20321 5764 20352
rect 5994 20340 6000 20352
rect 6052 20340 6058 20392
rect 8478 20389 8484 20392
rect 8472 20380 8484 20389
rect 8404 20352 8484 20380
rect 5721 20315 5779 20321
rect 5721 20281 5733 20315
rect 5767 20281 5779 20315
rect 5721 20275 5779 20281
rect 5813 20315 5871 20321
rect 5813 20281 5825 20315
rect 5859 20281 5871 20315
rect 5813 20275 5871 20281
rect 6273 20315 6331 20321
rect 6273 20281 6285 20315
rect 6319 20312 6331 20315
rect 7098 20312 7104 20324
rect 6319 20284 7104 20312
rect 6319 20281 6331 20284
rect 6273 20275 6331 20281
rect 4614 20244 4620 20256
rect 3191 20216 4375 20244
rect 4575 20216 4620 20244
rect 3191 20213 3203 20216
rect 3145 20207 3203 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 5077 20247 5135 20253
rect 5077 20213 5089 20247
rect 5123 20244 5135 20247
rect 5258 20244 5264 20256
rect 5123 20216 5264 20244
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 5258 20204 5264 20216
rect 5316 20244 5322 20256
rect 5828 20244 5856 20275
rect 7098 20272 7104 20284
rect 7156 20272 7162 20324
rect 7745 20315 7803 20321
rect 7745 20281 7757 20315
rect 7791 20312 7803 20315
rect 8404 20312 8432 20352
rect 8472 20343 8484 20352
rect 8478 20340 8484 20343
rect 8536 20340 8542 20392
rect 7791 20284 8432 20312
rect 7791 20281 7803 20284
rect 7745 20275 7803 20281
rect 6641 20247 6699 20253
rect 6641 20244 6653 20247
rect 5316 20216 6653 20244
rect 5316 20204 5322 20216
rect 6641 20213 6653 20216
rect 6687 20244 6699 20247
rect 6822 20244 6828 20256
rect 6687 20216 6828 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7466 20244 7472 20256
rect 7423 20216 7472 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 9582 20244 9588 20256
rect 9543 20216 9588 20244
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 1452 20012 1593 20040
rect 1452 20000 1458 20012
rect 1581 20009 1593 20012
rect 1627 20009 1639 20043
rect 1581 20003 1639 20009
rect 3697 20043 3755 20049
rect 3697 20009 3709 20043
rect 3743 20040 3755 20043
rect 3970 20040 3976 20052
rect 3743 20012 3976 20040
rect 3743 20009 3755 20012
rect 3697 20003 3755 20009
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4338 20040 4344 20052
rect 4251 20012 4344 20040
rect 4338 20000 4344 20012
rect 4396 20040 4402 20052
rect 5902 20040 5908 20052
rect 4396 20012 5908 20040
rect 4396 20000 4402 20012
rect 5902 20000 5908 20012
rect 5960 20040 5966 20052
rect 6181 20043 6239 20049
rect 6181 20040 6193 20043
rect 5960 20012 6193 20040
rect 5960 20000 5966 20012
rect 6181 20009 6193 20012
rect 6227 20009 6239 20043
rect 6181 20003 6239 20009
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6696 20012 6837 20040
rect 6696 20000 6702 20012
rect 6825 20009 6837 20012
rect 6871 20040 6883 20043
rect 7006 20040 7012 20052
rect 6871 20012 7012 20040
rect 6871 20009 6883 20012
rect 6825 20003 6883 20009
rect 7006 20000 7012 20012
rect 7064 20040 7070 20052
rect 9398 20040 9404 20052
rect 7064 20012 7972 20040
rect 9359 20012 9404 20040
rect 7064 20000 7070 20012
rect 4706 19972 4712 19984
rect 4667 19944 4712 19972
rect 4706 19932 4712 19944
rect 4764 19932 4770 19984
rect 5068 19975 5126 19981
rect 5068 19941 5080 19975
rect 5114 19972 5126 19975
rect 5258 19972 5264 19984
rect 5114 19944 5264 19972
rect 5114 19941 5126 19944
rect 5068 19935 5126 19941
rect 5258 19932 5264 19944
rect 5316 19932 5322 19984
rect 5442 19932 5448 19984
rect 5500 19972 5506 19984
rect 6656 19972 6684 20000
rect 7834 19972 7840 19984
rect 5500 19944 6684 19972
rect 7795 19944 7840 19972
rect 5500 19932 5506 19944
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 7944 19981 7972 20012
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12069 20043 12127 20049
rect 12069 20040 12081 20043
rect 12032 20012 12081 20040
rect 12032 20000 12038 20012
rect 12069 20009 12081 20012
rect 12115 20009 12127 20043
rect 12069 20003 12127 20009
rect 7929 19975 7987 19981
rect 7929 19941 7941 19975
rect 7975 19941 7987 19975
rect 7929 19935 7987 19941
rect 10594 19864 10600 19916
rect 10652 19904 10658 19916
rect 10962 19913 10968 19916
rect 10689 19907 10747 19913
rect 10689 19904 10701 19907
rect 10652 19876 10701 19904
rect 10652 19864 10658 19876
rect 10689 19873 10701 19876
rect 10735 19873 10747 19907
rect 10956 19904 10968 19913
rect 10923 19876 10968 19904
rect 10689 19867 10747 19873
rect 10956 19867 10968 19876
rect 10962 19864 10968 19867
rect 11020 19864 11026 19916
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 4801 19839 4859 19845
rect 4801 19836 4813 19839
rect 4764 19808 4813 19836
rect 4764 19796 4770 19808
rect 4801 19805 4813 19808
rect 4847 19805 4859 19839
rect 4801 19799 4859 19805
rect 7837 19839 7895 19845
rect 7837 19805 7849 19839
rect 7883 19836 7895 19839
rect 7926 19836 7932 19848
rect 7883 19808 7932 19836
rect 7883 19805 7895 19808
rect 7837 19799 7895 19805
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 7098 19728 7104 19780
rect 7156 19768 7162 19780
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 7156 19740 7389 19768
rect 7156 19728 7162 19740
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7377 19731 7435 19737
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 5258 19496 5264 19508
rect 5219 19468 5264 19496
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 6638 19496 6644 19508
rect 6551 19468 6644 19496
rect 6638 19456 6644 19468
rect 6696 19496 6702 19508
rect 7926 19496 7932 19508
rect 6696 19468 7932 19496
rect 6696 19456 6702 19468
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 10652 19468 10701 19496
rect 10652 19456 10658 19468
rect 10689 19465 10701 19468
rect 10735 19496 10747 19499
rect 10778 19496 10784 19508
rect 10735 19468 10784 19496
rect 10735 19465 10747 19468
rect 10689 19459 10747 19465
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 4982 19320 4988 19372
rect 5040 19360 5046 19372
rect 5810 19360 5816 19372
rect 5040 19332 5816 19360
rect 5040 19320 5046 19332
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 1946 19252 1952 19304
rect 2004 19292 2010 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 2004 19264 2237 19292
rect 2004 19252 2010 19264
rect 2225 19261 2237 19264
rect 2271 19292 2283 19295
rect 2317 19295 2375 19301
rect 2317 19292 2329 19295
rect 2271 19264 2329 19292
rect 2271 19261 2283 19264
rect 2225 19255 2283 19261
rect 2317 19261 2329 19264
rect 2363 19292 2375 19295
rect 3510 19292 3516 19304
rect 2363 19264 3516 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 3510 19252 3516 19264
rect 3568 19292 3574 19304
rect 4706 19292 4712 19304
rect 3568 19264 4712 19292
rect 3568 19252 3574 19264
rect 4706 19252 4712 19264
rect 4764 19292 4770 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 4764 19264 4905 19292
rect 4764 19252 4770 19264
rect 4893 19261 4905 19264
rect 4939 19292 4951 19295
rect 5534 19292 5540 19304
rect 4939 19264 5540 19292
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 5534 19252 5540 19264
rect 5592 19292 5598 19304
rect 6822 19292 6828 19304
rect 5592 19264 6828 19292
rect 5592 19252 5598 19264
rect 6822 19252 6828 19264
rect 6880 19292 6886 19304
rect 7374 19292 7380 19304
rect 6880 19264 7380 19292
rect 6880 19252 6886 19264
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7834 19252 7840 19304
rect 7892 19292 7898 19304
rect 9383 19295 9441 19301
rect 9383 19292 9395 19295
rect 7892 19264 9395 19292
rect 7892 19252 7898 19264
rect 9383 19261 9395 19264
rect 9429 19261 9441 19295
rect 9383 19255 9441 19261
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9916 19264 9965 19292
rect 9916 19252 9922 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 2590 19233 2596 19236
rect 2584 19224 2596 19233
rect 2551 19196 2596 19224
rect 2584 19187 2596 19196
rect 2590 19184 2596 19187
rect 2648 19184 2654 19236
rect 7006 19184 7012 19236
rect 7064 19233 7070 19236
rect 7064 19227 7128 19233
rect 7064 19193 7082 19227
rect 7116 19224 7128 19227
rect 8757 19227 8815 19233
rect 8757 19224 8769 19227
rect 7116 19196 8769 19224
rect 7116 19193 7128 19196
rect 7064 19187 7128 19193
rect 8757 19193 8769 19196
rect 8803 19224 8815 19227
rect 9582 19224 9588 19236
rect 8803 19196 9588 19224
rect 8803 19193 8815 19196
rect 8757 19187 8815 19193
rect 7064 19184 7070 19187
rect 9582 19184 9588 19196
rect 9640 19184 9646 19236
rect 9674 19184 9680 19236
rect 9732 19224 9738 19236
rect 9732 19196 9777 19224
rect 9732 19184 9738 19196
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 3970 19156 3976 19168
rect 3743 19128 3976 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 8205 19159 8263 19165
rect 8205 19156 8217 19159
rect 6972 19128 8217 19156
rect 6972 19116 6978 19128
rect 8205 19125 8217 19128
rect 8251 19125 8263 19159
rect 8205 19119 8263 19125
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19156 9275 19159
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9263 19128 9873 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9861 19125 9873 19128
rect 9907 19156 9919 19159
rect 10042 19156 10048 19168
rect 9907 19128 10048 19156
rect 9907 19125 9919 19128
rect 9861 19119 9919 19125
rect 10042 19116 10048 19128
rect 10100 19156 10106 19168
rect 10502 19156 10508 19168
rect 10100 19128 10508 19156
rect 10100 19116 10106 19128
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11057 19159 11115 19165
rect 11057 19156 11069 19159
rect 11020 19128 11069 19156
rect 11020 19116 11026 19128
rect 11057 19125 11069 19128
rect 11103 19125 11115 19159
rect 11057 19119 11115 19125
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 4798 18952 4804 18964
rect 4759 18924 4804 18952
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 6822 18952 6828 18964
rect 6783 18924 6828 18952
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 7285 18955 7343 18961
rect 7285 18921 7297 18955
rect 7331 18952 7343 18955
rect 7834 18952 7840 18964
rect 7331 18924 7840 18952
rect 7331 18921 7343 18924
rect 7285 18915 7343 18921
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 9214 18912 9220 18964
rect 9272 18952 9278 18964
rect 9309 18955 9367 18961
rect 9309 18952 9321 18955
rect 9272 18924 9321 18952
rect 9272 18912 9278 18924
rect 9309 18921 9321 18924
rect 9355 18952 9367 18955
rect 9674 18952 9680 18964
rect 9355 18924 9680 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 7742 18884 7748 18896
rect 7703 18856 7748 18884
rect 7742 18844 7748 18856
rect 7800 18844 7806 18896
rect 7926 18884 7932 18896
rect 7887 18856 7932 18884
rect 7926 18844 7932 18856
rect 7984 18844 7990 18896
rect 10226 18884 10232 18896
rect 10187 18856 10232 18884
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 7006 18776 7012 18828
rect 7064 18816 7070 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7064 18788 8033 18816
rect 7064 18776 7070 18788
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 2958 18708 2964 18760
rect 3016 18748 3022 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3016 18720 4077 18748
rect 3016 18708 3022 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 10137 18751 10195 18757
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10137 18711 10195 18717
rect 7466 18680 7472 18692
rect 7427 18652 7472 18680
rect 7466 18640 7472 18652
rect 7524 18640 7530 18692
rect 10152 18680 10180 18711
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 11146 18680 11152 18692
rect 10152 18652 11152 18680
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 2590 18612 2596 18624
rect 2455 18584 2596 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 9769 18615 9827 18621
rect 9769 18612 9781 18615
rect 9732 18584 9781 18612
rect 9732 18572 9738 18584
rect 9769 18581 9781 18584
rect 9815 18581 9827 18615
rect 9769 18575 9827 18581
rect 10594 18572 10600 18624
rect 10652 18612 10658 18624
rect 10962 18612 10968 18624
rect 10652 18584 10968 18612
rect 10652 18572 10658 18584
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 7742 18408 7748 18420
rect 6687 18380 7748 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 9953 18411 10011 18417
rect 9953 18377 9965 18411
rect 9999 18408 10011 18411
rect 10226 18408 10232 18420
rect 9999 18380 10232 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 10226 18368 10232 18380
rect 10284 18408 10290 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 10284 18380 10885 18408
rect 10284 18368 10290 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 11146 18408 11152 18420
rect 11020 18380 11152 18408
rect 11020 18368 11026 18380
rect 11146 18368 11152 18380
rect 11204 18408 11210 18420
rect 11241 18411 11299 18417
rect 11241 18408 11253 18411
rect 11204 18380 11253 18408
rect 11204 18368 11210 18380
rect 11241 18377 11253 18380
rect 11287 18377 11299 18411
rect 11241 18371 11299 18377
rect 1964 18272 1992 18368
rect 4893 18343 4951 18349
rect 4893 18309 4905 18343
rect 4939 18340 4951 18343
rect 5166 18340 5172 18352
rect 4939 18312 5172 18340
rect 4939 18309 4951 18312
rect 4893 18303 4951 18309
rect 5166 18300 5172 18312
rect 5224 18300 5230 18352
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 7285 18343 7343 18349
rect 7285 18340 7297 18343
rect 7064 18312 7297 18340
rect 7064 18300 7070 18312
rect 7285 18309 7297 18312
rect 7331 18309 7343 18343
rect 7285 18303 7343 18309
rect 7466 18300 7472 18352
rect 7524 18340 7530 18352
rect 7926 18340 7932 18352
rect 7524 18312 7932 18340
rect 7524 18300 7530 18312
rect 7926 18300 7932 18312
rect 7984 18340 7990 18352
rect 8297 18343 8355 18349
rect 8297 18340 8309 18343
rect 7984 18312 8309 18340
rect 7984 18300 7990 18312
rect 8297 18309 8309 18312
rect 8343 18309 8355 18343
rect 8297 18303 8355 18309
rect 8754 18300 8760 18352
rect 8812 18340 8818 18352
rect 9306 18340 9312 18352
rect 8812 18312 9312 18340
rect 8812 18300 8818 18312
rect 9306 18300 9312 18312
rect 9364 18300 9370 18352
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 1964 18244 2053 18272
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 4798 18232 4804 18284
rect 4856 18272 4862 18284
rect 5261 18275 5319 18281
rect 5261 18272 5273 18275
rect 4856 18244 5273 18272
rect 4856 18232 4862 18244
rect 5261 18241 5273 18244
rect 5307 18272 5319 18275
rect 7653 18275 7711 18281
rect 7653 18272 7665 18275
rect 5307 18244 7665 18272
rect 5307 18241 5319 18244
rect 5261 18235 5319 18241
rect 7653 18241 7665 18244
rect 7699 18241 7711 18275
rect 7653 18235 7711 18241
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18204 4399 18207
rect 5442 18204 5448 18216
rect 4387 18176 5448 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 5442 18164 5448 18176
rect 5500 18164 5506 18216
rect 7668 18204 7696 18235
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 8849 18275 8907 18281
rect 8849 18272 8861 18275
rect 8536 18244 8861 18272
rect 8536 18232 8542 18244
rect 8849 18241 8861 18244
rect 8895 18241 8907 18275
rect 8849 18235 8907 18241
rect 8573 18207 8631 18213
rect 8573 18204 8585 18207
rect 7668 18176 8585 18204
rect 8496 18148 8524 18176
rect 8573 18173 8585 18176
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 9364 18176 9413 18204
rect 9364 18164 9370 18176
rect 9401 18173 9413 18176
rect 9447 18204 9459 18207
rect 10505 18207 10563 18213
rect 10505 18204 10517 18207
rect 9447 18176 10517 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 10505 18173 10517 18176
rect 10551 18173 10563 18207
rect 10505 18167 10563 18173
rect 1946 18096 1952 18148
rect 2004 18136 2010 18148
rect 2286 18139 2344 18145
rect 2286 18136 2298 18139
rect 2004 18108 2298 18136
rect 2004 18096 2010 18108
rect 2286 18105 2298 18108
rect 2332 18105 2344 18139
rect 2286 18099 2344 18105
rect 4709 18139 4767 18145
rect 4709 18105 4721 18139
rect 4755 18136 4767 18139
rect 5074 18136 5080 18148
rect 4755 18108 5080 18136
rect 4755 18105 4767 18108
rect 4709 18099 4767 18105
rect 5074 18096 5080 18108
rect 5132 18136 5138 18148
rect 5353 18139 5411 18145
rect 5353 18136 5365 18139
rect 5132 18108 5365 18136
rect 5132 18096 5138 18108
rect 5353 18105 5365 18108
rect 5399 18136 5411 18139
rect 8021 18139 8079 18145
rect 8021 18136 8033 18139
rect 5399 18108 8033 18136
rect 5399 18105 5411 18108
rect 5353 18099 5411 18105
rect 8021 18105 8033 18108
rect 8067 18105 8079 18139
rect 8021 18099 8079 18105
rect 2590 18028 2596 18080
rect 2648 18068 2654 18080
rect 3421 18071 3479 18077
rect 3421 18068 3433 18071
rect 2648 18040 3433 18068
rect 2648 18028 2654 18040
rect 3421 18037 3433 18040
rect 3467 18037 3479 18071
rect 8036 18068 8064 18099
rect 8478 18096 8484 18148
rect 8536 18096 8542 18148
rect 8757 18139 8815 18145
rect 8757 18105 8769 18139
rect 8803 18136 8815 18139
rect 10134 18136 10140 18148
rect 8803 18108 10140 18136
rect 8803 18105 8815 18108
rect 8757 18099 8815 18105
rect 8772 18068 8800 18099
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 10229 18139 10287 18145
rect 10229 18105 10241 18139
rect 10275 18105 10287 18139
rect 10229 18099 10287 18105
rect 8036 18040 8800 18068
rect 3421 18031 3479 18037
rect 9490 18028 9496 18080
rect 9548 18068 9554 18080
rect 9677 18071 9735 18077
rect 9677 18068 9689 18071
rect 9548 18040 9689 18068
rect 9548 18028 9554 18040
rect 9677 18037 9689 18040
rect 9723 18068 9735 18071
rect 10244 18068 10272 18099
rect 10410 18068 10416 18080
rect 9723 18040 10272 18068
rect 10371 18040 10416 18068
rect 9723 18037 9735 18040
rect 9677 18031 9735 18037
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 5353 17867 5411 17873
rect 5353 17833 5365 17867
rect 5399 17864 5411 17867
rect 5718 17864 5724 17876
rect 5399 17836 5724 17864
rect 5399 17833 5411 17836
rect 5353 17827 5411 17833
rect 5718 17824 5724 17836
rect 5776 17824 5782 17876
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 9861 17867 9919 17873
rect 9861 17864 9873 17867
rect 9824 17836 9873 17864
rect 9824 17824 9830 17836
rect 9861 17833 9873 17836
rect 9907 17864 9919 17867
rect 10410 17864 10416 17876
rect 9907 17836 10416 17864
rect 9907 17833 9919 17836
rect 9861 17827 9919 17833
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 10652 17836 12265 17864
rect 10652 17824 10658 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 12253 17827 12311 17833
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 2961 17799 3019 17805
rect 2961 17796 2973 17799
rect 2924 17768 2973 17796
rect 2924 17756 2930 17768
rect 2961 17765 2973 17768
rect 3007 17765 3019 17799
rect 2961 17759 3019 17765
rect 5442 17756 5448 17808
rect 5500 17796 5506 17808
rect 8570 17796 8576 17808
rect 5500 17768 5545 17796
rect 8531 17768 8576 17796
rect 5500 17756 5506 17768
rect 8570 17756 8576 17768
rect 8628 17756 8634 17808
rect 1946 17688 1952 17740
rect 2004 17728 2010 17740
rect 2004 17700 3096 17728
rect 2004 17688 2010 17700
rect 3068 17672 3096 17700
rect 5074 17688 5080 17740
rect 5132 17728 5138 17740
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 5132 17700 5181 17728
rect 5132 17688 5138 17700
rect 5169 17697 5181 17700
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7432 17700 8401 17728
rect 7432 17688 7438 17700
rect 8389 17697 8401 17700
rect 8435 17728 8447 17731
rect 9582 17728 9588 17740
rect 8435 17700 9588 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10318 17728 10324 17740
rect 9916 17700 10324 17728
rect 9916 17688 9922 17700
rect 10318 17688 10324 17700
rect 10376 17728 10382 17740
rect 10781 17731 10839 17737
rect 10781 17728 10793 17731
rect 10376 17700 10793 17728
rect 10376 17688 10382 17700
rect 10781 17697 10793 17700
rect 10827 17728 10839 17731
rect 11140 17731 11198 17737
rect 11140 17728 11152 17731
rect 10827 17700 11152 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 11140 17697 11152 17700
rect 11186 17728 11198 17731
rect 12158 17728 12164 17740
rect 11186 17700 12164 17728
rect 11186 17697 11198 17700
rect 11140 17691 11198 17697
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 3050 17620 3056 17672
rect 3108 17660 3114 17672
rect 8662 17660 8668 17672
rect 3108 17632 3153 17660
rect 8623 17632 8668 17660
rect 3108 17620 3114 17632
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 1765 17595 1823 17601
rect 1765 17561 1777 17595
rect 1811 17592 1823 17595
rect 2222 17592 2228 17604
rect 1811 17564 2228 17592
rect 1811 17561 1823 17564
rect 1765 17555 1823 17561
rect 2222 17552 2228 17564
rect 2280 17592 2286 17604
rect 2590 17592 2596 17604
rect 2280 17564 2596 17592
rect 2280 17552 2286 17564
rect 2590 17552 2596 17564
rect 2648 17552 2654 17604
rect 10778 17552 10784 17604
rect 10836 17592 10842 17604
rect 10888 17592 10916 17623
rect 10836 17564 10916 17592
rect 10836 17552 10842 17564
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2041 17527 2099 17533
rect 2041 17524 2053 17527
rect 2004 17496 2053 17524
rect 2004 17484 2010 17496
rect 2041 17493 2053 17496
rect 2087 17493 2099 17527
rect 2498 17524 2504 17536
rect 2459 17496 2504 17524
rect 2041 17487 2099 17493
rect 2498 17484 2504 17496
rect 2556 17484 2562 17536
rect 4893 17527 4951 17533
rect 4893 17493 4905 17527
rect 4939 17524 4951 17527
rect 4982 17524 4988 17536
rect 4939 17496 4988 17524
rect 4939 17493 4951 17496
rect 4893 17487 4951 17493
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 6972 17496 8125 17524
rect 6972 17484 6978 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9766 17524 9772 17536
rect 9355 17496 9772 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 1946 17320 1952 17332
rect 1719 17292 1952 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2041 17323 2099 17329
rect 2041 17289 2053 17323
rect 2087 17320 2099 17323
rect 2958 17320 2964 17332
rect 2087 17292 2964 17320
rect 2087 17289 2099 17292
rect 2041 17283 2099 17289
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 3510 17320 3516 17332
rect 3471 17292 3516 17320
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 5077 17323 5135 17329
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 5442 17320 5448 17332
rect 5123 17292 5448 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7745 17323 7803 17329
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 8570 17320 8576 17332
rect 7791 17292 8576 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 8570 17280 8576 17292
rect 8628 17320 8634 17332
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 8628 17292 9321 17320
rect 8628 17280 8634 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 9309 17283 9367 17289
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 10962 17320 10968 17332
rect 10919 17292 10968 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 2225 17255 2283 17261
rect 2225 17221 2237 17255
rect 2271 17221 2283 17255
rect 2225 17215 2283 17221
rect 2038 17144 2044 17196
rect 2096 17184 2102 17196
rect 2240 17184 2268 17215
rect 2590 17184 2596 17196
rect 2096 17156 2596 17184
rect 2096 17144 2102 17156
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 3528 17184 3556 17280
rect 8113 17255 8171 17261
rect 8113 17221 8125 17255
rect 8159 17252 8171 17255
rect 8662 17252 8668 17264
rect 8159 17224 8668 17252
rect 8159 17221 8171 17224
rect 8113 17215 8171 17221
rect 8662 17212 8668 17224
rect 8720 17212 8726 17264
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3528 17156 3709 17184
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 8202 17184 8208 17196
rect 7248 17156 8208 17184
rect 7248 17144 7254 17156
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9858 17184 9864 17196
rect 9171 17156 9864 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 2498 17116 2504 17128
rect 2459 17088 2504 17116
rect 2498 17076 2504 17088
rect 2556 17076 2562 17128
rect 3970 17125 3976 17128
rect 3964 17116 3976 17125
rect 3931 17088 3976 17116
rect 3964 17079 3976 17088
rect 3970 17076 3976 17079
rect 4028 17076 4034 17128
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11195 17088 11928 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 2222 17008 2228 17060
rect 2280 17048 2286 17060
rect 2777 17051 2835 17057
rect 2777 17048 2789 17051
rect 2280 17020 2789 17048
rect 2280 17008 2286 17020
rect 2777 17017 2789 17020
rect 2823 17017 2835 17051
rect 2777 17011 2835 17017
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 5350 17048 5356 17060
rect 3016 17020 5356 17048
rect 3016 17008 3022 17020
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 9398 17048 9404 17060
rect 8803 17020 9404 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 9398 17008 9404 17020
rect 9456 17048 9462 17060
rect 9585 17051 9643 17057
rect 9585 17048 9597 17051
rect 9456 17020 9597 17048
rect 9456 17008 9462 17020
rect 9585 17017 9597 17020
rect 9631 17017 9643 17051
rect 9766 17048 9772 17060
rect 9727 17020 9772 17048
rect 9585 17011 9643 17017
rect 9766 17008 9772 17020
rect 9824 17008 9830 17060
rect 10321 17051 10379 17057
rect 10321 17017 10333 17051
rect 10367 17048 10379 17051
rect 10778 17048 10784 17060
rect 10367 17020 10784 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 11422 17048 11428 17060
rect 11383 17020 11428 17048
rect 11422 17008 11428 17020
rect 11480 17008 11486 17060
rect 11900 17057 11928 17088
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12437 17051 12495 17057
rect 12437 17048 12449 17051
rect 11931 17020 12449 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12437 17017 12449 17020
rect 12483 17017 12495 17051
rect 12437 17011 12495 17017
rect 2682 16980 2688 16992
rect 2643 16952 2688 16980
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 3145 16983 3203 16989
rect 3145 16980 3157 16983
rect 2924 16952 3157 16980
rect 2924 16940 2930 16952
rect 3145 16949 3157 16952
rect 3191 16949 3203 16983
rect 5718 16980 5724 16992
rect 5679 16952 5724 16980
rect 3145 16943 3203 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 10686 16980 10692 16992
rect 10647 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16980 10750 16992
rect 11333 16983 11391 16989
rect 11333 16980 11345 16983
rect 10744 16952 11345 16980
rect 10744 16940 10750 16952
rect 11333 16949 11345 16952
rect 11379 16949 11391 16983
rect 11440 16980 11468 17008
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11440 16952 12173 16980
rect 11333 16943 11391 16949
rect 12161 16949 12173 16952
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 1673 16779 1731 16785
rect 1673 16745 1685 16779
rect 1719 16776 1731 16779
rect 2682 16776 2688 16788
rect 1719 16748 2688 16776
rect 1719 16745 1731 16748
rect 1673 16739 1731 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 3789 16779 3847 16785
rect 3789 16745 3801 16779
rect 3835 16776 3847 16779
rect 3970 16776 3976 16788
rect 3835 16748 3976 16776
rect 3835 16745 3847 16748
rect 3789 16739 3847 16745
rect 2130 16668 2136 16720
rect 2188 16708 2194 16720
rect 2317 16711 2375 16717
rect 2317 16708 2329 16711
rect 2188 16680 2329 16708
rect 2188 16668 2194 16680
rect 2317 16677 2329 16680
rect 2363 16677 2375 16711
rect 3804 16708 3832 16739
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 5442 16776 5448 16788
rect 4396 16748 5448 16776
rect 4396 16736 4402 16748
rect 4614 16708 4620 16720
rect 2317 16671 2375 16677
rect 2424 16680 3832 16708
rect 4575 16680 4620 16708
rect 2038 16600 2044 16652
rect 2096 16640 2102 16652
rect 2096 16612 2268 16640
rect 2096 16600 2102 16612
rect 2240 16581 2268 16612
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2314 16532 2320 16584
rect 2372 16572 2378 16584
rect 2424 16581 2452 16680
rect 4614 16668 4620 16680
rect 4672 16668 4678 16720
rect 4724 16717 4752 16748
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 9306 16776 9312 16788
rect 9267 16748 9312 16776
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 12158 16776 12164 16788
rect 12119 16748 12164 16776
rect 12158 16736 12164 16748
rect 12216 16736 12222 16788
rect 4709 16711 4767 16717
rect 4709 16677 4721 16711
rect 4755 16677 4767 16711
rect 5074 16708 5080 16720
rect 5035 16680 5080 16708
rect 4709 16671 4767 16677
rect 5074 16668 5080 16680
rect 5132 16668 5138 16720
rect 5460 16708 5488 16736
rect 5874 16711 5932 16717
rect 5874 16708 5886 16711
rect 5460 16680 5886 16708
rect 5874 16677 5886 16680
rect 5920 16708 5932 16711
rect 5994 16708 6000 16720
rect 5920 16680 6000 16708
rect 5920 16677 5932 16680
rect 5874 16671 5932 16677
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 2590 16600 2596 16652
rect 2648 16640 2654 16652
rect 4430 16640 4436 16652
rect 2648 16612 2728 16640
rect 4391 16612 4436 16640
rect 2648 16600 2654 16612
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 2372 16544 2421 16572
rect 2372 16532 2378 16544
rect 2409 16541 2421 16544
rect 2455 16541 2467 16575
rect 2700 16572 2728 16612
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 5592 16612 5641 16640
rect 5592 16600 5598 16612
rect 5629 16609 5641 16612
rect 5675 16609 5687 16643
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 5629 16603 5687 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 9324 16640 9352 16736
rect 11037 16643 11095 16649
rect 11037 16640 11049 16643
rect 9324 16612 9628 16640
rect 3418 16572 3424 16584
rect 2700 16544 3424 16572
rect 2409 16535 2467 16541
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 9600 16572 9628 16612
rect 10704 16612 11049 16640
rect 9950 16572 9956 16584
rect 9600 16544 9956 16572
rect 9950 16532 9956 16544
rect 10008 16572 10014 16584
rect 10704 16572 10732 16612
rect 11037 16609 11049 16612
rect 11083 16640 11095 16643
rect 11422 16640 11428 16652
rect 11083 16612 11428 16640
rect 11083 16609 11095 16612
rect 11037 16603 11095 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 10008 16544 10732 16572
rect 10008 16532 10014 16544
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 10836 16544 10881 16572
rect 10836 16532 10842 16544
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 1857 16439 1915 16445
rect 1857 16436 1869 16439
rect 1820 16408 1869 16436
rect 1820 16396 1826 16408
rect 1857 16405 1869 16408
rect 1903 16405 1915 16439
rect 1857 16399 1915 16405
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3145 16439 3203 16445
rect 3145 16436 3157 16439
rect 3108 16408 3157 16436
rect 3108 16396 3114 16408
rect 3145 16405 3157 16408
rect 3191 16436 3203 16439
rect 3510 16436 3516 16448
rect 3191 16408 3516 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 4154 16436 4160 16448
rect 4115 16408 4160 16436
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 5316 16408 7021 16436
rect 5316 16396 5322 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7650 16436 7656 16448
rect 7611 16408 7656 16436
rect 7009 16399 7067 16405
rect 7650 16396 7656 16408
rect 7708 16396 7714 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 2225 16235 2283 16241
rect 2225 16201 2237 16235
rect 2271 16232 2283 16235
rect 2314 16232 2320 16244
rect 2271 16204 2320 16232
rect 2271 16201 2283 16204
rect 2225 16195 2283 16201
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 2498 16232 2504 16244
rect 2459 16204 2504 16232
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 3145 16235 3203 16241
rect 3145 16232 3157 16235
rect 2832 16204 3157 16232
rect 2832 16192 2838 16204
rect 3145 16201 3157 16204
rect 3191 16201 3203 16235
rect 3145 16195 3203 16201
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4246 16232 4252 16244
rect 4203 16204 4252 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4246 16192 4252 16204
rect 4304 16232 4310 16244
rect 4614 16232 4620 16244
rect 4304 16204 4620 16232
rect 4304 16192 4310 16204
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 5592 16204 5641 16232
rect 5592 16192 5598 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 5994 16232 6000 16244
rect 5955 16204 6000 16232
rect 5629 16195 5687 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 9398 16232 9404 16244
rect 9359 16204 9404 16232
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 11241 16235 11299 16241
rect 11241 16201 11253 16235
rect 11287 16232 11299 16235
rect 11422 16232 11428 16244
rect 11287 16204 11428 16232
rect 11287 16201 11299 16204
rect 11241 16195 11299 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 4709 16167 4767 16173
rect 4709 16133 4721 16167
rect 4755 16164 4767 16167
rect 4798 16164 4804 16176
rect 4755 16136 4804 16164
rect 4755 16133 4767 16136
rect 4709 16127 4767 16133
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 7374 16164 7380 16176
rect 7335 16136 7380 16164
rect 7374 16124 7380 16136
rect 7432 16124 7438 16176
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16096 3019 16099
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 3007 16068 3617 16096
rect 3007 16065 3019 16068
rect 2961 16059 3019 16065
rect 3605 16065 3617 16068
rect 3651 16096 3663 16099
rect 4062 16096 4068 16108
rect 3651 16068 4068 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 5258 16096 5264 16108
rect 5219 16068 5264 16096
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 7834 16096 7840 16108
rect 7747 16068 7840 16096
rect 7834 16056 7840 16068
rect 7892 16096 7898 16108
rect 8297 16099 8355 16105
rect 8297 16096 8309 16099
rect 7892 16068 8309 16096
rect 7892 16056 7898 16068
rect 8297 16065 8309 16068
rect 8343 16065 8355 16099
rect 9950 16096 9956 16108
rect 9911 16068 9956 16096
rect 8297 16059 8355 16065
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 4982 16028 4988 16040
rect 4943 16000 4988 16028
rect 4982 15988 4988 16000
rect 5040 16028 5046 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 5040 16000 6377 16028
rect 5040 15988 5046 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 16028 7251 16031
rect 7926 16028 7932 16040
rect 7239 16000 7932 16028
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 7926 15988 7932 16000
rect 7984 16028 7990 16040
rect 8478 16028 8484 16040
rect 7984 16000 8484 16028
rect 7984 15988 7990 16000
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 3510 15920 3516 15972
rect 3568 15960 3574 15972
rect 3697 15963 3755 15969
rect 3697 15960 3709 15963
rect 3568 15932 3709 15960
rect 3568 15920 3574 15932
rect 3697 15929 3709 15932
rect 3743 15929 3755 15963
rect 5166 15960 5172 15972
rect 5127 15932 5172 15960
rect 3697 15923 3755 15929
rect 5166 15920 5172 15932
rect 5224 15920 5230 15972
rect 7650 15920 7656 15972
rect 7708 15960 7714 15972
rect 7837 15963 7895 15969
rect 7837 15960 7849 15963
rect 7708 15932 7849 15960
rect 7708 15920 7714 15932
rect 7837 15929 7849 15932
rect 7883 15929 7895 15963
rect 7837 15923 7895 15929
rect 9217 15963 9275 15969
rect 9217 15929 9229 15963
rect 9263 15960 9275 15963
rect 9677 15963 9735 15969
rect 9677 15960 9689 15963
rect 9263 15932 9689 15960
rect 9263 15929 9275 15932
rect 9217 15923 9275 15929
rect 9677 15929 9689 15932
rect 9723 15960 9735 15963
rect 10042 15960 10048 15972
rect 9723 15932 10048 15960
rect 9723 15929 9735 15932
rect 9677 15923 9735 15929
rect 10042 15920 10048 15932
rect 10100 15960 10106 15972
rect 10226 15960 10232 15972
rect 10100 15932 10232 15960
rect 10100 15920 10106 15932
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 3602 15892 3608 15904
rect 3563 15864 3608 15892
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 4430 15892 4436 15904
rect 4391 15864 4436 15892
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 9398 15892 9404 15904
rect 8352 15864 9404 15892
rect 8352 15852 8358 15864
rect 9398 15852 9404 15864
rect 9456 15892 9462 15904
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9456 15864 9873 15892
rect 9456 15852 9462 15864
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 9861 15855 9919 15861
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10836 15864 10885 15892
rect 10836 15852 10842 15864
rect 10873 15861 10885 15864
rect 10919 15892 10931 15895
rect 11054 15892 11060 15904
rect 10919 15864 11060 15892
rect 10919 15861 10931 15864
rect 10873 15855 10931 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 3418 15688 3424 15700
rect 3379 15660 3424 15688
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 4338 15688 4344 15700
rect 4299 15660 4344 15688
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 5166 15648 5172 15700
rect 5224 15688 5230 15700
rect 5353 15691 5411 15697
rect 5353 15688 5365 15691
rect 5224 15660 5365 15688
rect 5224 15648 5230 15660
rect 5353 15657 5365 15660
rect 5399 15657 5411 15691
rect 8478 15688 8484 15700
rect 8439 15660 8484 15688
rect 5353 15651 5411 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 1578 15580 1584 15632
rect 1636 15620 1642 15632
rect 2593 15623 2651 15629
rect 2593 15620 2605 15623
rect 1636 15592 2605 15620
rect 1636 15580 1642 15592
rect 2593 15589 2605 15592
rect 2639 15589 2651 15623
rect 2593 15583 2651 15589
rect 3145 15623 3203 15629
rect 3145 15589 3157 15623
rect 3191 15620 3203 15623
rect 3602 15620 3608 15632
rect 3191 15592 3608 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 3602 15580 3608 15592
rect 3660 15580 3666 15632
rect 4709 15623 4767 15629
rect 4709 15589 4721 15623
rect 4755 15620 4767 15623
rect 5077 15623 5135 15629
rect 5077 15620 5089 15623
rect 4755 15592 5089 15620
rect 4755 15589 4767 15592
rect 4709 15583 4767 15589
rect 5077 15589 5089 15592
rect 5123 15620 5135 15623
rect 5258 15620 5264 15632
rect 5123 15592 5264 15620
rect 5123 15589 5135 15592
rect 5077 15583 5135 15589
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 10229 15623 10287 15629
rect 10229 15589 10241 15623
rect 10275 15620 10287 15623
rect 10410 15620 10416 15632
rect 10275 15592 10416 15620
rect 10275 15589 10287 15592
rect 10229 15583 10287 15589
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7368 15555 7426 15561
rect 7368 15552 7380 15555
rect 6972 15524 7380 15552
rect 6972 15512 6978 15524
rect 7368 15521 7380 15524
rect 7414 15552 7426 15555
rect 8202 15552 8208 15564
rect 7414 15524 8208 15552
rect 7414 15521 7426 15524
rect 7368 15515 7426 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 11514 15561 11520 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10008 15524 10333 15552
rect 10008 15512 10014 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 11508 15515 11520 15561
rect 11572 15552 11578 15564
rect 11572 15524 11608 15552
rect 11514 15512 11520 15515
rect 11572 15512 11578 15524
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2682 15484 2688 15496
rect 2643 15456 2688 15484
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 5902 15484 5908 15496
rect 5592 15456 5908 15484
rect 5592 15444 5598 15456
rect 5902 15444 5908 15456
rect 5960 15484 5966 15496
rect 7006 15484 7012 15496
rect 5960 15456 7012 15484
rect 5960 15444 5966 15456
rect 7006 15444 7012 15456
rect 7064 15484 7070 15496
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 7064 15456 7113 15484
rect 7064 15444 7070 15456
rect 7101 15453 7113 15456
rect 7147 15453 7159 15487
rect 7101 15447 7159 15453
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10042 15484 10048 15496
rect 9732 15456 10048 15484
rect 9732 15444 9738 15456
rect 10042 15444 10048 15456
rect 10100 15484 10106 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 10100 15456 10149 15484
rect 10100 15444 10106 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 11112 15456 11253 15484
rect 11112 15444 11118 15456
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 1857 15419 1915 15425
rect 1857 15385 1869 15419
rect 1903 15416 1915 15419
rect 2130 15416 2136 15428
rect 1903 15388 2136 15416
rect 1903 15385 1915 15388
rect 1857 15379 1915 15385
rect 2130 15376 2136 15388
rect 2188 15376 2194 15428
rect 9766 15416 9772 15428
rect 9727 15388 9772 15416
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 9398 15348 9404 15360
rect 9359 15320 9404 15348
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12621 15351 12679 15357
rect 12621 15348 12633 15351
rect 12492 15320 12633 15348
rect 12492 15308 12498 15320
rect 12621 15317 12633 15320
rect 12667 15317 12679 15351
rect 12621 15311 12679 15317
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 2222 15144 2228 15156
rect 2179 15116 2228 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 2222 15104 2228 15116
rect 2280 15144 2286 15156
rect 2682 15144 2688 15156
rect 2280 15116 2688 15144
rect 2280 15104 2286 15116
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 7101 15147 7159 15153
rect 7101 15144 7113 15147
rect 7064 15116 7113 15144
rect 7064 15104 7070 15116
rect 7101 15113 7113 15116
rect 7147 15113 7159 15147
rect 7834 15144 7840 15156
rect 7795 15116 7840 15144
rect 7101 15107 7159 15113
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 10008 15116 10057 15144
rect 10008 15104 10014 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 10045 15107 10103 15113
rect 11514 15104 11520 15156
rect 11572 15144 11578 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 11572 15116 11621 15144
rect 11572 15104 11578 15116
rect 11609 15113 11621 15116
rect 11655 15113 11667 15147
rect 11609 15107 11667 15113
rect 2498 15036 2504 15088
rect 2556 15076 2562 15088
rect 2774 15076 2780 15088
rect 2556 15048 2780 15076
rect 2556 15036 2562 15048
rect 2774 15036 2780 15048
rect 2832 15076 2838 15088
rect 2961 15079 3019 15085
rect 2961 15076 2973 15079
rect 2832 15048 2973 15076
rect 2832 15036 2838 15048
rect 2961 15045 2973 15048
rect 3007 15045 3019 15079
rect 2961 15039 3019 15045
rect 4709 15079 4767 15085
rect 4709 15045 4721 15079
rect 4755 15076 4767 15079
rect 4982 15076 4988 15088
rect 4755 15048 4988 15076
rect 4755 15045 4767 15048
rect 4709 15039 4767 15045
rect 4982 15036 4988 15048
rect 5040 15036 5046 15088
rect 5350 15076 5356 15088
rect 5092 15048 5356 15076
rect 3418 15008 3424 15020
rect 2792 14980 3424 15008
rect 2792 14949 2820 14980
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 5092 15017 5120 15048
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4571 14980 5089 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 5077 14977 5089 14980
rect 5123 14977 5135 15011
rect 5258 15008 5264 15020
rect 5219 14980 5264 15008
rect 5077 14971 5135 14977
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3510 14940 3516 14952
rect 3200 14912 3516 14940
rect 3200 14900 3206 14912
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 5629 14943 5687 14949
rect 5629 14940 5641 14943
rect 4212 14912 5641 14940
rect 4212 14900 4218 14912
rect 5184 14881 5212 14912
rect 5629 14909 5641 14912
rect 5675 14909 5687 14943
rect 8110 14940 8116 14952
rect 8071 14912 8116 14940
rect 5629 14903 5687 14909
rect 8110 14900 8116 14912
rect 8168 14940 8174 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8168 14912 8769 14940
rect 8168 14900 8174 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 5169 14875 5227 14881
rect 5169 14841 5181 14875
rect 5215 14841 5227 14875
rect 5169 14835 5227 14841
rect 6822 14832 6828 14884
rect 6880 14872 6886 14884
rect 6880 14844 7696 14872
rect 6880 14832 6886 14844
rect 1578 14764 1584 14816
rect 1636 14804 1642 14816
rect 1673 14807 1731 14813
rect 1673 14804 1685 14807
rect 1636 14776 1685 14804
rect 1636 14764 1642 14776
rect 1673 14773 1685 14776
rect 1719 14773 1731 14807
rect 3418 14804 3424 14816
rect 3379 14776 3424 14804
rect 1673 14767 1731 14773
rect 3418 14764 3424 14776
rect 3476 14804 3482 14816
rect 3881 14807 3939 14813
rect 3881 14804 3893 14807
rect 3476 14776 3893 14804
rect 3476 14764 3482 14776
rect 3881 14773 3893 14776
rect 3927 14773 3939 14807
rect 3881 14767 3939 14773
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6178 14804 6184 14816
rect 5868 14776 6184 14804
rect 5868 14764 5874 14776
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 7668 14813 7696 14844
rect 8202 14832 8208 14884
rect 8260 14872 8266 14884
rect 8389 14875 8447 14881
rect 8389 14872 8401 14875
rect 8260 14844 8401 14872
rect 8260 14832 8266 14844
rect 8389 14841 8401 14844
rect 8435 14872 8447 14875
rect 8478 14872 8484 14884
rect 8435 14844 8484 14872
rect 8435 14841 8447 14844
rect 8389 14835 8447 14841
rect 8478 14832 8484 14844
rect 8536 14872 8542 14884
rect 9125 14875 9183 14881
rect 9125 14872 9137 14875
rect 8536 14844 9137 14872
rect 8536 14832 8542 14844
rect 9125 14841 9137 14844
rect 9171 14841 9183 14875
rect 9125 14835 9183 14841
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 7699 14776 8309 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 8297 14773 8309 14776
rect 8343 14804 8355 14807
rect 8754 14804 8760 14816
rect 8343 14776 8760 14804
rect 8343 14773 8355 14776
rect 8297 14767 8355 14773
rect 8754 14764 8760 14776
rect 8812 14764 8818 14816
rect 9769 14807 9827 14813
rect 9769 14773 9781 14807
rect 9815 14804 9827 14807
rect 10042 14804 10048 14816
rect 9815 14776 10048 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10410 14804 10416 14816
rect 10371 14776 10416 14804
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 11112 14776 11253 14804
rect 11112 14764 11118 14776
rect 11241 14773 11253 14776
rect 11287 14773 11299 14807
rect 11241 14767 11299 14773
rect 11514 14764 11520 14816
rect 11572 14804 11578 14816
rect 12618 14804 12624 14816
rect 11572 14776 12624 14804
rect 11572 14764 11578 14776
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 1452 14572 1593 14600
rect 1452 14560 1458 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 1581 14563 1639 14569
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2774 14600 2780 14612
rect 2179 14572 2780 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 5626 14560 5632 14612
rect 5684 14600 5690 14612
rect 6178 14600 6184 14612
rect 5684 14572 6184 14600
rect 5684 14560 5690 14572
rect 6178 14560 6184 14572
rect 6236 14600 6242 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6236 14572 6653 14600
rect 6236 14560 6242 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 6641 14563 6699 14569
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 7432 14572 7481 14600
rect 7432 14560 7438 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8352 14572 8401 14600
rect 8352 14560 8358 14572
rect 8389 14569 8401 14572
rect 8435 14600 8447 14603
rect 8846 14600 8852 14612
rect 8435 14572 8852 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 12676 14572 13461 14600
rect 12676 14560 12682 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13449 14563 13507 14569
rect 1486 14492 1492 14544
rect 1544 14532 1550 14544
rect 3234 14532 3240 14544
rect 1544 14504 3240 14532
rect 1544 14492 1550 14504
rect 3234 14492 3240 14504
rect 3292 14492 3298 14544
rect 4798 14492 4804 14544
rect 4856 14532 4862 14544
rect 5077 14535 5135 14541
rect 5077 14532 5089 14535
rect 4856 14504 5089 14532
rect 4856 14492 4862 14504
rect 5077 14501 5089 14504
rect 5123 14501 5135 14535
rect 5077 14495 5135 14501
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 5534 14532 5540 14544
rect 5316 14504 5540 14532
rect 5316 14492 5322 14504
rect 5534 14492 5540 14504
rect 5592 14532 5598 14544
rect 5905 14535 5963 14541
rect 5905 14532 5917 14535
rect 5592 14504 5917 14532
rect 5592 14492 5598 14504
rect 5905 14501 5917 14504
rect 5951 14532 5963 14535
rect 6733 14535 6791 14541
rect 6733 14532 6745 14535
rect 5951 14504 6745 14532
rect 5951 14501 5963 14504
rect 5905 14495 5963 14501
rect 6733 14501 6745 14504
rect 6779 14501 6791 14535
rect 6733 14495 6791 14501
rect 8018 14492 8024 14544
rect 8076 14532 8082 14544
rect 8205 14535 8263 14541
rect 8205 14532 8217 14535
rect 8076 14504 8217 14532
rect 8076 14492 8082 14504
rect 8205 14501 8217 14504
rect 8251 14532 8263 14535
rect 8570 14532 8576 14544
rect 8251 14504 8576 14532
rect 8251 14501 8263 14504
rect 8205 14495 8263 14501
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 8662 14492 8668 14544
rect 8720 14532 8726 14544
rect 9674 14532 9680 14544
rect 8720 14504 9680 14532
rect 8720 14492 8726 14504
rect 9674 14492 9680 14504
rect 9732 14532 9738 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9732 14504 10057 14532
rect 9732 14492 9738 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 12342 14541 12348 14544
rect 10229 14535 10287 14541
rect 10229 14532 10241 14535
rect 10192 14504 10241 14532
rect 10192 14492 10198 14504
rect 10229 14501 10241 14504
rect 10275 14501 10287 14535
rect 12336 14532 12348 14541
rect 12303 14504 12348 14532
rect 10229 14495 10287 14501
rect 12336 14495 12348 14504
rect 12342 14492 12348 14495
rect 12400 14492 12406 14544
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 12066 14464 12072 14476
rect 11112 14436 12072 14464
rect 11112 14424 11118 14436
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 4982 14396 4988 14408
rect 4943 14368 4988 14396
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 5166 14396 5172 14408
rect 5127 14368 5172 14396
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 6638 14396 6644 14408
rect 6599 14368 6644 14396
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 5629 14331 5687 14337
rect 5629 14297 5641 14331
rect 5675 14328 5687 14331
rect 5718 14328 5724 14340
rect 5675 14300 5724 14328
rect 5675 14297 5687 14300
rect 5629 14291 5687 14297
rect 5718 14288 5724 14300
rect 5776 14328 5782 14340
rect 6181 14331 6239 14337
rect 6181 14328 6193 14331
rect 5776 14300 6193 14328
rect 5776 14288 5782 14300
rect 6181 14297 6193 14300
rect 6227 14297 6239 14331
rect 6181 14291 6239 14297
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 7929 14331 7987 14337
rect 7929 14328 7941 14331
rect 7708 14300 7941 14328
rect 7708 14288 7714 14300
rect 7929 14297 7941 14300
rect 7975 14297 7987 14331
rect 7929 14291 7987 14297
rect 9769 14331 9827 14337
rect 9769 14297 9781 14331
rect 9815 14328 9827 14331
rect 10410 14328 10416 14340
rect 9815 14300 10416 14328
rect 9815 14297 9827 14300
rect 9769 14291 9827 14297
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 2961 14263 3019 14269
rect 2961 14229 2973 14263
rect 3007 14260 3019 14263
rect 3142 14260 3148 14272
rect 3007 14232 3148 14260
rect 3007 14229 3019 14232
rect 2961 14223 3019 14229
rect 3142 14220 3148 14232
rect 3200 14220 3206 14272
rect 4614 14260 4620 14272
rect 4575 14232 4620 14260
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7466 14260 7472 14272
rect 7239 14232 7472 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 3418 14056 3424 14068
rect 3375 14028 3424 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 8662 14056 8668 14068
rect 8352 14028 8668 14056
rect 8352 14016 8358 14028
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 8812 14028 9321 14056
rect 8812 14016 8818 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 9766 14056 9772 14068
rect 9679 14028 9772 14056
rect 9309 14019 9367 14025
rect 9766 14016 9772 14028
rect 9824 14056 9830 14068
rect 10134 14056 10140 14068
rect 9824 14028 10140 14056
rect 9824 14016 9830 14028
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 11241 14059 11299 14065
rect 11241 14025 11253 14059
rect 11287 14056 11299 14059
rect 11422 14056 11428 14068
rect 11287 14028 11428 14056
rect 11287 14025 11299 14028
rect 11241 14019 11299 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12342 14056 12348 14068
rect 12207 14028 12348 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 5258 13988 5264 14000
rect 5219 13960 5264 13988
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 2222 13920 2228 13932
rect 1412 13892 2228 13920
rect 1412 13861 1440 13892
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 3881 13923 3939 13929
rect 3881 13920 3893 13923
rect 2832 13892 3893 13920
rect 2832 13880 2838 13892
rect 3881 13889 3893 13892
rect 3927 13889 3939 13923
rect 5718 13920 5724 13932
rect 5679 13892 5724 13920
rect 3881 13883 3939 13889
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 6196 13864 6224 14016
rect 7006 13988 7012 14000
rect 6967 13960 7012 13988
rect 7006 13948 7012 13960
rect 7064 13948 7070 14000
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 12621 13991 12679 13997
rect 12621 13988 12633 13991
rect 12124 13960 12633 13988
rect 12124 13948 12130 13960
rect 12621 13957 12633 13960
rect 12667 13957 12679 13991
rect 12621 13951 12679 13957
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7524 13892 7573 13920
rect 7524 13880 7530 13892
rect 7561 13889 7573 13892
rect 7607 13920 7619 13923
rect 8294 13920 8300 13932
rect 7607 13892 8300 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 3510 13852 3516 13864
rect 3292 13824 3516 13852
rect 3292 13812 3298 13824
rect 3510 13812 3516 13824
rect 3568 13852 3574 13864
rect 3605 13855 3663 13861
rect 3605 13852 3617 13855
rect 3568 13824 3617 13852
rect 3568 13812 3574 13824
rect 3605 13821 3617 13824
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 4663 13824 5089 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5077 13821 5089 13824
rect 5123 13852 5135 13855
rect 5166 13852 5172 13864
rect 5123 13824 5172 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5166 13812 5172 13824
rect 5224 13852 5230 13864
rect 5224 13824 5856 13852
rect 5224 13812 5230 13824
rect 2682 13744 2688 13796
rect 2740 13784 2746 13796
rect 3050 13784 3056 13796
rect 2740 13756 3056 13784
rect 2740 13744 2746 13756
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 3145 13787 3203 13793
rect 3145 13753 3157 13787
rect 3191 13784 3203 13787
rect 3786 13784 3792 13796
rect 3191 13756 3792 13784
rect 3191 13753 3203 13756
rect 3145 13747 3203 13753
rect 3252 13728 3280 13756
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 5828 13793 5856 13824
rect 6178 13812 6184 13864
rect 6236 13812 6242 13864
rect 6638 13852 6644 13864
rect 6551 13824 6644 13852
rect 6638 13812 6644 13824
rect 6696 13852 6702 13864
rect 8018 13852 8024 13864
rect 6696 13824 6868 13852
rect 6696 13812 6702 13824
rect 5813 13787 5871 13793
rect 5813 13753 5825 13787
rect 5859 13784 5871 13787
rect 6086 13784 6092 13796
rect 5859 13756 6092 13784
rect 5859 13753 5871 13756
rect 5813 13747 5871 13753
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 6840 13784 6868 13824
rect 7116 13824 8024 13852
rect 6914 13784 6920 13796
rect 6840 13756 6920 13784
rect 6914 13744 6920 13756
rect 6972 13744 6978 13796
rect 7116 13728 7144 13824
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8536 13824 8677 13852
rect 8536 13812 8542 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 9858 13852 9864 13864
rect 9819 13824 9864 13852
rect 8665 13815 8723 13821
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10128 13787 10186 13793
rect 10128 13753 10140 13787
rect 10174 13784 10186 13787
rect 10318 13784 10324 13796
rect 10174 13756 10324 13784
rect 10174 13753 10186 13756
rect 10128 13747 10186 13753
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 2774 13716 2780 13728
rect 2735 13688 2780 13716
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 3234 13676 3240 13728
rect 3292 13676 3298 13728
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5721 13719 5779 13725
rect 5721 13716 5733 13719
rect 5408 13688 5733 13716
rect 5408 13676 5414 13688
rect 5721 13685 5733 13688
rect 5767 13685 5779 13719
rect 5721 13679 5779 13685
rect 7098 13676 7104 13728
rect 7156 13676 7162 13728
rect 7374 13676 7380 13728
rect 7432 13716 7438 13728
rect 7469 13719 7527 13725
rect 7469 13716 7481 13719
rect 7432 13688 7481 13716
rect 7432 13676 7438 13688
rect 7469 13685 7481 13688
rect 7515 13685 7527 13719
rect 7469 13679 7527 13685
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4798 13512 4804 13524
rect 4663 13484 4804 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 4982 13512 4988 13524
rect 4943 13484 4988 13512
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7929 13515 7987 13521
rect 7929 13512 7941 13515
rect 6972 13484 7941 13512
rect 6972 13472 6978 13484
rect 7929 13481 7941 13484
rect 7975 13481 7987 13515
rect 10318 13512 10324 13524
rect 10279 13484 10324 13512
rect 7929 13475 7987 13481
rect 10318 13472 10324 13484
rect 10376 13512 10382 13524
rect 10597 13515 10655 13521
rect 10597 13512 10609 13515
rect 10376 13484 10609 13512
rect 10376 13472 10382 13484
rect 10597 13481 10609 13484
rect 10643 13481 10655 13515
rect 10597 13475 10655 13481
rect 2222 13404 2228 13456
rect 2280 13444 2286 13456
rect 2682 13444 2688 13456
rect 2280 13416 2688 13444
rect 2280 13404 2286 13416
rect 2682 13404 2688 13416
rect 2740 13444 2746 13456
rect 2869 13447 2927 13453
rect 2869 13444 2881 13447
rect 2740 13416 2881 13444
rect 2740 13404 2746 13416
rect 2869 13413 2881 13416
rect 2915 13413 2927 13447
rect 2869 13407 2927 13413
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 5690 13447 5748 13453
rect 5690 13444 5702 13447
rect 5592 13416 5702 13444
rect 5592 13404 5598 13416
rect 5690 13413 5702 13416
rect 5736 13413 5748 13447
rect 5690 13407 5748 13413
rect 5902 13404 5908 13456
rect 5960 13404 5966 13456
rect 11324 13447 11382 13453
rect 11324 13413 11336 13447
rect 11370 13444 11382 13447
rect 11514 13444 11520 13456
rect 11370 13416 11520 13444
rect 11370 13413 11382 13416
rect 11324 13407 11382 13413
rect 11514 13404 11520 13416
rect 11572 13444 11578 13456
rect 12342 13444 12348 13456
rect 11572 13416 12348 13444
rect 11572 13404 11578 13416
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 5445 13379 5503 13385
rect 3007 13348 3188 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3050 13308 3056 13320
rect 2915 13280 3056 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 2225 13243 2283 13249
rect 2225 13209 2237 13243
rect 2271 13240 2283 13243
rect 2682 13240 2688 13252
rect 2271 13212 2688 13240
rect 2271 13209 2283 13212
rect 2225 13203 2283 13209
rect 2682 13200 2688 13212
rect 2740 13240 2746 13252
rect 3160 13240 3188 13348
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 5920 13376 5948 13404
rect 5491 13348 5948 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 11054 13308 11060 13320
rect 11015 13280 11060 13308
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 3329 13243 3387 13249
rect 3329 13240 3341 13243
rect 2740 13212 3341 13240
rect 2740 13200 2746 13212
rect 3329 13209 3341 13212
rect 3375 13209 3387 13243
rect 3329 13203 3387 13209
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 2038 13172 2044 13184
rect 1719 13144 2044 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 2038 13132 2044 13144
rect 2096 13172 2102 13184
rect 2409 13175 2467 13181
rect 2409 13172 2421 13175
rect 2096 13144 2421 13172
rect 2096 13132 2102 13144
rect 2409 13141 2421 13144
rect 2455 13141 2467 13175
rect 5350 13172 5356 13184
rect 5311 13144 5356 13172
rect 2409 13135 2467 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 6825 13175 6883 13181
rect 6825 13172 6837 13175
rect 6144 13144 6837 13172
rect 6144 13132 6150 13144
rect 6825 13141 6837 13144
rect 6871 13141 6883 13175
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 6825 13135 6883 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12492 13144 12537 13172
rect 12492 13132 12498 13144
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 6917 12971 6975 12977
rect 6917 12968 6929 12971
rect 5408 12940 6929 12968
rect 5408 12928 5414 12940
rect 6917 12937 6929 12940
rect 6963 12937 6975 12971
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 6917 12931 6975 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10318 12968 10324 12980
rect 9999 12940 10324 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 2961 12903 3019 12909
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 3050 12900 3056 12912
rect 3007 12872 3056 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 3050 12860 3056 12872
rect 3108 12860 3114 12912
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 5813 12903 5871 12909
rect 5813 12900 5825 12903
rect 5592 12872 5825 12900
rect 5592 12860 5598 12872
rect 5813 12869 5825 12872
rect 5859 12869 5871 12903
rect 5813 12863 5871 12869
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 5828 12832 5856 12863
rect 5994 12860 6000 12912
rect 6052 12900 6058 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 6052 12872 6561 12900
rect 6052 12860 6058 12872
rect 6549 12869 6561 12872
rect 6595 12900 6607 12903
rect 6595 12872 7328 12900
rect 6595 12869 6607 12872
rect 6549 12863 6607 12869
rect 7300 12841 7328 12872
rect 6181 12835 6239 12841
rect 6181 12832 6193 12835
rect 2740 12804 3188 12832
rect 5828 12804 6193 12832
rect 2740 12792 2746 12804
rect 3050 12764 3056 12776
rect 3011 12736 3056 12764
rect 3050 12724 3056 12736
rect 3108 12724 3114 12776
rect 3160 12764 3188 12804
rect 6181 12801 6193 12804
rect 6227 12801 6239 12835
rect 6181 12795 6239 12801
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 3309 12767 3367 12773
rect 3309 12764 3321 12767
rect 3160 12736 3321 12764
rect 3309 12733 3321 12736
rect 3355 12733 3367 12767
rect 3309 12727 3367 12733
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 5500 12736 5549 12764
rect 5500 12724 5506 12736
rect 5537 12733 5549 12736
rect 5583 12764 5595 12767
rect 5902 12764 5908 12776
rect 5583 12736 5908 12764
rect 5583 12733 5595 12736
rect 5537 12727 5595 12733
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6196 12764 6224 12795
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 6196 12736 7481 12764
rect 7469 12733 7481 12736
rect 7515 12733 7527 12767
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 7469 12727 7527 12733
rect 8220 12736 8585 12764
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 2130 12696 2136 12708
rect 2043 12668 2136 12696
rect 2130 12656 2136 12668
rect 2188 12696 2194 12708
rect 3142 12696 3148 12708
rect 2188 12668 3148 12696
rect 2188 12656 2194 12668
rect 3142 12656 3148 12668
rect 3200 12696 3206 12708
rect 3200 12668 4476 12696
rect 3200 12656 3206 12668
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 2222 12588 2228 12640
rect 2280 12628 2286 12640
rect 4448 12637 4476 12668
rect 8220 12640 8248 12736
rect 8573 12733 8585 12736
rect 8619 12764 8631 12767
rect 9858 12764 9864 12776
rect 8619 12736 9864 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9858 12724 9864 12736
rect 9916 12764 9922 12776
rect 11054 12764 11060 12776
rect 9916 12736 11060 12764
rect 9916 12724 9922 12736
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8818 12699 8876 12705
rect 8818 12696 8830 12699
rect 8352 12668 8830 12696
rect 8352 12656 8358 12668
rect 8818 12665 8830 12668
rect 8864 12665 8876 12699
rect 8818 12659 8876 12665
rect 2501 12631 2559 12637
rect 2501 12628 2513 12631
rect 2280 12600 2513 12628
rect 2280 12588 2286 12600
rect 2501 12597 2513 12600
rect 2547 12597 2559 12631
rect 2501 12591 2559 12597
rect 4433 12631 4491 12637
rect 4433 12597 4445 12631
rect 4479 12597 4491 12631
rect 4433 12591 4491 12597
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7282 12628 7288 12640
rect 7064 12600 7288 12628
rect 7064 12588 7070 12600
rect 7282 12588 7288 12600
rect 7340 12628 7346 12640
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 7340 12600 7389 12628
rect 7340 12588 7346 12600
rect 7377 12597 7389 12600
rect 7423 12597 7435 12631
rect 7377 12591 7435 12597
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 8260 12600 8401 12628
rect 8260 12588 8266 12600
rect 8389 12597 8401 12600
rect 8435 12597 8447 12631
rect 8389 12591 8447 12597
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1912 12396 1961 12424
rect 1912 12384 1918 12396
rect 1949 12393 1961 12396
rect 1995 12424 2007 12427
rect 2299 12427 2357 12433
rect 2299 12424 2311 12427
rect 1995 12396 2311 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2299 12393 2311 12396
rect 2345 12393 2357 12427
rect 2299 12387 2357 12393
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3237 12427 3295 12433
rect 3237 12424 3249 12427
rect 3108 12396 3249 12424
rect 3108 12384 3114 12396
rect 3237 12393 3249 12396
rect 3283 12424 3295 12427
rect 5442 12424 5448 12436
rect 3283 12396 5448 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8570 12424 8576 12436
rect 8352 12396 8576 12424
rect 8352 12384 8358 12396
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 1673 12359 1731 12365
rect 1673 12325 1685 12359
rect 1719 12356 1731 12359
rect 2130 12356 2136 12368
rect 1719 12328 2136 12356
rect 1719 12325 1731 12328
rect 1673 12319 1731 12325
rect 2130 12316 2136 12328
rect 2188 12316 2194 12368
rect 2406 12316 2412 12368
rect 2464 12356 2470 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2464 12328 2789 12356
rect 2464 12316 2470 12328
rect 2777 12325 2789 12328
rect 2823 12356 2835 12359
rect 2823 12328 3004 12356
rect 2823 12325 2835 12328
rect 2777 12319 2835 12325
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2866 12220 2872 12232
rect 2827 12192 2872 12220
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 2976 12152 3004 12328
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 4982 12356 4988 12368
rect 4672 12328 4988 12356
rect 4672 12316 4678 12328
rect 4982 12316 4988 12328
rect 5040 12316 5046 12368
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 7837 12359 7895 12365
rect 7837 12356 7849 12359
rect 7524 12328 7849 12356
rect 7524 12316 7530 12328
rect 7837 12325 7849 12328
rect 7883 12325 7895 12359
rect 7837 12319 7895 12325
rect 10042 12316 10048 12368
rect 10100 12356 10106 12368
rect 10321 12359 10379 12365
rect 10321 12356 10333 12359
rect 10100 12328 10333 12356
rect 10100 12316 10106 12328
rect 10321 12325 10333 12328
rect 10367 12325 10379 12359
rect 10321 12319 10379 12325
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5258 12288 5264 12300
rect 4847 12260 5264 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 4816 12220 4844 12251
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 7650 12288 7656 12300
rect 7611 12260 7656 12288
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10413 12291 10471 12297
rect 10413 12288 10425 12291
rect 10008 12260 10425 12288
rect 10008 12248 10014 12260
rect 10413 12257 10425 12260
rect 10459 12288 10471 12291
rect 10459 12260 11652 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 4672 12192 4844 12220
rect 4672 12180 4678 12192
rect 4890 12180 4896 12232
rect 4948 12220 4954 12232
rect 5077 12223 5135 12229
rect 5077 12220 5089 12223
rect 4948 12192 5089 12220
rect 4948 12180 4954 12192
rect 5077 12189 5089 12192
rect 5123 12189 5135 12223
rect 7926 12220 7932 12232
rect 7887 12192 7932 12220
rect 5077 12183 5135 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 10226 12220 10232 12232
rect 9456 12192 10232 12220
rect 9456 12180 9462 12192
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10652 12192 10793 12220
rect 10652 12180 10658 12192
rect 10781 12189 10793 12192
rect 10827 12220 10839 12223
rect 11514 12220 11520 12232
rect 10827 12192 11520 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 11624 12220 11652 12260
rect 12618 12220 12624 12232
rect 11624 12192 12624 12220
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 7374 12152 7380 12164
rect 2832 12124 3004 12152
rect 7335 12124 7380 12152
rect 2832 12112 2838 12124
rect 7374 12112 7380 12124
rect 7432 12112 7438 12164
rect 11149 12155 11207 12161
rect 11149 12152 11161 12155
rect 10704 12124 11161 12152
rect 10704 12096 10732 12124
rect 11149 12121 11161 12124
rect 11195 12121 11207 12155
rect 11149 12115 11207 12121
rect 4522 12084 4528 12096
rect 4483 12056 4528 12084
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 9861 12087 9919 12093
rect 9861 12053 9873 12087
rect 9907 12084 9919 12087
rect 10686 12084 10692 12096
rect 9907 12056 10692 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 2682 11880 2688 11892
rect 2643 11852 2688 11880
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 2924 11852 4353 11880
rect 2924 11840 2930 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4890 11880 4896 11892
rect 4851 11852 4896 11880
rect 4341 11843 4399 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 5040 11852 5273 11880
rect 5040 11840 5046 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 7650 11880 7656 11892
rect 6319 11852 7656 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 7745 11883 7803 11889
rect 7745 11849 7757 11883
rect 7791 11880 7803 11883
rect 8202 11880 8208 11892
rect 7791 11852 8208 11880
rect 7791 11849 7803 11852
rect 7745 11843 7803 11849
rect 7852 11756 7880 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 8628 11852 9229 11880
rect 8628 11840 8634 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 10413 11815 10471 11821
rect 10413 11781 10425 11815
rect 10459 11812 10471 11815
rect 11054 11812 11060 11824
rect 10459 11784 11060 11812
rect 10459 11781 10471 11784
rect 10413 11775 10471 11781
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 7834 11744 7840 11756
rect 7747 11716 7840 11744
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10134 11744 10140 11756
rect 9732 11716 10140 11744
rect 9732 11704 9738 11716
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3050 11676 3056 11688
rect 3007 11648 3056 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 10686 11676 10692 11688
rect 10647 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 3228 11611 3286 11617
rect 3228 11577 3240 11611
rect 3274 11608 3286 11611
rect 3326 11608 3332 11620
rect 3274 11580 3332 11608
rect 3274 11577 3286 11580
rect 3228 11571 3286 11577
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 7377 11611 7435 11617
rect 7377 11577 7389 11611
rect 7423 11608 7435 11611
rect 7926 11608 7932 11620
rect 7423 11580 7932 11608
rect 7423 11577 7435 11580
rect 7377 11571 7435 11577
rect 7926 11568 7932 11580
rect 7984 11608 7990 11620
rect 8082 11611 8140 11617
rect 8082 11608 8094 11611
rect 7984 11580 8094 11608
rect 7984 11568 7990 11580
rect 8082 11577 8094 11580
rect 8128 11577 8140 11611
rect 8082 11571 8140 11577
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9732 11580 10149 11608
rect 9732 11568 9738 11580
rect 10137 11577 10149 11580
rect 10183 11608 10195 11611
rect 10226 11608 10232 11620
rect 10183 11580 10232 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 10594 11568 10600 11620
rect 10652 11608 10658 11620
rect 10965 11611 11023 11617
rect 10965 11608 10977 11611
rect 10652 11580 10977 11608
rect 10652 11568 10658 11580
rect 10965 11577 10977 11580
rect 11011 11577 11023 11611
rect 10965 11571 11023 11577
rect 2317 11543 2375 11549
rect 2317 11509 2329 11543
rect 2363 11540 2375 11543
rect 2774 11540 2780 11552
rect 2363 11512 2780 11540
rect 2363 11509 2375 11512
rect 2317 11503 2375 11509
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 6641 11543 6699 11549
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 7466 11540 7472 11552
rect 6687 11512 7472 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10042 11540 10048 11552
rect 9907 11512 10048 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10870 11540 10876 11552
rect 10831 11512 10876 11540
rect 10870 11500 10876 11512
rect 10928 11540 10934 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 10928 11512 11345 11540
rect 10928 11500 10934 11512
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11333 11503 11391 11509
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12802 11540 12808 11552
rect 12483 11512 12808 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 1452 11308 1593 11336
rect 1452 11296 1458 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 1581 11299 1639 11305
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2866 11336 2872 11348
rect 2363 11308 2872 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3050 11336 3056 11348
rect 3011 11308 3056 11336
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 4525 11339 4583 11345
rect 4525 11305 4537 11339
rect 4571 11336 4583 11339
rect 4614 11336 4620 11348
rect 4571 11308 4620 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 6638 11336 6644 11348
rect 4948 11308 6644 11336
rect 4948 11296 4954 11308
rect 6638 11296 6644 11308
rect 6696 11336 6702 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6696 11308 6837 11336
rect 6696 11296 6702 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7616 11308 7665 11336
rect 7616 11296 7622 11308
rect 7653 11305 7665 11308
rect 7699 11336 7711 11339
rect 7834 11336 7840 11348
rect 7699 11308 7840 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8481 11339 8539 11345
rect 8481 11336 8493 11339
rect 8444 11308 8493 11336
rect 8444 11296 8450 11308
rect 8481 11305 8493 11308
rect 8527 11305 8539 11339
rect 9950 11336 9956 11348
rect 9911 11308 9956 11336
rect 8481 11299 8539 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 13078 11336 13084 11348
rect 12176 11308 13084 11336
rect 5712 11271 5770 11277
rect 5712 11237 5724 11271
rect 5758 11268 5770 11271
rect 6086 11268 6092 11280
rect 5758 11240 6092 11268
rect 5758 11237 5770 11240
rect 5712 11231 5770 11237
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 10962 11268 10968 11280
rect 10923 11240 10968 11268
rect 10962 11228 10968 11240
rect 11020 11268 11026 11280
rect 12051 11271 12109 11277
rect 12051 11268 12063 11271
rect 11020 11240 12063 11268
rect 11020 11228 11026 11240
rect 12051 11237 12063 11240
rect 12097 11237 12109 11271
rect 12051 11231 12109 11237
rect 5442 11200 5448 11212
rect 5403 11172 5448 11200
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10594 11200 10600 11212
rect 10192 11172 10600 11200
rect 10192 11160 10198 11172
rect 10594 11160 10600 11172
rect 10652 11200 10658 11212
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10652 11172 11069 11200
rect 10652 11160 10658 11172
rect 11057 11169 11069 11172
rect 11103 11200 11115 11203
rect 12176 11200 12204 11308
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 12529 11271 12587 11277
rect 12529 11268 12541 11271
rect 12400 11240 12541 11268
rect 12400 11228 12406 11240
rect 12529 11237 12541 11240
rect 12575 11237 12587 11271
rect 12529 11231 12587 11237
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 12676 11240 12721 11268
rect 12676 11228 12682 11240
rect 12710 11200 12716 11212
rect 11103 11172 12204 11200
rect 12544 11172 12716 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 3326 11064 3332 11076
rect 3287 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 7650 11024 7656 11076
rect 7708 11064 7714 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 7708 11036 8033 11064
rect 7708 11024 7714 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8404 11064 8432 11095
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8536 11104 8585 11132
rect 8536 11092 8542 11104
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 12544 11141 12572 11172
rect 12710 11160 12716 11172
rect 12768 11200 12774 11212
rect 12894 11200 12900 11212
rect 12768 11172 12900 11200
rect 12768 11160 12774 11172
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10376 11104 10885 11132
rect 10376 11092 10382 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 8021 11027 8079 11033
rect 8220 11036 8432 11064
rect 10505 11067 10563 11073
rect 7374 10956 7380 11008
rect 7432 10996 7438 11008
rect 8220 10996 8248 11036
rect 10505 11033 10517 11067
rect 10551 11064 10563 11067
rect 11885 11067 11943 11073
rect 10551 11036 11284 11064
rect 10551 11033 10563 11036
rect 10505 11027 10563 11033
rect 11256 11008 11284 11036
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 12636 11064 12664 11092
rect 11931 11036 12664 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 7432 10968 8248 10996
rect 7432 10956 7438 10968
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 11425 10999 11483 11005
rect 11425 10996 11437 10999
rect 11296 10968 11437 10996
rect 11296 10956 11302 10968
rect 11425 10965 11437 10968
rect 11471 10965 11483 10999
rect 13078 10996 13084 11008
rect 13039 10968 13084 10996
rect 11425 10959 11483 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6086 10792 6092 10804
rect 6047 10764 6092 10792
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8536 10764 8953 10792
rect 8536 10752 8542 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10962 10792 10968 10804
rect 9815 10764 10968 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12342 10792 12348 10804
rect 12115 10764 12348 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 10134 10724 10140 10736
rect 10095 10696 10140 10724
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10318 10684 10324 10736
rect 10376 10724 10382 10736
rect 10413 10727 10471 10733
rect 10413 10724 10425 10727
rect 10376 10696 10425 10724
rect 10376 10684 10382 10696
rect 10413 10693 10425 10696
rect 10459 10693 10471 10727
rect 10413 10687 10471 10693
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 11146 10724 11152 10736
rect 10827 10696 11152 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10724 12587 10727
rect 13354 10724 13360 10736
rect 12575 10696 13360 10724
rect 12575 10693 12587 10696
rect 12529 10687 12587 10693
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 7558 10656 7564 10668
rect 7519 10628 7564 10656
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 11238 10656 11244 10668
rect 11199 10628 11244 10656
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 12434 10656 12440 10668
rect 11388 10628 12440 10656
rect 11388 10616 11394 10628
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4522 10588 4528 10600
rect 4304 10560 4528 10588
rect 4304 10548 4310 10560
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10588 12866 10600
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 12860 10560 13461 10588
rect 12860 10548 12866 10560
rect 13449 10557 13461 10560
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 7101 10523 7159 10529
rect 7101 10489 7113 10523
rect 7147 10520 7159 10523
rect 7828 10523 7886 10529
rect 7828 10520 7840 10523
rect 7147 10492 7840 10520
rect 7147 10489 7159 10492
rect 7101 10483 7159 10489
rect 7828 10489 7840 10492
rect 7874 10520 7886 10523
rect 8110 10520 8116 10532
rect 7874 10492 8116 10520
rect 7874 10489 7886 10492
rect 7828 10483 7886 10489
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 11054 10480 11060 10532
rect 11112 10520 11118 10532
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 11112 10492 11253 10520
rect 11112 10480 11118 10492
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11241 10483 11299 10489
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 4982 10452 4988 10464
rect 4571 10424 4988 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 6914 10452 6920 10464
rect 5675 10424 6920 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12768 10424 13001 10452
rect 12768 10412 12774 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1762 10248 1768 10260
rect 1719 10220 1768 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 8386 10248 8392 10260
rect 8347 10220 8392 10248
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8536 10220 8677 10248
rect 8536 10208 8542 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 8665 10211 8723 10217
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 9824 10220 10425 10248
rect 9824 10208 9830 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 10965 10251 11023 10257
rect 10965 10217 10977 10251
rect 11011 10248 11023 10251
rect 11330 10248 11336 10260
rect 11011 10220 11336 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 6638 10189 6644 10192
rect 4617 10183 4675 10189
rect 4617 10180 4629 10183
rect 4304 10152 4629 10180
rect 4304 10140 4310 10152
rect 4617 10149 4629 10152
rect 4663 10149 4675 10183
rect 6632 10180 6644 10189
rect 6599 10152 6644 10180
rect 4617 10143 4675 10149
rect 6632 10143 6644 10152
rect 6638 10140 6644 10143
rect 6696 10140 6702 10192
rect 11054 10140 11060 10192
rect 11112 10180 11118 10192
rect 11241 10183 11299 10189
rect 11241 10180 11253 10183
rect 11112 10152 11253 10180
rect 11112 10140 11118 10152
rect 11241 10149 11253 10152
rect 11287 10149 11299 10183
rect 11241 10143 11299 10149
rect 11790 10140 11796 10192
rect 11848 10180 11854 10192
rect 11977 10183 12035 10189
rect 11977 10180 11989 10183
rect 11848 10152 11989 10180
rect 11848 10140 11854 10152
rect 11977 10149 11989 10152
rect 12023 10149 12035 10183
rect 11977 10143 12035 10149
rect 12069 10183 12127 10189
rect 12069 10149 12081 10183
rect 12115 10180 12127 10183
rect 12158 10180 12164 10192
rect 12115 10152 12164 10180
rect 12115 10149 12127 10152
rect 12069 10143 12127 10149
rect 12158 10140 12164 10152
rect 12216 10180 12222 10192
rect 13078 10180 13084 10192
rect 12216 10152 13084 10180
rect 12216 10140 12222 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 13354 10180 13360 10192
rect 13315 10152 13360 10180
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 13538 10180 13544 10192
rect 13499 10152 13544 10180
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4396 10084 4445 10112
rect 4396 10072 4402 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 6362 10112 6368 10124
rect 5592 10084 6368 10112
rect 5592 10072 5598 10084
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10008 10084 10517 10112
rect 10008 10072 10014 10084
rect 10505 10081 10517 10084
rect 10551 10112 10563 10115
rect 10594 10112 10600 10124
rect 10551 10084 10600 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 12492 10084 13645 10112
rect 12492 10072 12498 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 10284 10016 10333 10044
rect 10284 10004 10290 10016
rect 10321 10013 10333 10016
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 11388 10016 11897 10044
rect 11388 10004 11394 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 4062 9976 4068 9988
rect 3927 9948 4068 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10870 9976 10876 9988
rect 9999 9948 10876 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10870 9936 10876 9948
rect 10928 9936 10934 9988
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 13081 9979 13139 9985
rect 13081 9976 13093 9979
rect 12584 9948 13093 9976
rect 12584 9936 12590 9948
rect 13081 9945 13093 9948
rect 13127 9945 13139 9979
rect 13081 9939 13139 9945
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3142 9908 3148 9920
rect 3007 9880 3148 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 4154 9908 4160 9920
rect 4115 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 5166 9908 5172 9920
rect 5127 9880 5172 9908
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8110 9908 8116 9920
rect 7791 9880 8116 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 11514 9908 11520 9920
rect 11475 9880 11520 9908
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12710 9908 12716 9920
rect 12483 9880 12716 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 12860 9880 12905 9908
rect 12860 9868 12866 9880
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 6089 9707 6147 9713
rect 3292 9676 3832 9704
rect 3292 9664 3298 9676
rect 3804 9648 3832 9676
rect 6089 9673 6101 9707
rect 6135 9704 6147 9707
rect 6638 9704 6644 9716
rect 6135 9676 6644 9704
rect 6135 9673 6147 9676
rect 6089 9667 6147 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 8478 9704 8484 9716
rect 8439 9676 8484 9704
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 9861 9707 9919 9713
rect 9861 9704 9873 9707
rect 9824 9676 9873 9704
rect 9824 9664 9830 9676
rect 9861 9673 9873 9676
rect 9907 9673 9919 9707
rect 10226 9704 10232 9716
rect 10187 9676 10232 9704
rect 9861 9667 9919 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10594 9704 10600 9716
rect 10555 9676 10600 9704
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 11425 9707 11483 9713
rect 11425 9704 11437 9707
rect 11388 9676 11437 9704
rect 11388 9664 11394 9676
rect 11425 9673 11437 9676
rect 11471 9673 11483 9707
rect 11425 9667 11483 9673
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 12713 9707 12771 9713
rect 12713 9704 12725 9707
rect 11572 9676 12725 9704
rect 11572 9664 11578 9676
rect 12713 9673 12725 9676
rect 12759 9704 12771 9707
rect 13538 9704 13544 9716
rect 12759 9676 13544 9704
rect 12759 9673 12771 9676
rect 12713 9667 12771 9673
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3786 9596 3792 9648
rect 3844 9596 3850 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 3988 9608 4537 9636
rect 3988 9580 4016 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 6362 9636 6368 9648
rect 6323 9608 6368 9636
rect 4525 9599 4583 9605
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 7466 9636 7472 9648
rect 7427 9608 7472 9636
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 3510 9568 3516 9580
rect 2976 9540 3516 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1762 9500 1768 9512
rect 1443 9472 1768 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 2976 9500 3004 9540
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3970 9528 3976 9580
rect 4028 9528 4034 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4120 9540 4997 9568
rect 4120 9528 4126 9540
rect 4985 9537 4997 9540
rect 5031 9568 5043 9571
rect 5074 9568 5080 9580
rect 5031 9540 5080 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8496 9568 8524 9664
rect 11790 9636 11796 9648
rect 11751 9608 11796 9636
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12158 9636 12164 9648
rect 12119 9608 12164 9636
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 12250 9596 12256 9648
rect 12308 9636 12314 9648
rect 12434 9636 12440 9648
rect 12308 9608 12440 9636
rect 12308 9596 12314 9608
rect 12434 9596 12440 9608
rect 12492 9636 12498 9648
rect 12989 9639 13047 9645
rect 12989 9636 13001 9639
rect 12492 9608 13001 9636
rect 12492 9596 12498 9608
rect 12989 9605 13001 9608
rect 13035 9605 13047 9639
rect 12989 9599 13047 9605
rect 8067 9540 8524 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 2455 9472 3004 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 3108 9472 5120 9500
rect 3108 9460 3114 9472
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 2866 9432 2872 9444
rect 2823 9404 2872 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 2866 9392 2872 9404
rect 2924 9432 2930 9444
rect 3234 9432 3240 9444
rect 2924 9404 3240 9432
rect 2924 9392 2930 9404
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 4982 9432 4988 9444
rect 4943 9404 4988 9432
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 5092 9441 5120 9472
rect 7944 9472 8769 9500
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5166 9432 5172 9444
rect 5123 9404 5172 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 7745 9435 7803 9441
rect 7745 9401 7757 9435
rect 7791 9401 7803 9435
rect 7745 9395 7803 9401
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 3050 9364 3056 9376
rect 2096 9336 3056 9364
rect 2096 9324 2102 9336
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 3200 9336 3433 9364
rect 3200 9324 3206 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 3421 9327 3479 9333
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4338 9364 4344 9376
rect 4203 9336 4344 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 4764 9336 5457 9364
rect 4764 9324 4770 9336
rect 5445 9333 5457 9336
rect 5491 9364 5503 9367
rect 5810 9364 5816 9376
rect 5491 9336 5816 9364
rect 5491 9333 5503 9336
rect 5445 9327 5503 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9364 7254 9376
rect 7760 9364 7788 9395
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 7944 9441 7972 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 13357 9503 13415 9509
rect 13357 9500 13369 9503
rect 10192 9472 13369 9500
rect 10192 9460 10198 9472
rect 13357 9469 13369 9472
rect 13403 9500 13415 9503
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13403 9472 13921 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 7929 9435 7987 9441
rect 7929 9432 7941 9435
rect 7892 9404 7941 9432
rect 7892 9392 7898 9404
rect 7929 9401 7941 9404
rect 7975 9401 7987 9435
rect 7929 9395 7987 9401
rect 13538 9364 13544 9376
rect 7248 9336 7788 9364
rect 13499 9336 13544 9364
rect 7248 9324 7254 9336
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2832 9132 2973 9160
rect 2832 9120 2838 9132
rect 2961 9129 2973 9132
rect 3007 9160 3019 9163
rect 4062 9160 4068 9172
rect 3007 9132 4068 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5224 9132 5641 9160
rect 5224 9120 5230 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 6914 9160 6920 9172
rect 6875 9132 6920 9160
rect 5629 9123 5687 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11204 9132 11897 9160
rect 11204 9120 11210 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 13504 9132 13645 9160
rect 13504 9120 13510 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 1673 9095 1731 9101
rect 1673 9061 1685 9095
rect 1719 9092 1731 9095
rect 3050 9092 3056 9104
rect 1719 9064 2912 9092
rect 3011 9064 3056 9092
rect 1719 9061 1731 9064
rect 1673 9055 1731 9061
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 2774 9024 2780 9036
rect 2648 8996 2780 9024
rect 2648 8984 2654 8996
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 2884 9024 2912 9064
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 4494 9095 4552 9101
rect 4494 9092 4506 9095
rect 3568 9064 4506 9092
rect 3568 9052 3574 9064
rect 4494 9061 4506 9064
rect 4540 9092 4552 9095
rect 4706 9092 4712 9104
rect 4540 9064 4712 9092
rect 4540 9061 4552 9064
rect 4494 9055 4552 9061
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 7926 9052 7932 9104
rect 7984 9092 7990 9104
rect 8021 9095 8079 9101
rect 8021 9092 8033 9095
rect 7984 9064 8033 9092
rect 7984 9052 7990 9064
rect 8021 9061 8033 9064
rect 8067 9061 8079 9095
rect 8021 9055 8079 9061
rect 10229 9095 10287 9101
rect 10229 9061 10241 9095
rect 10275 9092 10287 9095
rect 10594 9092 10600 9104
rect 10275 9064 10600 9092
rect 10275 9061 10287 9064
rect 10229 9055 10287 9061
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 11977 9095 12035 9101
rect 11977 9061 11989 9095
rect 12023 9092 12035 9095
rect 12342 9092 12348 9104
rect 12023 9064 12348 9092
rect 12023 9061 12035 9064
rect 11977 9055 12035 9061
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 13170 9092 13176 9104
rect 13131 9064 13176 9092
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 3881 9027 3939 9033
rect 2884 8996 3004 9024
rect 2976 8968 3004 8996
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4062 9024 4068 9036
rect 3927 8996 4068 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4338 9024 4344 9036
rect 4295 8996 4344 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 5534 9024 5540 9036
rect 4396 8996 5540 9024
rect 4396 8984 4402 8996
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9916 8996 10057 9024
rect 9916 8984 9922 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11480 8996 11713 9024
rect 11480 8984 11486 8996
rect 11701 8993 11713 8996
rect 11747 9024 11759 9027
rect 12250 9024 12256 9036
rect 11747 8996 12256 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12894 9033 12900 9036
rect 12886 9027 12900 9033
rect 12886 9024 12898 9027
rect 12452 8996 12898 9024
rect 2958 8956 2964 8968
rect 2919 8928 2964 8956
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 8110 8956 8116 8968
rect 8071 8928 8116 8956
rect 7929 8919 7987 8925
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 3142 8888 3148 8900
rect 2740 8860 3148 8888
rect 2740 8848 2746 8860
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3602 8848 3608 8900
rect 3660 8888 3666 8900
rect 4062 8888 4068 8900
rect 3660 8860 4068 8888
rect 3660 8848 3666 8860
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 7561 8891 7619 8897
rect 7561 8857 7573 8891
rect 7607 8888 7619 8891
rect 7834 8888 7840 8900
rect 7607 8860 7840 8888
rect 7607 8857 7619 8860
rect 7561 8851 7619 8857
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 7944 8888 7972 8919
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 12452 8956 12480 8996
rect 12886 8993 12898 8996
rect 12886 8987 12900 8993
rect 12894 8984 12900 8987
rect 12952 8984 12958 9036
rect 11440 8928 12480 8956
rect 8202 8888 8208 8900
rect 7944 8860 8208 8888
rect 8202 8848 8208 8860
rect 8260 8888 8266 8900
rect 11440 8897 11468 8928
rect 8849 8891 8907 8897
rect 8849 8888 8861 8891
rect 8260 8860 8861 8888
rect 8260 8848 8266 8860
rect 8849 8857 8861 8860
rect 8895 8857 8907 8891
rect 8849 8851 8907 8857
rect 11425 8891 11483 8897
rect 11425 8857 11437 8891
rect 11471 8857 11483 8891
rect 11425 8851 11483 8857
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8820 2559 8823
rect 2774 8820 2780 8832
rect 2547 8792 2780 8820
rect 2547 8789 2559 8792
rect 2501 8783 2559 8789
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 9766 8820 9772 8832
rect 9727 8792 9772 8820
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3568 8588 3893 8616
rect 3568 8576 3574 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 5040 8588 5273 8616
rect 5040 8576 5046 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 6917 8619 6975 8625
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 7006 8616 7012 8628
rect 6963 8588 7012 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8202 8616 8208 8628
rect 8163 8588 8208 8616
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 12894 8616 12900 8628
rect 12855 8588 12900 8616
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 5077 8551 5135 8557
rect 5077 8517 5089 8551
rect 5123 8548 5135 8551
rect 5994 8548 6000 8560
rect 5123 8520 6000 8548
rect 5123 8517 5135 8520
rect 5077 8511 5135 8517
rect 5644 8489 5672 8520
rect 5994 8508 6000 8520
rect 6052 8548 6058 8560
rect 6270 8548 6276 8560
rect 6052 8520 6276 8548
rect 6052 8508 6058 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 8846 8508 8852 8560
rect 8904 8548 8910 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 8904 8520 8953 8548
rect 8904 8508 8910 8520
rect 8941 8517 8953 8520
rect 8987 8517 8999 8551
rect 8941 8511 8999 8517
rect 11425 8551 11483 8557
rect 11425 8517 11437 8551
rect 11471 8548 11483 8551
rect 11514 8548 11520 8560
rect 11471 8520 11520 8548
rect 11471 8517 11483 8520
rect 11425 8511 11483 8517
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5629 8443 5687 8449
rect 5810 8440 5816 8452
rect 5868 8480 5874 8492
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5868 8452 6193 8480
rect 5868 8440 5874 8452
rect 6181 8449 6193 8452
rect 6227 8480 6239 8483
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 6227 8452 7481 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7834 8480 7840 8492
rect 7795 8452 7840 8480
rect 7469 8443 7527 8449
rect 7834 8440 7840 8452
rect 7892 8480 7898 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 7892 8452 8677 8480
rect 7892 8440 7898 8452
rect 8665 8449 8677 8452
rect 8711 8480 8723 8483
rect 8711 8452 9444 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 1964 8288 1992 8375
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2205 8415 2263 8421
rect 2205 8412 2217 8415
rect 2096 8384 2217 8412
rect 2096 8372 2102 8384
rect 2205 8381 2217 8384
rect 2251 8381 2263 8415
rect 2205 8375 2263 8381
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 6972 8384 7205 8412
rect 6972 8372 6978 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 8260 8384 9229 8412
rect 8260 8372 8266 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 6362 8304 6368 8356
rect 6420 8344 6426 8356
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 6420 8316 6653 8344
rect 6420 8304 6426 8316
rect 6641 8313 6653 8316
rect 6687 8344 6699 8347
rect 7374 8344 7380 8356
rect 6687 8316 7380 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 9416 8353 9444 8452
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8412 11299 8415
rect 11606 8412 11612 8424
rect 11287 8384 11612 8412
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 11606 8372 11612 8384
rect 11664 8412 11670 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11664 8384 11805 8412
rect 11664 8372 11670 8384
rect 11793 8381 11805 8384
rect 11839 8412 11851 8415
rect 11974 8412 11980 8424
rect 11839 8384 11980 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 13078 8412 13084 8424
rect 13039 8384 13084 8412
rect 13078 8372 13084 8384
rect 13136 8412 13142 8424
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 13136 8384 13645 8412
rect 13136 8372 13142 8384
rect 13633 8381 13645 8384
rect 13679 8381 13691 8415
rect 13633 8375 13691 8381
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8313 9459 8347
rect 9401 8307 9459 8313
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 9548 8316 9593 8344
rect 9548 8304 9554 8316
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 1946 8276 1952 8288
rect 1903 8248 1952 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 3326 8276 3332 8288
rect 2740 8248 3332 8276
rect 2740 8236 2746 8248
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 4338 8276 4344 8288
rect 4299 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 4709 8279 4767 8285
rect 4709 8245 4721 8279
rect 4755 8276 4767 8279
rect 5718 8276 5724 8288
rect 4755 8248 5724 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 5718 8236 5724 8248
rect 5776 8276 5782 8288
rect 6086 8276 6092 8288
rect 5776 8248 6092 8276
rect 5776 8236 5782 8248
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 10229 8279 10287 8285
rect 10229 8276 10241 8279
rect 9640 8248 10241 8276
rect 9640 8236 9646 8248
rect 10229 8245 10241 8248
rect 10275 8276 10287 8279
rect 10318 8276 10324 8288
rect 10275 8248 10324 8276
rect 10275 8245 10287 8248
rect 10229 8239 10287 8245
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 10594 8276 10600 8288
rect 10555 8248 10600 8276
rect 10594 8236 10600 8248
rect 10652 8236 10658 8288
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12342 8276 12348 8288
rect 12299 8248 12348 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 13262 8276 13268 8288
rect 13223 8248 13268 8276
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2590 8072 2596 8084
rect 1995 8044 2596 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2832 8044 2973 8072
rect 2832 8032 2838 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3970 8072 3976 8084
rect 3559 8044 3976 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 2038 7964 2044 8016
rect 2096 8004 2102 8016
rect 2225 8007 2283 8013
rect 2225 8004 2237 8007
rect 2096 7976 2237 8004
rect 2096 7964 2102 7976
rect 2225 7973 2237 7976
rect 2271 7973 2283 8007
rect 2225 7967 2283 7973
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 2884 7908 3065 7936
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 2884 7868 2912 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 2740 7840 2912 7868
rect 2961 7871 3019 7877
rect 2740 7828 2746 7840
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3528 7868 3556 8035
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 4982 8072 4988 8084
rect 4856 8044 4988 8072
rect 4856 8032 4862 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 5868 8044 6377 8072
rect 5868 8032 5874 8044
rect 6365 8041 6377 8044
rect 6411 8072 6423 8075
rect 6917 8075 6975 8081
rect 6917 8072 6929 8075
rect 6411 8044 6929 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6917 8041 6929 8044
rect 6963 8041 6975 8075
rect 6917 8035 6975 8041
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 8110 8072 8116 8084
rect 7607 8044 8116 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8680 8044 9137 8072
rect 5252 8007 5310 8013
rect 5252 7973 5264 8007
rect 5298 8004 5310 8007
rect 5442 8004 5448 8016
rect 5298 7976 5448 8004
rect 5298 7973 5310 7976
rect 5252 7967 5310 7973
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 8386 8004 8392 8016
rect 8347 7976 8392 8004
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 8570 8004 8576 8016
rect 8531 7976 8576 8004
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 8680 8013 8708 8044
rect 9125 8041 9137 8044
rect 9171 8072 9183 8075
rect 9490 8072 9496 8084
rect 9171 8044 9496 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9490 8032 9496 8044
rect 9548 8072 9554 8084
rect 11422 8072 11428 8084
rect 9548 8044 10364 8072
rect 11383 8044 11428 8072
rect 9548 8032 9554 8044
rect 8665 8007 8723 8013
rect 8665 7973 8677 8007
rect 8711 7973 8723 8007
rect 8665 7967 8723 7973
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8680 7936 8708 7967
rect 9858 7964 9864 8016
rect 9916 8004 9922 8016
rect 10336 8013 10364 8044
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 10229 8007 10287 8013
rect 10229 8004 10241 8007
rect 9916 7976 10241 8004
rect 9916 7964 9922 7976
rect 10229 7973 10241 7976
rect 10275 7973 10287 8007
rect 10229 7967 10287 7973
rect 10321 8007 10379 8013
rect 10321 7973 10333 8007
rect 10367 8004 10379 8007
rect 10502 8004 10508 8016
rect 10367 7976 10508 8004
rect 10367 7973 10379 7976
rect 10321 7967 10379 7973
rect 10502 7964 10508 7976
rect 10560 8004 10566 8016
rect 10560 7976 13216 8004
rect 10560 7964 10566 7976
rect 10042 7936 10048 7948
rect 7975 7908 8708 7936
rect 10003 7908 10048 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 12060 7939 12118 7945
rect 12060 7905 12072 7939
rect 12106 7936 12118 7939
rect 12342 7936 12348 7948
rect 12106 7908 12348 7936
rect 12106 7905 12118 7908
rect 12060 7899 12118 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 3007 7840 3556 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4396 7840 4997 7868
rect 4396 7828 4402 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 4985 7831 5043 7837
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7732 4399 7735
rect 4798 7732 4804 7744
rect 4387 7704 4804 7732
rect 4387 7701 4399 7704
rect 4341 7695 4399 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5000 7732 5028 7831
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 9769 7803 9827 7809
rect 9769 7769 9781 7803
rect 9815 7800 9827 7803
rect 10594 7800 10600 7812
rect 9815 7772 10600 7800
rect 9815 7769 9827 7772
rect 9769 7763 9827 7769
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 13188 7809 13216 7976
rect 13173 7803 13231 7809
rect 13173 7769 13185 7803
rect 13219 7769 13231 7803
rect 13173 7763 13231 7769
rect 5258 7732 5264 7744
rect 5000 7704 5264 7732
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8294 7732 8300 7744
rect 8159 7704 8300 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9582 7732 9588 7744
rect 9539 7704 9588 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 10686 7732 10692 7744
rect 10647 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2682 7528 2688 7540
rect 2547 7500 2688 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2832 7500 3157 7528
rect 2832 7488 2838 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4304 7500 4353 7528
rect 4304 7488 4310 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 8628 7500 8769 7528
rect 8628 7488 8634 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 8757 7491 8815 7497
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 9125 7463 9183 7469
rect 9125 7460 9137 7463
rect 8444 7432 9137 7460
rect 8444 7420 8450 7432
rect 9125 7429 9137 7432
rect 9171 7429 9183 7463
rect 9125 7423 9183 7429
rect 9769 7463 9827 7469
rect 9769 7429 9781 7463
rect 9815 7460 9827 7463
rect 9858 7460 9864 7472
rect 9815 7432 9864 7460
rect 9815 7429 9827 7432
rect 9769 7423 9827 7429
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 6472 7364 6960 7392
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2498 7324 2504 7336
rect 1443 7296 2504 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 3835 7296 4905 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 4893 7293 4905 7296
rect 4939 7324 4951 7327
rect 5442 7324 5448 7336
rect 4939 7296 5448 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5442 7284 5448 7296
rect 5500 7324 5506 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5500 7296 5641 7324
rect 5500 7284 5506 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 198 7216 204 7268
rect 256 7256 262 7268
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 256 7228 4077 7256
rect 256 7216 262 7228
rect 4065 7225 4077 7228
rect 4111 7256 4123 7259
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4111 7228 4813 7256
rect 4111 7225 4123 7228
rect 4065 7219 4123 7225
rect 4801 7225 4813 7228
rect 4847 7256 4859 7259
rect 6472 7256 6500 7364
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 4847 7228 6500 7256
rect 6564 7296 6837 7324
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 5258 7188 5264 7200
rect 2832 7160 2877 7188
rect 5219 7160 5264 7188
rect 2832 7148 2838 7160
rect 5258 7148 5264 7160
rect 5316 7188 5322 7200
rect 6564 7197 6592 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6932 7324 6960 7364
rect 7374 7324 7380 7336
rect 6932 7296 7380 7324
rect 6825 7287 6883 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 9858 7324 9864 7336
rect 9819 7296 9864 7324
rect 9858 7284 9864 7296
rect 9916 7324 9922 7336
rect 10686 7324 10692 7336
rect 9916 7296 10692 7324
rect 9916 7284 9922 7296
rect 10686 7284 10692 7296
rect 10744 7324 10750 7336
rect 11790 7324 11796 7336
rect 10744 7296 11796 7324
rect 10744 7284 10750 7296
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 7070 7259 7128 7265
rect 7070 7256 7082 7259
rect 6972 7228 7082 7256
rect 6972 7216 6978 7228
rect 7070 7225 7082 7228
rect 7116 7225 7128 7259
rect 7070 7219 7128 7225
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 10106 7259 10164 7265
rect 10106 7256 10118 7259
rect 9640 7228 10118 7256
rect 9640 7216 9646 7228
rect 10106 7225 10118 7228
rect 10152 7225 10164 7259
rect 10106 7219 10164 7225
rect 11422 7216 11428 7268
rect 11480 7256 11486 7268
rect 12728 7256 12756 7287
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 11480 7228 13277 7256
rect 11480 7216 11486 7228
rect 13265 7225 13277 7228
rect 13311 7225 13323 7259
rect 13265 7219 13323 7225
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 5316 7160 6561 7188
rect 5316 7148 5322 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 8202 7188 8208 7200
rect 8163 7160 8208 7188
rect 6549 7151 6607 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 10376 7160 11253 7188
rect 10376 7148 10382 7160
rect 11241 7157 11253 7160
rect 11287 7157 11299 7191
rect 11241 7151 11299 7157
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12342 7188 12348 7200
rect 12299 7160 12348 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 14182 7188 14188 7200
rect 12943 7160 14188 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 5442 6984 5448 6996
rect 5403 6956 5448 6984
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 6914 6984 6920 6996
rect 6875 6956 6920 6984
rect 6914 6944 6920 6956
rect 6972 6984 6978 6996
rect 7558 6984 7564 6996
rect 6972 6956 7564 6984
rect 6972 6944 6978 6956
rect 7558 6944 7564 6956
rect 7616 6984 7622 6996
rect 8481 6987 8539 6993
rect 8481 6984 8493 6987
rect 7616 6956 8493 6984
rect 7616 6944 7622 6956
rect 8481 6953 8493 6956
rect 8527 6953 8539 6987
rect 8481 6947 8539 6953
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10042 6984 10048 6996
rect 9999 6956 10048 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 9493 6919 9551 6925
rect 2556 6888 2912 6916
rect 2556 6876 2562 6888
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1670 6848 1676 6860
rect 1443 6820 1676 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2685 6851 2743 6857
rect 2685 6848 2697 6851
rect 1912 6820 2697 6848
rect 1912 6808 1918 6820
rect 2685 6817 2697 6820
rect 2731 6848 2743 6851
rect 2774 6848 2780 6860
rect 2731 6820 2780 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 2884 6848 2912 6888
rect 9493 6885 9505 6919
rect 9539 6916 9551 6919
rect 10502 6916 10508 6928
rect 9539 6888 10508 6916
rect 9539 6885 9551 6888
rect 9493 6879 9551 6885
rect 10502 6876 10508 6888
rect 10560 6925 10566 6928
rect 10560 6919 10624 6925
rect 10560 6885 10578 6919
rect 10612 6885 10624 6919
rect 10560 6879 10624 6885
rect 10560 6876 10566 6879
rect 4338 6857 4344 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 2884 6820 3801 6848
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 4332 6848 4344 6857
rect 4299 6820 4344 6848
rect 3789 6811 3847 6817
rect 4332 6811 4344 6820
rect 4338 6808 4344 6811
rect 4396 6808 4402 6860
rect 7368 6851 7426 6857
rect 7368 6817 7380 6851
rect 7414 6848 7426 6851
rect 7650 6848 7656 6860
rect 7414 6820 7656 6848
rect 7414 6817 7426 6820
rect 7368 6811 7426 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8352 6820 9045 6848
rect 8352 6808 8358 6820
rect 9033 6817 9045 6820
rect 9079 6848 9091 6851
rect 9306 6848 9312 6860
rect 9079 6820 9312 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 12802 6848 12808 6860
rect 12763 6820 12808 6848
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1544 6752 1593 6780
rect 1544 6740 1550 6752
rect 1581 6749 1593 6752
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 2869 6743 2927 6749
rect 2774 6672 2780 6724
rect 2832 6712 2838 6724
rect 2884 6712 2912 6743
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 7098 6780 7104 6792
rect 7059 6752 7104 6780
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10226 6780 10232 6792
rect 9916 6752 10232 6780
rect 9916 6740 9922 6752
rect 10226 6740 10232 6752
rect 10284 6780 10290 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 10284 6752 10333 6780
rect 10284 6740 10290 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 2832 6684 2912 6712
rect 2832 6672 2838 6684
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2464 6616 2513 6644
rect 2464 6604 2470 6616
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 2501 6607 2559 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11296 6616 11713 6644
rect 11296 6604 11302 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 12989 6647 13047 6653
rect 12989 6613 13001 6647
rect 13035 6644 13047 6647
rect 13722 6644 13728 6656
rect 13035 6616 13728 6644
rect 13035 6613 13047 6616
rect 12989 6607 13047 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2314 6440 2320 6452
rect 2188 6412 2320 6440
rect 2188 6400 2194 6412
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 10502 6400 10508 6452
rect 10560 6440 10566 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10560 6412 10701 6440
rect 10560 6400 10566 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 10689 6403 10747 6409
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 12618 6440 12624 6452
rect 11931 6412 12624 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 9030 6372 9036 6384
rect 8991 6344 9036 6372
rect 9030 6332 9036 6344
rect 9088 6332 9094 6384
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 8895 6276 9628 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9600 6248 9628 6276
rect 1946 6236 1952 6248
rect 1859 6208 1952 6236
rect 1946 6196 1952 6208
rect 2004 6236 2010 6248
rect 2222 6245 2228 6248
rect 2216 6236 2228 6245
rect 2004 6208 2029 6236
rect 2183 6208 2228 6236
rect 2004 6196 2010 6208
rect 2216 6199 2228 6208
rect 2222 6196 2228 6199
rect 2280 6196 2286 6248
rect 4062 6236 4068 6248
rect 3252 6208 4068 6236
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6168 1915 6171
rect 1964 6168 1992 6196
rect 3252 6168 3280 6208
rect 4062 6196 4068 6208
rect 4120 6236 4126 6248
rect 4246 6236 4252 6248
rect 4120 6208 4252 6236
rect 4120 6196 4126 6208
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 6972 6208 7849 6236
rect 6972 6196 6978 6208
rect 7837 6205 7849 6208
rect 7883 6236 7895 6239
rect 8386 6236 8392 6248
rect 7883 6208 8392 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9306 6236 9312 6248
rect 9267 6208 9312 6236
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6236 11299 6239
rect 11900 6236 11928 6403
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 13357 6443 13415 6449
rect 13357 6440 13369 6443
rect 12860 6412 13369 6440
rect 12860 6400 12866 6412
rect 13357 6409 13369 6412
rect 13403 6409 13415 6443
rect 13357 6403 13415 6409
rect 11287 6208 11928 6236
rect 12437 6239 12495 6245
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12483 6208 13001 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12989 6205 13001 6208
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 4338 6168 4344 6180
rect 1903 6140 3280 6168
rect 3344 6140 4344 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 3344 6109 3372 6140
rect 4338 6128 4344 6140
rect 4396 6168 4402 6180
rect 4433 6171 4491 6177
rect 4433 6168 4445 6171
rect 4396 6140 4445 6168
rect 4396 6128 4402 6140
rect 4433 6137 4445 6140
rect 4479 6137 4491 6171
rect 4433 6131 4491 6137
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 9447 6171 9505 6177
rect 9447 6168 9459 6171
rect 8904 6140 9459 6168
rect 8904 6128 8910 6140
rect 9447 6137 9459 6140
rect 9493 6137 9505 6171
rect 9447 6131 9505 6137
rect 9950 6128 9956 6180
rect 10008 6168 10014 6180
rect 10410 6168 10416 6180
rect 10008 6140 10416 6168
rect 10008 6128 10014 6140
rect 10410 6128 10416 6140
rect 10468 6168 10474 6180
rect 12452 6168 12480 6199
rect 10468 6140 12480 6168
rect 10468 6128 10474 6140
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 2740 6072 3341 6100
rect 2740 6060 2746 6072
rect 3329 6069 3341 6072
rect 3375 6069 3387 6103
rect 3329 6063 3387 6069
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 4246 6100 4252 6112
rect 4203 6072 4252 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 4246 6060 4252 6072
rect 4304 6100 4310 6112
rect 5258 6100 5264 6112
rect 4304 6072 5264 6100
rect 4304 6060 4310 6072
rect 5258 6060 5264 6072
rect 5316 6100 5322 6112
rect 7098 6100 7104 6112
rect 5316 6072 7104 6100
rect 5316 6060 5322 6072
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 7650 6100 7656 6112
rect 7607 6072 7656 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8754 6100 8760 6112
rect 8067 6072 8760 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10321 6103 10379 6109
rect 10321 6100 10333 6103
rect 10284 6072 10333 6100
rect 10284 6060 10290 6072
rect 10321 6069 10333 6072
rect 10367 6069 10379 6103
rect 10321 6063 10379 6069
rect 11425 6103 11483 6109
rect 11425 6069 11437 6103
rect 11471 6100 11483 6103
rect 12066 6100 12072 6112
rect 11471 6072 12072 6100
rect 11471 6069 11483 6072
rect 11425 6063 11483 6069
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 12621 6103 12679 6109
rect 12621 6069 12633 6103
rect 12667 6100 12679 6103
rect 12986 6100 12992 6112
rect 12667 6072 12992 6100
rect 12667 6069 12679 6072
rect 12621 6063 12679 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 2222 5856 2228 5908
rect 2280 5896 2286 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 2280 5868 2329 5896
rect 2280 5856 2286 5868
rect 2317 5865 2329 5868
rect 2363 5896 2375 5899
rect 3418 5896 3424 5908
rect 2363 5868 3424 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8904 5868 8953 5896
rect 8904 5856 8910 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9858 5896 9864 5908
rect 9088 5868 9864 5896
rect 9088 5856 9094 5868
rect 9858 5856 9864 5868
rect 9916 5896 9922 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 9916 5868 10241 5896
rect 9916 5856 9922 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 10229 5859 10287 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12676 5868 12909 5896
rect 12676 5856 12682 5868
rect 12897 5865 12909 5868
rect 12943 5865 12955 5899
rect 12897 5859 12955 5865
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 8294 5828 8300 5840
rect 7432 5800 8300 5828
rect 7432 5788 7438 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 9824 5800 10057 5828
rect 9824 5788 9830 5800
rect 10045 5797 10057 5800
rect 10091 5797 10103 5831
rect 10318 5828 10324 5840
rect 10279 5800 10324 5828
rect 10045 5791 10103 5797
rect 10318 5788 10324 5800
rect 10376 5828 10382 5840
rect 10502 5828 10508 5840
rect 10376 5800 10508 5828
rect 10376 5788 10382 5800
rect 10502 5788 10508 5800
rect 10560 5788 10566 5840
rect 11784 5831 11842 5837
rect 11784 5797 11796 5831
rect 11830 5828 11842 5831
rect 12158 5828 12164 5840
rect 11830 5800 12164 5828
rect 11830 5797 11842 5800
rect 11784 5791 11842 5797
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 2133 5763 2191 5769
rect 2133 5760 2145 5763
rect 2004 5732 2145 5760
rect 2004 5720 2010 5732
rect 2133 5729 2145 5732
rect 2179 5760 2191 5763
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 2179 5732 4537 5760
rect 2179 5729 2191 5732
rect 2133 5723 2191 5729
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 6822 5760 6828 5772
rect 6687 5732 6828 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8113 5763 8171 5769
rect 8113 5760 8125 5763
rect 7984 5732 8125 5760
rect 7984 5720 7990 5732
rect 8113 5729 8125 5732
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 2409 5695 2467 5701
rect 2409 5692 2421 5695
rect 1820 5664 2421 5692
rect 1820 5652 1826 5664
rect 2409 5661 2421 5664
rect 2455 5692 2467 5695
rect 2682 5692 2688 5704
rect 2455 5664 2688 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 7650 5692 7656 5704
rect 7563 5664 7656 5692
rect 7650 5652 7656 5664
rect 7708 5692 7714 5704
rect 8386 5692 8392 5704
rect 7708 5664 8392 5692
rect 7708 5652 7714 5664
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11480 5664 11529 5692
rect 11480 5652 11486 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 1854 5624 1860 5636
rect 1815 5596 1860 5624
rect 1854 5584 1860 5596
rect 1912 5584 1918 5636
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 2832 5596 3801 5624
rect 2832 5584 2838 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 9769 5627 9827 5633
rect 9769 5593 9781 5627
rect 9815 5624 9827 5627
rect 10870 5624 10876 5636
rect 9815 5596 10876 5624
rect 9815 5593 9827 5596
rect 9769 5587 9827 5593
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5556 2927 5559
rect 3234 5556 3240 5568
rect 2915 5528 3240 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 7098 5556 7104 5568
rect 6871 5528 7104 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7837 5559 7895 5565
rect 7837 5525 7849 5559
rect 7883 5556 7895 5559
rect 8294 5556 8300 5568
rect 7883 5528 8300 5556
rect 7883 5525 7895 5528
rect 7837 5519 7895 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 10689 5559 10747 5565
rect 10689 5556 10701 5559
rect 10468 5528 10701 5556
rect 10468 5516 10474 5528
rect 10689 5525 10701 5528
rect 10735 5525 10747 5559
rect 10689 5519 10747 5525
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 1762 5352 1768 5364
rect 1723 5324 1768 5352
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 1946 5352 1952 5364
rect 1907 5324 1952 5352
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 6822 5352 6828 5364
rect 6687 5324 6828 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 7064 5324 7113 5352
rect 7064 5312 7070 5324
rect 7101 5321 7113 5324
rect 7147 5321 7159 5355
rect 7101 5315 7159 5321
rect 3513 5287 3571 5293
rect 3513 5284 3525 5287
rect 2424 5256 3525 5284
rect 2424 5225 2452 5256
rect 3513 5253 3525 5256
rect 3559 5284 3571 5287
rect 4801 5287 4859 5293
rect 4801 5284 4813 5287
rect 3559 5256 4813 5284
rect 3559 5253 3571 5256
rect 3513 5247 3571 5253
rect 4801 5253 4813 5256
rect 4847 5253 4859 5287
rect 4801 5247 4859 5253
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5216 4031 5219
rect 4062 5216 4068 5228
rect 4019 5188 4068 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 7116 5216 7144 5315
rect 7374 5312 7380 5364
rect 7432 5352 7438 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 7432 5324 7481 5352
rect 7432 5312 7438 5324
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 7469 5315 7527 5321
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 9824 5324 10885 5352
rect 9824 5312 9830 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 11977 5355 12035 5361
rect 11977 5321 11989 5355
rect 12023 5352 12035 5355
rect 12158 5352 12164 5364
rect 12023 5324 12164 5352
rect 12023 5321 12035 5324
rect 11977 5315 12035 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 7742 5284 7748 5296
rect 7703 5256 7748 5284
rect 7742 5244 7748 5256
rect 7800 5244 7806 5296
rect 9950 5284 9956 5296
rect 9911 5256 9956 5284
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 10413 5219 10471 5225
rect 7116 5188 7604 5216
rect 2314 5108 2320 5160
rect 2372 5148 2378 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2372 5120 2513 5148
rect 2372 5108 2378 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 7466 5148 7472 5160
rect 5767 5120 7472 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 4065 5083 4123 5089
rect 4065 5080 4077 5083
rect 3476 5052 4077 5080
rect 3476 5040 3482 5052
rect 4065 5049 4077 5052
rect 4111 5049 4123 5083
rect 7190 5080 7196 5092
rect 4065 5043 4123 5049
rect 4264 5052 7196 5080
rect 2406 5012 2412 5024
rect 2367 4984 2412 5012
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 2866 5012 2872 5024
rect 2827 4984 2872 5012
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 3142 4972 3148 5024
rect 3200 5012 3206 5024
rect 3329 5015 3387 5021
rect 3329 5012 3341 5015
rect 3200 4984 3341 5012
rect 3200 4972 3206 4984
rect 3329 4981 3341 4984
rect 3375 5012 3387 5015
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3375 4984 3985 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 3973 4981 3985 4984
rect 4019 5012 4031 5015
rect 4264 5012 4292 5052
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 7576 5080 7604 5188
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 10594 5216 10600 5228
rect 10459 5188 10600 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 8018 5148 8024 5160
rect 7979 5120 8024 5148
rect 8018 5108 8024 5120
rect 8076 5148 8082 5160
rect 8478 5148 8484 5160
rect 8076 5120 8484 5148
rect 8076 5108 8082 5120
rect 8478 5108 8484 5120
rect 8536 5148 8542 5160
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8536 5120 8677 5148
rect 8536 5108 8542 5120
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9447 5120 9781 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 9769 5117 9781 5120
rect 9815 5148 9827 5151
rect 10502 5148 10508 5160
rect 9815 5120 10508 5148
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12492 5120 13001 5148
rect 12492 5108 12498 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 8205 5083 8263 5089
rect 8205 5080 8217 5083
rect 7576 5052 8217 5080
rect 8205 5049 8217 5052
rect 8251 5049 8263 5083
rect 8205 5043 8263 5049
rect 8297 5083 8355 5089
rect 8297 5049 8309 5083
rect 8343 5080 8355 5083
rect 8386 5080 8392 5092
rect 8343 5052 8392 5080
rect 8343 5049 8355 5052
rect 8297 5043 8355 5049
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 10410 5080 10416 5092
rect 10371 5052 10416 5080
rect 10410 5040 10416 5052
rect 10468 5040 10474 5092
rect 4430 5012 4436 5024
rect 4019 4984 4292 5012
rect 4391 4984 4436 5012
rect 4019 4981 4031 4984
rect 3973 4975 4031 4981
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5442 5012 5448 5024
rect 5307 4984 5448 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 5626 5012 5632 5024
rect 5587 4984 5632 5012
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 6273 5015 6331 5021
rect 6273 4981 6285 5015
rect 6319 5012 6331 5015
rect 7006 5012 7012 5024
rect 6319 4984 7012 5012
rect 6319 4981 6331 4984
rect 6273 4975 6331 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 11422 5012 11428 5024
rect 10284 4984 11428 5012
rect 10284 4972 10290 4984
rect 11422 4972 11428 4984
rect 11480 5012 11486 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11480 4984 11529 5012
rect 11480 4972 11486 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12584 4984 12633 5012
rect 12584 4972 12590 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 1946 4808 1952 4820
rect 1859 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4808 2010 4820
rect 2314 4808 2320 4820
rect 2004 4780 2320 4808
rect 2004 4768 2010 4780
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2682 4808 2688 4820
rect 2643 4780 2688 4808
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 4062 4808 4068 4820
rect 3559 4780 4068 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 5997 4811 6055 4817
rect 5997 4777 6009 4811
rect 6043 4808 6055 4811
rect 6638 4808 6644 4820
rect 6043 4780 6644 4808
rect 6043 4777 6055 4780
rect 5997 4771 6055 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 6825 4811 6883 4817
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 6871 4780 7481 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 7469 4777 7481 4780
rect 7515 4808 7527 4811
rect 7742 4808 7748 4820
rect 7515 4780 7748 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 9858 4808 9864 4820
rect 9819 4780 9864 4808
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 10962 4768 10968 4780
rect 11020 4808 11026 4820
rect 11146 4808 11152 4820
rect 11020 4780 11152 4808
rect 11020 4768 11026 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 2332 4740 2360 4768
rect 2777 4743 2835 4749
rect 2777 4740 2789 4743
rect 2332 4712 2789 4740
rect 2777 4709 2789 4712
rect 2823 4709 2835 4743
rect 2777 4703 2835 4709
rect 4617 4743 4675 4749
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 4798 4740 4804 4752
rect 4663 4712 4804 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 4798 4700 4804 4712
rect 4856 4740 4862 4752
rect 4982 4740 4988 4752
rect 4856 4712 4988 4740
rect 4856 4700 4862 4712
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 7558 4740 7564 4752
rect 7519 4712 7564 4740
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 10686 4700 10692 4752
rect 10744 4740 10750 4752
rect 10781 4743 10839 4749
rect 10781 4740 10793 4743
rect 10744 4712 10793 4740
rect 10744 4700 10750 4712
rect 10781 4709 10793 4712
rect 10827 4709 10839 4743
rect 10781 4703 10839 4709
rect 4338 4632 4344 4684
rect 4396 4672 4402 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 4396 4644 4445 4672
rect 4396 4632 4402 4644
rect 4433 4641 4445 4644
rect 4479 4672 4491 4675
rect 4890 4672 4896 4684
rect 4479 4644 4896 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5776 4644 5825 4672
rect 5776 4632 5782 4644
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 7742 4672 7748 4684
rect 7340 4644 7748 4672
rect 7340 4632 7346 4644
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 8478 4672 8484 4684
rect 8439 4644 8484 4672
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9732 4644 10333 4672
rect 9732 4632 9738 4644
rect 10321 4641 10333 4644
rect 10367 4672 10379 4675
rect 11974 4672 11980 4684
rect 10367 4644 11100 4672
rect 11935 4644 11980 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 2222 4536 2228 4548
rect 2183 4508 2228 4536
rect 2222 4496 2228 4508
rect 2280 4496 2286 4548
rect 4154 4536 4160 4548
rect 4115 4508 4160 4536
rect 4154 4496 4160 4508
rect 4212 4496 4218 4548
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3476 4440 3801 4468
rect 3476 4428 3482 4440
rect 3789 4437 3801 4440
rect 3835 4468 3847 4471
rect 4724 4468 4752 4567
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7432 4576 7481 4604
rect 7432 4564 7438 4576
rect 7469 4573 7481 4576
rect 7515 4604 7527 4607
rect 9398 4604 9404 4616
rect 7515 4576 9404 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 10594 4604 10600 4616
rect 9539 4576 10600 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 11072 4613 11100 4644
rect 11974 4632 11980 4644
rect 12032 4672 12038 4684
rect 12710 4672 12716 4684
rect 12032 4644 12716 4672
rect 12032 4632 12038 4644
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11238 4604 11244 4616
rect 11103 4576 11244 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 5721 4539 5779 4545
rect 5721 4505 5733 4539
rect 5767 4536 5779 4539
rect 6914 4536 6920 4548
rect 5767 4508 6920 4536
rect 5767 4505 5779 4508
rect 5721 4499 5779 4505
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 8386 4536 8392 4548
rect 8299 4508 8392 4536
rect 8386 4496 8392 4508
rect 8444 4536 8450 4548
rect 9582 4536 9588 4548
rect 8444 4508 9588 4536
rect 8444 4496 8450 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 10410 4496 10416 4548
rect 10468 4536 10474 4548
rect 10505 4539 10563 4545
rect 10505 4536 10517 4539
rect 10468 4508 10517 4536
rect 10468 4496 10474 4508
rect 10505 4505 10517 4508
rect 10551 4505 10563 4539
rect 10505 4499 10563 4505
rect 3835 4440 4752 4468
rect 5261 4471 5319 4477
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 5442 4468 5448 4480
rect 5307 4440 5448 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 6457 4471 6515 4477
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6503 4440 7021 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 7009 4437 7021 4440
rect 7055 4468 7067 4471
rect 7190 4468 7196 4480
rect 7055 4440 7196 4468
rect 7055 4437 7067 4440
rect 7009 4431 7067 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 8662 4468 8668 4480
rect 8623 4440 8668 4468
rect 8662 4428 8668 4440
rect 8720 4428 8726 4480
rect 9125 4471 9183 4477
rect 9125 4437 9137 4471
rect 9171 4468 9183 4471
rect 9306 4468 9312 4480
rect 9171 4440 9312 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 12161 4471 12219 4477
rect 12161 4468 12173 4471
rect 11112 4440 12173 4468
rect 11112 4428 11118 4440
rect 12161 4437 12173 4440
rect 12207 4437 12219 4471
rect 12161 4431 12219 4437
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 13265 4471 13323 4477
rect 13265 4468 13277 4471
rect 12308 4440 13277 4468
rect 12308 4428 12314 4440
rect 13265 4437 13277 4440
rect 13311 4437 13323 4471
rect 13265 4431 13323 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 1946 4224 1952 4276
rect 2004 4264 2010 4276
rect 3697 4267 3755 4273
rect 3697 4264 3709 4267
rect 2004 4236 3709 4264
rect 2004 4224 2010 4236
rect 3697 4233 3709 4236
rect 3743 4233 3755 4267
rect 4338 4264 4344 4276
rect 4299 4236 4344 4264
rect 3697 4227 3755 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 5261 4267 5319 4273
rect 5261 4233 5273 4267
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 5276 4140 5304 4227
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 5776 4236 6193 4264
rect 5776 4224 5782 4236
rect 6181 4233 6193 4236
rect 6227 4264 6239 4267
rect 6822 4264 6828 4276
rect 6227 4236 6828 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7558 4264 7564 4276
rect 7156 4236 7564 4264
rect 7156 4224 7162 4236
rect 7558 4224 7564 4236
rect 7616 4264 7622 4276
rect 7837 4267 7895 4273
rect 7837 4264 7849 4267
rect 7616 4236 7849 4264
rect 7616 4224 7622 4236
rect 7837 4233 7849 4236
rect 7883 4233 7895 4267
rect 7837 4227 7895 4233
rect 8297 4267 8355 4273
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8478 4264 8484 4276
rect 8343 4236 8484 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 9677 4267 9735 4273
rect 9677 4233 9689 4267
rect 9723 4264 9735 4267
rect 9723 4236 10640 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 6641 4199 6699 4205
rect 6641 4196 6653 4199
rect 5368 4168 6653 4196
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 5166 4128 5172 4140
rect 4212 4100 5172 4128
rect 4212 4088 4218 4100
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2363 4032 2728 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 2406 3992 2412 4004
rect 1903 3964 2412 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 2406 3952 2412 3964
rect 2464 3992 2470 4004
rect 2562 3995 2620 4001
rect 2562 3992 2574 3995
rect 2464 3964 2574 3992
rect 2464 3952 2470 3964
rect 2562 3961 2574 3964
rect 2608 3961 2620 3995
rect 2562 3955 2620 3961
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 2700 3924 2728 4032
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5368 4060 5396 4168
rect 6641 4165 6653 4168
rect 6687 4196 6699 4199
rect 7374 4196 7380 4208
rect 6687 4168 7380 4196
rect 6687 4165 6699 4168
rect 6641 4159 6699 4165
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 10045 4199 10103 4205
rect 10045 4165 10057 4199
rect 10091 4165 10103 4199
rect 10045 4159 10103 4165
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4128 5690 4140
rect 6899 4131 6957 4137
rect 6899 4128 6911 4131
rect 5684 4100 6911 4128
rect 5684 4088 5690 4100
rect 6899 4097 6911 4100
rect 6945 4097 6957 4131
rect 6899 4091 6957 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7558 4128 7564 4140
rect 7515 4100 7564 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7558 4088 7564 4100
rect 7616 4128 7622 4140
rect 8202 4128 8208 4140
rect 7616 4100 8208 4128
rect 7616 4088 7622 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9306 4128 9312 4140
rect 8987 4100 9312 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9306 4088 9312 4100
rect 9364 4128 9370 4140
rect 10060 4128 10088 4159
rect 10612 4137 10640 4236
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 10965 4267 11023 4273
rect 10965 4264 10977 4267
rect 10744 4236 10977 4264
rect 10744 4224 10750 4236
rect 10965 4233 10977 4236
rect 11011 4233 11023 4267
rect 11974 4264 11980 4276
rect 11935 4236 11980 4264
rect 10965 4227 11023 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 13170 4264 13176 4276
rect 13131 4236 13176 4264
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 9364 4100 10088 4128
rect 10597 4131 10655 4137
rect 9364 4088 9370 4100
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11054 4088 11060 4140
rect 11112 4088 11118 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 11204 4100 11345 4128
rect 11204 4088 11210 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 5132 4032 5396 4060
rect 5132 4020 5138 4032
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 8463 4063 8521 4069
rect 8463 4060 8475 4063
rect 7432 4032 8475 4060
rect 7432 4020 7438 4032
rect 8463 4029 8475 4032
rect 8509 4060 8521 4063
rect 9398 4060 9404 4072
rect 8509 4032 9404 4060
rect 8509 4029 8521 4032
rect 8463 4023 8521 4029
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 5813 3995 5871 4001
rect 5813 3992 5825 3995
rect 5000 3964 5825 3992
rect 5000 3936 5028 3964
rect 5813 3961 5825 3964
rect 5859 3961 5871 3995
rect 5813 3955 5871 3961
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 6972 3964 7205 3992
rect 6972 3952 6978 3964
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7193 3955 7251 3961
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 8938 3992 8944 4004
rect 8352 3964 8944 3992
rect 8352 3952 8358 3964
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3961 9091 3995
rect 9692 3992 9720 4023
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 11072 4060 11100 4088
rect 9824 4032 11100 4060
rect 9824 4020 9830 4032
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12618 4060 12624 4072
rect 12492 4032 12624 4060
rect 12492 4020 12498 4032
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 9033 3955 9091 3961
rect 9600 3964 9720 3992
rect 10321 3995 10379 4001
rect 4338 3924 4344 3936
rect 2271 3896 4344 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4798 3924 4804 3936
rect 4755 3896 4804 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 7064 3896 7389 3924
rect 7064 3884 7070 3896
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 9048 3924 9076 3955
rect 9600 3936 9628 3964
rect 10321 3961 10333 3995
rect 10367 3961 10379 3995
rect 10321 3955 10379 3961
rect 8720 3896 9076 3924
rect 9493 3927 9551 3933
rect 8720 3884 8726 3896
rect 9493 3893 9505 3927
rect 9539 3924 9551 3927
rect 9582 3924 9588 3936
rect 9539 3896 9588 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9732 3896 9781 3924
rect 9732 3884 9738 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 9769 3887 9827 3893
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10336 3924 10364 3955
rect 12710 3952 12716 4004
rect 12768 3992 12774 4004
rect 13541 3995 13599 4001
rect 13541 3992 13553 3995
rect 12768 3964 13553 3992
rect 12768 3952 12774 3964
rect 13541 3961 13553 3964
rect 13587 3961 13599 3995
rect 13541 3955 13599 3961
rect 10100 3896 10364 3924
rect 10505 3927 10563 3933
rect 10100 3884 10106 3896
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10686 3924 10692 3936
rect 10551 3896 10692 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 12618 3924 12624 3936
rect 12579 3896 12624 3924
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 7558 3720 7564 3732
rect 6840 3692 7564 3720
rect 2958 3652 2964 3664
rect 2919 3624 2964 3652
rect 2958 3612 2964 3624
rect 3016 3612 3022 3664
rect 5442 3661 5448 3664
rect 5436 3652 5448 3661
rect 5355 3624 5448 3652
rect 5436 3615 5448 3624
rect 5500 3652 5506 3664
rect 6840 3652 6868 3692
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8202 3720 8208 3732
rect 8163 3692 8208 3720
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8757 3723 8815 3729
rect 8757 3689 8769 3723
rect 8803 3720 8815 3723
rect 8846 3720 8852 3732
rect 8803 3692 8852 3720
rect 8803 3689 8815 3692
rect 8757 3683 8815 3689
rect 8846 3680 8852 3692
rect 8904 3720 8910 3732
rect 11609 3723 11667 3729
rect 11609 3720 11621 3723
rect 8904 3692 11621 3720
rect 8904 3680 8910 3692
rect 11609 3689 11621 3692
rect 11655 3720 11667 3723
rect 11655 3692 13492 3720
rect 11655 3689 11667 3692
rect 11609 3683 11667 3689
rect 7098 3652 7104 3664
rect 5500 3624 6868 3652
rect 7059 3624 7104 3652
rect 5442 3612 5448 3615
rect 5500 3612 5506 3624
rect 7098 3612 7104 3624
rect 7156 3612 7162 3664
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 7926 3652 7932 3664
rect 7524 3624 7932 3652
rect 7524 3612 7530 3624
rect 7926 3612 7932 3624
rect 7984 3652 7990 3664
rect 8021 3655 8079 3661
rect 8021 3652 8033 3655
rect 7984 3624 8033 3652
rect 7984 3612 7990 3624
rect 8021 3621 8033 3624
rect 8067 3621 8079 3655
rect 8021 3615 8079 3621
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8996 3624 9045 3652
rect 8996 3612 9002 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9398 3652 9404 3664
rect 9359 3624 9404 3652
rect 9033 3615 9091 3621
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 10042 3652 10048 3664
rect 10003 3624 10048 3652
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 10410 3612 10416 3664
rect 10468 3661 10474 3664
rect 10468 3655 10532 3661
rect 10468 3621 10486 3655
rect 10520 3621 10532 3655
rect 10468 3615 10532 3621
rect 10468 3612 10474 3615
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13320 3624 13365 3652
rect 13320 3612 13326 3624
rect 2976 3584 3004 3612
rect 3142 3584 3148 3596
rect 2976 3556 3148 3584
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 4028 3556 4077 3584
rect 4028 3544 4034 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2590 3516 2596 3528
rect 1820 3488 2596 3516
rect 1820 3476 1826 3488
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3485 3111 3519
rect 4080 3516 4108 3547
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4396 3556 4629 3584
rect 4396 3544 4402 3556
rect 4617 3553 4629 3556
rect 4663 3584 4675 3587
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 4663 3556 5181 3584
rect 4663 3553 4675 3556
rect 4617 3547 4675 3553
rect 5169 3553 5181 3556
rect 5215 3584 5227 3587
rect 6270 3584 6276 3596
rect 5215 3556 6276 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 7116 3584 7144 3612
rect 8294 3584 8300 3596
rect 7116 3556 8300 3584
rect 8294 3544 8300 3556
rect 8352 3584 8358 3596
rect 8662 3584 8668 3596
rect 8352 3556 8668 3584
rect 8352 3544 8358 3556
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 13078 3584 13084 3596
rect 13039 3556 13084 3584
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 13354 3584 13360 3596
rect 13267 3556 13360 3584
rect 13354 3544 13360 3556
rect 13412 3584 13418 3596
rect 13464 3584 13492 3692
rect 13412 3556 13492 3584
rect 13412 3544 13418 3556
rect 4706 3516 4712 3528
rect 4080 3488 4712 3516
rect 3053 3479 3111 3485
rect 2501 3451 2559 3457
rect 2501 3417 2513 3451
rect 2547 3448 2559 3451
rect 2682 3448 2688 3460
rect 2547 3420 2688 3448
rect 2547 3417 2559 3420
rect 2501 3411 2559 3417
rect 2682 3408 2688 3420
rect 2740 3408 2746 3460
rect 2317 3383 2375 3389
rect 2317 3349 2329 3383
rect 2363 3380 2375 3383
rect 2406 3380 2412 3392
rect 2363 3352 2412 3380
rect 2363 3349 2375 3352
rect 2317 3343 2375 3349
rect 2406 3340 2412 3352
rect 2464 3380 2470 3392
rect 3068 3380 3096 3479
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12492 3488 12537 3516
rect 12492 3476 12498 3488
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 6972 3420 7757 3448
rect 6972 3408 6978 3420
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 12802 3448 12808 3460
rect 12763 3420 12808 3448
rect 7745 3411 7803 3417
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 3418 3380 3424 3392
rect 2464 3352 3424 3380
rect 2464 3340 2470 3352
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 4062 3380 4068 3392
rect 3927 3352 4068 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4982 3380 4988 3392
rect 4943 3352 4988 3380
rect 4982 3340 4988 3352
rect 5040 3380 5046 3392
rect 6549 3383 6607 3389
rect 6549 3380 6561 3383
rect 5040 3352 6561 3380
rect 5040 3340 5046 3352
rect 6549 3349 6561 3352
rect 6595 3349 6607 3383
rect 6549 3343 6607 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 2832 3148 2877 3176
rect 2832 3136 2838 3148
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3200 3148 3709 3176
rect 3200 3136 3206 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6917 3179 6975 3185
rect 6917 3176 6929 3179
rect 5776 3148 6929 3176
rect 5776 3136 5782 3148
rect 6917 3145 6929 3148
rect 6963 3145 6975 3179
rect 6917 3139 6975 3145
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8202 3176 8208 3188
rect 7975 3148 8208 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9640 3148 10057 3176
rect 9640 3136 9646 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 10410 3136 10416 3188
rect 10468 3176 10474 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10468 3148 10977 3176
rect 10468 3136 10474 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 13354 3176 13360 3188
rect 13315 3148 13360 3176
rect 10965 3139 11023 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 6270 3108 6276 3120
rect 1452 3080 2636 3108
rect 6183 3080 6276 3108
rect 1452 3068 1458 3080
rect 1578 3040 1584 3052
rect 1539 3012 1584 3040
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 2608 3049 2636 3080
rect 6270 3068 6276 3080
rect 6328 3108 6334 3120
rect 8481 3111 8539 3117
rect 8481 3108 8493 3111
rect 6328 3080 8493 3108
rect 6328 3068 6334 3080
rect 8481 3077 8493 3080
rect 8527 3108 8539 3111
rect 8527 3080 8708 3108
rect 8527 3077 8539 3080
rect 8481 3071 8539 3077
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 3050 3040 3056 3052
rect 2639 3012 3056 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 3050 3000 3056 3012
rect 3108 3040 3114 3052
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 3108 3012 3157 3040
rect 3108 3000 3114 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6687 3012 7481 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 7469 3009 7481 3012
rect 7515 3040 7527 3043
rect 7558 3040 7564 3052
rect 7515 3012 7564 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 8680 3049 8708 3080
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 12161 3111 12219 3117
rect 12161 3108 12173 3111
rect 10928 3080 12173 3108
rect 10928 3068 10934 3080
rect 12161 3077 12173 3080
rect 12207 3077 12219 3111
rect 12161 3071 12219 3077
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 12176 3040 12204 3071
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 13725 3111 13783 3117
rect 13725 3108 13737 3111
rect 13136 3080 13737 3108
rect 13136 3068 13142 3080
rect 13725 3077 13737 3080
rect 13771 3077 13783 3111
rect 13725 3071 13783 3077
rect 13262 3040 13268 3052
rect 12176 3012 13268 3040
rect 8665 3003 8723 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2866 2972 2872 2984
rect 1443 2944 2872 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3970 2972 3976 2984
rect 3068 2944 3976 2972
rect 3068 2916 3096 2944
rect 3970 2932 3976 2944
rect 4028 2972 4034 2984
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 4028 2944 4077 2972
rect 4028 2932 4034 2944
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2972 4307 2975
rect 4338 2972 4344 2984
rect 4295 2944 4344 2972
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4516 2975 4574 2981
rect 4516 2941 4528 2975
rect 4562 2972 4574 2975
rect 4982 2972 4988 2984
rect 4562 2944 4988 2972
rect 4562 2941 4574 2944
rect 4516 2935 4574 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 7190 2972 7196 2984
rect 7151 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 2958 2904 2964 2916
rect 2271 2876 2964 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 3050 2864 3056 2916
rect 3108 2864 3114 2916
rect 3234 2904 3240 2916
rect 3195 2876 3240 2904
rect 3234 2864 3240 2876
rect 3292 2864 3298 2916
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 3418 2904 3424 2916
rect 3375 2876 3424 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 3418 2864 3424 2876
rect 3476 2864 3482 2916
rect 7374 2904 7380 2916
rect 7335 2876 7380 2904
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 3252 2836 3280 2864
rect 2740 2808 3280 2836
rect 2740 2796 2746 2808
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5500 2808 5641 2836
rect 5500 2796 5506 2808
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 8680 2836 8708 3003
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 9306 2972 9312 2984
rect 8812 2944 9312 2972
rect 8812 2932 8818 2944
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11330 2972 11336 2984
rect 11195 2944 11336 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11330 2932 11336 2944
rect 11388 2972 11394 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11388 2944 11713 2972
rect 11388 2932 11394 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12492 2944 13001 2972
rect 12492 2932 12498 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 8846 2864 8852 2916
rect 8904 2913 8910 2916
rect 8904 2907 8968 2913
rect 8904 2873 8922 2907
rect 8956 2873 8968 2907
rect 8904 2867 8968 2873
rect 8904 2864 8910 2867
rect 10226 2836 10232 2848
rect 8680 2808 10232 2836
rect 5629 2799 5687 2805
rect 10226 2796 10232 2808
rect 10284 2836 10290 2848
rect 10597 2839 10655 2845
rect 10597 2836 10609 2839
rect 10284 2808 10609 2836
rect 10284 2796 10290 2808
rect 10597 2805 10609 2808
rect 10643 2805 10655 2839
rect 10597 2799 10655 2805
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 11514 2836 11520 2848
rect 11379 2808 11520 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 5534 2632 5540 2644
rect 5495 2604 5540 2632
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 7466 2632 7472 2644
rect 6411 2604 7472 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8294 2632 8300 2644
rect 8220 2604 8300 2632
rect 2038 2524 2044 2576
rect 2096 2564 2102 2576
rect 2961 2567 3019 2573
rect 2961 2564 2973 2567
rect 2096 2536 2973 2564
rect 2096 2524 2102 2536
rect 566 2320 572 2372
rect 624 2360 630 2372
rect 2240 2369 2268 2536
rect 2961 2533 2973 2536
rect 3007 2533 3019 2567
rect 2961 2527 3019 2533
rect 3050 2524 3056 2576
rect 3108 2524 3114 2576
rect 3513 2567 3571 2573
rect 3513 2533 3525 2567
rect 3559 2564 3571 2567
rect 4062 2564 4068 2576
rect 3559 2536 4068 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3068 2496 3096 2524
rect 2823 2468 3096 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 2225 2363 2283 2369
rect 2225 2360 2237 2363
rect 624 2332 2237 2360
rect 624 2320 630 2332
rect 2225 2329 2237 2332
rect 2271 2329 2283 2363
rect 2225 2323 2283 2329
rect 2501 2363 2559 2369
rect 2501 2329 2513 2363
rect 2547 2360 2559 2363
rect 2682 2360 2688 2372
rect 2547 2332 2688 2360
rect 2547 2329 2559 2332
rect 2501 2323 2559 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 1949 2295 2007 2301
rect 1949 2261 1961 2295
rect 1995 2292 2007 2295
rect 2792 2292 2820 2459
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3528 2428 3556 2527
rect 4062 2524 4068 2536
rect 4120 2564 4126 2576
rect 4402 2567 4460 2573
rect 4402 2564 4414 2567
rect 4120 2536 4414 2564
rect 4120 2524 4126 2536
rect 4402 2533 4414 2536
rect 4448 2564 4460 2567
rect 5442 2564 5448 2576
rect 4448 2536 5448 2564
rect 4448 2533 4460 2536
rect 4402 2527 4460 2533
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 3927 2468 4169 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4157 2465 4169 2468
rect 4203 2496 4215 2499
rect 4246 2496 4252 2508
rect 4203 2468 4252 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 7834 2496 7840 2508
rect 7392 2468 7840 2496
rect 7392 2440 7420 2468
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 3099 2400 3556 2428
rect 6733 2431 6791 2437
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7374 2428 7380 2440
rect 6779 2400 7380 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8220 2428 8248 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10100 2604 10425 2632
rect 10100 2592 10106 2604
rect 10413 2601 10425 2604
rect 10459 2632 10471 2635
rect 11057 2635 11115 2641
rect 11057 2632 11069 2635
rect 10459 2604 11069 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 11057 2601 11069 2604
rect 11103 2601 11115 2635
rect 11330 2632 11336 2644
rect 11057 2595 11115 2601
rect 11164 2604 11336 2632
rect 11164 2573 11192 2604
rect 11330 2592 11336 2604
rect 11388 2632 11394 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11388 2604 11529 2632
rect 11388 2592 11394 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2533 11207 2567
rect 11149 2527 11207 2533
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8352 2468 8493 2496
rect 8352 2456 8358 2468
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8527 2468 9045 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 10870 2496 10876 2508
rect 10091 2468 10876 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2496 12682 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12676 2468 13185 2496
rect 12676 2456 12682 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 7607 2400 8401 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8389 2397 8401 2400
rect 8435 2428 8447 2431
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 8435 2400 9413 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 9401 2397 9413 2400
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 7006 2360 7012 2372
rect 6967 2332 7012 2360
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 8665 2363 8723 2369
rect 8665 2360 8677 2363
rect 8260 2332 8677 2360
rect 8260 2320 8266 2332
rect 8665 2329 8677 2332
rect 8711 2329 8723 2363
rect 10594 2360 10600 2372
rect 10555 2332 10600 2360
rect 8665 2323 8723 2329
rect 10594 2320 10600 2332
rect 10652 2320 10658 2372
rect 12802 2292 12808 2304
rect 1995 2264 2820 2292
rect 12763 2264 12808 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 6638 1368 6644 1420
rect 6696 1408 6702 1420
rect 8938 1408 8944 1420
rect 6696 1380 8944 1408
rect 6696 1368 6702 1380
rect 8938 1368 8944 1380
rect 8996 1368 9002 1420
<< via1 >>
rect 5540 37680 5592 37732
rect 6368 37680 6420 37732
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 12348 36864 12400 36916
rect 11336 36660 11388 36712
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 10968 36363 11020 36372
rect 10968 36329 10977 36363
rect 10977 36329 11011 36363
rect 11011 36329 11020 36363
rect 10968 36320 11020 36329
rect 13452 36320 13504 36372
rect 10784 36227 10836 36236
rect 10784 36193 10793 36227
rect 10793 36193 10827 36227
rect 10827 36193 10836 36227
rect 10784 36184 10836 36193
rect 12256 36184 12308 36236
rect 4344 36023 4396 36032
rect 4344 35989 4353 36023
rect 4353 35989 4387 36023
rect 4387 35989 4396 36023
rect 4344 35980 4396 35989
rect 4620 35980 4672 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 8208 35776 8260 35828
rect 9312 35776 9364 35828
rect 10692 35776 10744 35828
rect 11060 35776 11112 35828
rect 13728 35776 13780 35828
rect 3976 35708 4028 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 4528 35683 4580 35692
rect 4528 35649 4537 35683
rect 4537 35649 4571 35683
rect 4571 35649 4580 35683
rect 4528 35640 4580 35649
rect 4620 35683 4672 35692
rect 4620 35649 4629 35683
rect 4629 35649 4663 35683
rect 4663 35649 4672 35683
rect 4620 35640 4672 35649
rect 1768 35572 1820 35624
rect 8392 35615 8444 35624
rect 8392 35581 8401 35615
rect 8401 35581 8435 35615
rect 8435 35581 8444 35615
rect 8392 35572 8444 35581
rect 8576 35572 8628 35624
rect 11152 35615 11204 35624
rect 11152 35581 11161 35615
rect 11161 35581 11195 35615
rect 11195 35581 11204 35615
rect 11152 35572 11204 35581
rect 2228 35479 2280 35488
rect 2228 35445 2237 35479
rect 2237 35445 2271 35479
rect 2271 35445 2280 35479
rect 2228 35436 2280 35445
rect 4804 35436 4856 35488
rect 4988 35436 5040 35488
rect 9864 35479 9916 35488
rect 9864 35445 9873 35479
rect 9873 35445 9907 35479
rect 9907 35445 9916 35479
rect 9864 35436 9916 35445
rect 10692 35436 10744 35488
rect 12256 35436 12308 35488
rect 13268 35436 13320 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 7932 35232 7984 35284
rect 9496 35232 9548 35284
rect 9956 35232 10008 35284
rect 11152 35232 11204 35284
rect 11520 35232 11572 35284
rect 13360 35275 13412 35284
rect 13360 35241 13369 35275
rect 13369 35241 13403 35275
rect 13403 35241 13412 35275
rect 13360 35232 13412 35241
rect 2504 35164 2556 35216
rect 5448 35164 5500 35216
rect 7840 35096 7892 35148
rect 9772 35096 9824 35148
rect 10784 35139 10836 35148
rect 10784 35105 10793 35139
rect 10793 35105 10827 35139
rect 10827 35105 10836 35139
rect 10784 35096 10836 35105
rect 12072 35096 12124 35148
rect 13176 35139 13228 35148
rect 13176 35105 13185 35139
rect 13185 35105 13219 35139
rect 13219 35105 13228 35139
rect 13176 35096 13228 35105
rect 2228 35028 2280 35080
rect 2412 35028 2464 35080
rect 2964 35028 3016 35080
rect 4896 35028 4948 35080
rect 1768 34892 1820 34944
rect 2228 34935 2280 34944
rect 2228 34901 2237 34935
rect 2237 34901 2271 34935
rect 2271 34901 2280 34935
rect 2228 34892 2280 34901
rect 3240 34935 3292 34944
rect 3240 34901 3249 34935
rect 3249 34901 3283 34935
rect 3283 34901 3292 34935
rect 3240 34892 3292 34901
rect 4620 34892 4672 34944
rect 7012 34935 7064 34944
rect 7012 34901 7021 34935
rect 7021 34901 7055 34935
rect 7055 34901 7064 34935
rect 7012 34892 7064 34901
rect 8852 34892 8904 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 2504 34731 2556 34740
rect 2504 34697 2513 34731
rect 2513 34697 2547 34731
rect 2547 34697 2556 34731
rect 2504 34688 2556 34697
rect 3240 34688 3292 34740
rect 7840 34731 7892 34740
rect 7840 34697 7849 34731
rect 7849 34697 7883 34731
rect 7883 34697 7892 34731
rect 7840 34688 7892 34697
rect 8760 34688 8812 34740
rect 10324 34688 10376 34740
rect 13636 34731 13688 34740
rect 13636 34697 13645 34731
rect 13645 34697 13679 34731
rect 13679 34697 13688 34731
rect 13636 34688 13688 34697
rect 3148 34552 3200 34604
rect 3424 34552 3476 34604
rect 5080 34620 5132 34672
rect 6736 34620 6788 34672
rect 8484 34663 8536 34672
rect 8484 34629 8493 34663
rect 8493 34629 8527 34663
rect 8527 34629 8536 34663
rect 8484 34620 8536 34629
rect 4528 34552 4580 34604
rect 8852 34552 8904 34604
rect 4344 34484 4396 34536
rect 4620 34527 4672 34536
rect 4620 34493 4629 34527
rect 4629 34493 4663 34527
rect 4663 34493 4672 34527
rect 4620 34484 4672 34493
rect 5448 34527 5500 34536
rect 5448 34493 5457 34527
rect 5457 34493 5491 34527
rect 5491 34493 5500 34527
rect 5448 34484 5500 34493
rect 7104 34484 7156 34536
rect 8576 34484 8628 34536
rect 10140 34484 10192 34536
rect 11520 34484 11572 34536
rect 12072 34527 12124 34536
rect 12072 34493 12081 34527
rect 12081 34493 12115 34527
rect 12115 34493 12124 34527
rect 12072 34484 12124 34493
rect 13176 34527 13228 34536
rect 13176 34493 13185 34527
rect 13185 34493 13219 34527
rect 13219 34493 13228 34527
rect 13176 34484 13228 34493
rect 7012 34416 7064 34468
rect 7288 34416 7340 34468
rect 3240 34348 3292 34400
rect 4804 34348 4856 34400
rect 4896 34348 4948 34400
rect 6092 34348 6144 34400
rect 6920 34348 6972 34400
rect 11244 34416 11296 34468
rect 8852 34348 8904 34400
rect 9772 34391 9824 34400
rect 9772 34357 9781 34391
rect 9781 34357 9815 34391
rect 9815 34357 9824 34391
rect 9772 34348 9824 34357
rect 10416 34348 10468 34400
rect 10784 34348 10836 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 2228 34187 2280 34196
rect 2228 34153 2237 34187
rect 2237 34153 2271 34187
rect 2271 34153 2280 34187
rect 2228 34144 2280 34153
rect 5448 34144 5500 34196
rect 14188 34144 14240 34196
rect 2780 34076 2832 34128
rect 4620 34119 4672 34128
rect 4620 34085 4654 34119
rect 4654 34085 4672 34119
rect 4620 34076 4672 34085
rect 6920 34076 6972 34128
rect 2044 34051 2096 34060
rect 2044 34017 2053 34051
rect 2053 34017 2087 34051
rect 2087 34017 2096 34051
rect 2044 34008 2096 34017
rect 4160 34008 4212 34060
rect 4896 34008 4948 34060
rect 10232 34076 10284 34128
rect 9956 34051 10008 34060
rect 9956 34017 9990 34051
rect 9990 34017 10008 34051
rect 12716 34051 12768 34060
rect 9956 34008 10008 34017
rect 12716 34017 12725 34051
rect 12725 34017 12759 34051
rect 12759 34017 12768 34051
rect 12716 34008 12768 34017
rect 2964 33940 3016 33992
rect 6092 33940 6144 33992
rect 1768 33915 1820 33924
rect 1768 33881 1777 33915
rect 1777 33881 1811 33915
rect 1811 33881 1820 33915
rect 1768 33872 1820 33881
rect 4344 33804 4396 33856
rect 8852 33847 8904 33856
rect 8852 33813 8861 33847
rect 8861 33813 8895 33847
rect 8895 33813 8904 33847
rect 8852 33804 8904 33813
rect 9496 33804 9548 33856
rect 10968 33804 11020 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 2780 33600 2832 33652
rect 7104 33643 7156 33652
rect 7104 33609 7113 33643
rect 7113 33609 7147 33643
rect 7147 33609 7156 33643
rect 7104 33600 7156 33609
rect 11980 33600 12032 33652
rect 13636 33643 13688 33652
rect 13636 33609 13645 33643
rect 13645 33609 13679 33643
rect 13679 33609 13688 33643
rect 13636 33600 13688 33609
rect 1676 33396 1728 33448
rect 4160 33396 4212 33448
rect 4344 33439 4396 33448
rect 4344 33405 4378 33439
rect 4378 33405 4396 33439
rect 4344 33396 4396 33405
rect 6920 33396 6972 33448
rect 8208 33396 8260 33448
rect 8484 33439 8536 33448
rect 8484 33405 8493 33439
rect 8493 33405 8527 33439
rect 8527 33405 8536 33439
rect 8484 33396 8536 33405
rect 10232 33396 10284 33448
rect 13452 33439 13504 33448
rect 2964 33328 3016 33380
rect 1676 33260 1728 33312
rect 7104 33328 7156 33380
rect 7564 33371 7616 33380
rect 7564 33337 7573 33371
rect 7573 33337 7607 33371
rect 7607 33337 7616 33371
rect 7564 33328 7616 33337
rect 7656 33371 7708 33380
rect 7656 33337 7665 33371
rect 7665 33337 7699 33371
rect 7699 33337 7708 33371
rect 8852 33371 8904 33380
rect 7656 33328 7708 33337
rect 8852 33337 8886 33371
rect 8886 33337 8904 33371
rect 8852 33328 8904 33337
rect 6092 33260 6144 33312
rect 13452 33405 13461 33439
rect 13461 33405 13495 33439
rect 13495 33405 13504 33439
rect 13452 33396 13504 33405
rect 9680 33260 9732 33312
rect 10232 33260 10284 33312
rect 11428 33260 11480 33312
rect 12716 33303 12768 33312
rect 12716 33269 12725 33303
rect 12725 33269 12759 33303
rect 12759 33269 12768 33303
rect 12716 33260 12768 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 1676 33056 1728 33108
rect 4620 33099 4672 33108
rect 4620 33065 4629 33099
rect 4629 33065 4663 33099
rect 4663 33065 4672 33099
rect 4620 33056 4672 33065
rect 4712 33056 4764 33108
rect 5724 33056 5776 33108
rect 6736 33056 6788 33108
rect 7656 33056 7708 33108
rect 2688 32988 2740 33040
rect 2780 32988 2832 33040
rect 6644 32988 6696 33040
rect 8116 33031 8168 33040
rect 8116 32997 8125 33031
rect 8125 32997 8159 33031
rect 8159 32997 8168 33031
rect 8116 32988 8168 32997
rect 8852 33056 8904 33108
rect 10048 33056 10100 33108
rect 10968 33056 11020 33108
rect 8760 32988 8812 33040
rect 9680 32988 9732 33040
rect 9956 33031 10008 33040
rect 9956 32997 9965 33031
rect 9965 32997 9999 33031
rect 9999 32997 10008 33031
rect 9956 32988 10008 32997
rect 3148 32920 3200 32972
rect 4344 32920 4396 32972
rect 6184 32920 6236 32972
rect 3240 32852 3292 32904
rect 4896 32852 4948 32904
rect 6920 32920 6972 32972
rect 10232 32920 10284 32972
rect 10784 32920 10836 32972
rect 8116 32895 8168 32904
rect 2412 32827 2464 32836
rect 2412 32793 2421 32827
rect 2421 32793 2455 32827
rect 2455 32793 2464 32827
rect 2412 32784 2464 32793
rect 3516 32784 3568 32836
rect 8116 32861 8125 32895
rect 8125 32861 8159 32895
rect 8159 32861 8168 32895
rect 8116 32852 8168 32861
rect 6736 32784 6788 32836
rect 7288 32784 7340 32836
rect 6092 32759 6144 32768
rect 6092 32725 6101 32759
rect 6101 32725 6135 32759
rect 6135 32725 6144 32759
rect 6092 32716 6144 32725
rect 7104 32759 7156 32768
rect 7104 32725 7113 32759
rect 7113 32725 7147 32759
rect 7147 32725 7156 32759
rect 7104 32716 7156 32725
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 2044 32512 2096 32564
rect 4344 32512 4396 32564
rect 4620 32512 4672 32564
rect 8300 32555 8352 32564
rect 8300 32521 8309 32555
rect 8309 32521 8343 32555
rect 8343 32521 8352 32555
rect 8300 32512 8352 32521
rect 8392 32512 8444 32564
rect 8668 32512 8720 32564
rect 9496 32555 9548 32564
rect 3240 32444 3292 32496
rect 4896 32444 4948 32496
rect 5264 32487 5316 32496
rect 5264 32453 5273 32487
rect 5273 32453 5307 32487
rect 5307 32453 5316 32487
rect 5264 32444 5316 32453
rect 8760 32444 8812 32496
rect 1584 32419 1636 32428
rect 1584 32385 1593 32419
rect 1593 32385 1627 32419
rect 1627 32385 1636 32419
rect 1584 32376 1636 32385
rect 3976 32376 4028 32428
rect 5724 32419 5776 32428
rect 5724 32385 5733 32419
rect 5733 32385 5767 32419
rect 5767 32385 5776 32419
rect 5724 32376 5776 32385
rect 1400 32351 1452 32360
rect 1400 32317 1409 32351
rect 1409 32317 1443 32351
rect 1443 32317 1452 32351
rect 1400 32308 1452 32317
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 4160 32308 4212 32360
rect 5448 32308 5500 32360
rect 6000 32308 6052 32360
rect 3516 32240 3568 32292
rect 7656 32308 7708 32360
rect 9496 32521 9505 32555
rect 9505 32521 9539 32555
rect 9539 32521 9548 32555
rect 9496 32512 9548 32521
rect 10232 32512 10284 32564
rect 10784 32555 10836 32564
rect 10784 32521 10793 32555
rect 10793 32521 10827 32555
rect 10827 32521 10836 32555
rect 10784 32512 10836 32521
rect 12164 32512 12216 32564
rect 10048 32419 10100 32428
rect 10048 32385 10057 32419
rect 10057 32385 10091 32419
rect 10091 32385 10100 32419
rect 10048 32376 10100 32385
rect 10968 32351 11020 32360
rect 2964 32172 3016 32224
rect 8484 32240 8536 32292
rect 9404 32240 9456 32292
rect 10968 32317 10977 32351
rect 10977 32317 11011 32351
rect 11011 32317 11020 32351
rect 10968 32308 11020 32317
rect 5264 32172 5316 32224
rect 6092 32172 6144 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 1400 31968 1452 32020
rect 2044 32011 2096 32020
rect 2044 31977 2053 32011
rect 2053 31977 2087 32011
rect 2087 31977 2096 32011
rect 2044 31968 2096 31977
rect 2964 31968 3016 32020
rect 3976 31968 4028 32020
rect 5264 32011 5316 32020
rect 5264 31977 5273 32011
rect 5273 31977 5307 32011
rect 5307 31977 5316 32011
rect 5264 31968 5316 31977
rect 6184 31968 6236 32020
rect 6644 31968 6696 32020
rect 6736 31968 6788 32020
rect 7104 31968 7156 32020
rect 9404 32011 9456 32020
rect 9404 31977 9413 32011
rect 9413 31977 9447 32011
rect 9447 31977 9456 32011
rect 9404 31968 9456 31977
rect 3148 31900 3200 31952
rect 7196 31943 7248 31952
rect 7196 31909 7205 31943
rect 7205 31909 7239 31943
rect 7239 31909 7248 31943
rect 7196 31900 7248 31909
rect 7380 31943 7432 31952
rect 7380 31909 7389 31943
rect 7389 31909 7423 31943
rect 7423 31909 7432 31943
rect 7380 31900 7432 31909
rect 2872 31764 2924 31816
rect 3148 31764 3200 31816
rect 6644 31764 6696 31816
rect 7656 31900 7708 31952
rect 8116 31900 8168 31952
rect 9956 31900 10008 31952
rect 11152 31900 11204 31952
rect 11796 31943 11848 31952
rect 11796 31909 11805 31943
rect 11805 31909 11839 31943
rect 11839 31909 11848 31943
rect 11796 31900 11848 31909
rect 11888 31943 11940 31952
rect 11888 31909 11897 31943
rect 11897 31909 11931 31943
rect 11931 31909 11940 31943
rect 11888 31900 11940 31909
rect 8024 31832 8076 31884
rect 8852 31832 8904 31884
rect 10048 31832 10100 31884
rect 12440 31832 12492 31884
rect 9864 31764 9916 31816
rect 10232 31807 10284 31816
rect 10232 31773 10241 31807
rect 10241 31773 10275 31807
rect 10275 31773 10284 31807
rect 10232 31764 10284 31773
rect 9680 31696 9732 31748
rect 12164 31696 12216 31748
rect 8760 31628 8812 31680
rect 9312 31628 9364 31680
rect 9772 31671 9824 31680
rect 9772 31637 9781 31671
rect 9781 31637 9815 31671
rect 9815 31637 9824 31671
rect 9772 31628 9824 31637
rect 12624 31628 12676 31680
rect 12900 31671 12952 31680
rect 12900 31637 12909 31671
rect 12909 31637 12943 31671
rect 12943 31637 12952 31671
rect 12900 31628 12952 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 6644 31467 6696 31476
rect 6644 31433 6653 31467
rect 6653 31433 6687 31467
rect 6687 31433 6696 31467
rect 6644 31424 6696 31433
rect 7196 31424 7248 31476
rect 10048 31424 10100 31476
rect 10324 31424 10376 31476
rect 10508 31424 10560 31476
rect 12624 31424 12676 31476
rect 7380 31399 7432 31408
rect 7380 31365 7389 31399
rect 7389 31365 7423 31399
rect 7423 31365 7432 31399
rect 7380 31356 7432 31365
rect 8024 31356 8076 31408
rect 9956 31356 10008 31408
rect 12532 31399 12584 31408
rect 12532 31365 12541 31399
rect 12541 31365 12575 31399
rect 12575 31365 12584 31399
rect 12532 31356 12584 31365
rect 10048 31288 10100 31340
rect 11888 31288 11940 31340
rect 12348 31288 12400 31340
rect 10784 31220 10836 31272
rect 10876 31220 10928 31272
rect 11060 31220 11112 31272
rect 11244 31220 11296 31272
rect 11336 31220 11388 31272
rect 11796 31263 11848 31272
rect 11796 31229 11805 31263
rect 11805 31229 11839 31263
rect 11839 31229 11848 31263
rect 11796 31220 11848 31229
rect 12440 31220 12492 31272
rect 9312 31084 9364 31136
rect 9864 31084 9916 31136
rect 12900 31152 12952 31204
rect 11244 31084 11296 31136
rect 12164 31127 12216 31136
rect 12164 31093 12173 31127
rect 12173 31093 12207 31127
rect 12207 31093 12216 31127
rect 12164 31084 12216 31093
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 9956 30923 10008 30932
rect 9956 30889 9965 30923
rect 9965 30889 9999 30923
rect 9999 30889 10008 30923
rect 9956 30880 10008 30889
rect 10232 30923 10284 30932
rect 10232 30889 10241 30923
rect 10241 30889 10275 30923
rect 10275 30889 10284 30923
rect 10232 30880 10284 30889
rect 12440 30923 12492 30932
rect 12440 30889 12449 30923
rect 12449 30889 12483 30923
rect 12483 30889 12492 30923
rect 12440 30880 12492 30889
rect 1676 30855 1728 30864
rect 1676 30821 1685 30855
rect 1685 30821 1719 30855
rect 1719 30821 1728 30855
rect 1676 30812 1728 30821
rect 10784 30855 10836 30864
rect 10784 30821 10793 30855
rect 10793 30821 10827 30855
rect 10827 30821 10836 30855
rect 10784 30812 10836 30821
rect 11244 30812 11296 30864
rect 12348 30744 12400 30796
rect 1676 30676 1728 30728
rect 7380 30540 7432 30592
rect 9312 30583 9364 30592
rect 9312 30549 9321 30583
rect 9321 30549 9355 30583
rect 9355 30549 9364 30583
rect 9312 30540 9364 30549
rect 11244 30540 11296 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 1676 30379 1728 30388
rect 1676 30345 1685 30379
rect 1685 30345 1719 30379
rect 1719 30345 1728 30379
rect 1676 30336 1728 30345
rect 9312 30336 9364 30388
rect 7012 30268 7064 30320
rect 10140 30200 10192 30252
rect 10416 30200 10468 30252
rect 12164 30200 12216 30252
rect 4252 30132 4304 30184
rect 8208 30132 8260 30184
rect 7196 30107 7248 30116
rect 7196 30073 7205 30107
rect 7205 30073 7239 30107
rect 7239 30073 7248 30107
rect 7196 30064 7248 30073
rect 7380 30107 7432 30116
rect 7380 30073 7389 30107
rect 7389 30073 7423 30107
rect 7423 30073 7432 30107
rect 7380 30064 7432 30073
rect 9772 30064 9824 30116
rect 10140 30107 10192 30116
rect 10140 30073 10149 30107
rect 10149 30073 10183 30107
rect 10183 30073 10192 30107
rect 10140 30064 10192 30073
rect 11244 30132 11296 30184
rect 3424 29996 3476 30048
rect 4436 29996 4488 30048
rect 12164 30064 12216 30116
rect 12348 29996 12400 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 12624 29792 12676 29844
rect 5632 29724 5684 29776
rect 6092 29724 6144 29776
rect 6644 29724 6696 29776
rect 8116 29724 8168 29776
rect 10600 29767 10652 29776
rect 10600 29733 10609 29767
rect 10609 29733 10643 29767
rect 10643 29733 10652 29767
rect 10600 29724 10652 29733
rect 10876 29724 10928 29776
rect 4252 29656 4304 29708
rect 6276 29656 6328 29708
rect 7288 29656 7340 29708
rect 11980 29656 12032 29708
rect 12256 29656 12308 29708
rect 10876 29631 10928 29640
rect 7196 29520 7248 29572
rect 3424 29495 3476 29504
rect 3424 29461 3433 29495
rect 3433 29461 3467 29495
rect 3467 29461 3476 29495
rect 3424 29452 3476 29461
rect 5816 29452 5868 29504
rect 7288 29452 7340 29504
rect 7472 29495 7524 29504
rect 7472 29461 7481 29495
rect 7481 29461 7515 29495
rect 7515 29461 7524 29495
rect 10876 29597 10885 29631
rect 10885 29597 10919 29631
rect 10919 29597 10928 29631
rect 10876 29588 10928 29597
rect 12348 29588 12400 29640
rect 10048 29520 10100 29572
rect 7472 29452 7524 29461
rect 8484 29452 8536 29504
rect 10140 29452 10192 29504
rect 10692 29452 10744 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 7380 29248 7432 29300
rect 10232 29248 10284 29300
rect 10876 29248 10928 29300
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 10140 29180 10192 29232
rect 10784 29180 10836 29232
rect 4252 29155 4304 29164
rect 4252 29121 4261 29155
rect 4261 29121 4295 29155
rect 4295 29121 4304 29155
rect 4252 29112 4304 29121
rect 7564 29112 7616 29164
rect 9956 29112 10008 29164
rect 4436 28976 4488 29028
rect 4620 28976 4672 29028
rect 4988 28976 5040 29028
rect 5540 28976 5592 29028
rect 6000 28976 6052 29028
rect 6276 29019 6328 29028
rect 6276 28985 6285 29019
rect 6285 28985 6319 29019
rect 6319 28985 6328 29019
rect 6276 28976 6328 28985
rect 5632 28951 5684 28960
rect 5632 28917 5641 28951
rect 5641 28917 5675 28951
rect 5675 28917 5684 28951
rect 5632 28908 5684 28917
rect 7288 28976 7340 29028
rect 7748 28976 7800 29028
rect 8116 28976 8168 29028
rect 7104 28908 7156 28960
rect 7380 28951 7432 28960
rect 7380 28917 7389 28951
rect 7389 28917 7423 28951
rect 7423 28917 7432 28951
rect 7380 28908 7432 28917
rect 7840 28908 7892 28960
rect 8484 28976 8536 29028
rect 11980 28976 12032 29028
rect 11060 28908 11112 28960
rect 12348 28908 12400 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 7380 28704 7432 28756
rect 8300 28704 8352 28756
rect 10232 28747 10284 28756
rect 10232 28713 10241 28747
rect 10241 28713 10275 28747
rect 10275 28713 10284 28747
rect 10232 28704 10284 28713
rect 12348 28747 12400 28756
rect 12348 28713 12357 28747
rect 12357 28713 12391 28747
rect 12391 28713 12400 28747
rect 12348 28704 12400 28713
rect 1676 28679 1728 28688
rect 1676 28645 1685 28679
rect 1685 28645 1719 28679
rect 1719 28645 1728 28679
rect 1676 28636 1728 28645
rect 4068 28636 4120 28688
rect 4528 28636 4580 28688
rect 4804 28636 4856 28688
rect 5172 28636 5224 28688
rect 11244 28679 11296 28688
rect 11244 28645 11256 28679
rect 11256 28645 11296 28679
rect 11244 28636 11296 28645
rect 4436 28568 4488 28620
rect 1676 28500 1728 28552
rect 4528 28500 4580 28552
rect 5080 28500 5132 28552
rect 7748 28568 7800 28620
rect 11060 28568 11112 28620
rect 5908 28500 5960 28552
rect 7104 28543 7156 28552
rect 7104 28509 7113 28543
rect 7113 28509 7147 28543
rect 7147 28509 7156 28543
rect 7104 28500 7156 28509
rect 5448 28364 5500 28416
rect 5632 28364 5684 28416
rect 7840 28364 7892 28416
rect 9864 28364 9916 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 5908 28203 5960 28212
rect 5908 28169 5917 28203
rect 5917 28169 5951 28203
rect 5951 28169 5960 28203
rect 5908 28160 5960 28169
rect 7840 28160 7892 28212
rect 4896 28092 4948 28144
rect 7472 28024 7524 28076
rect 10232 28160 10284 28212
rect 10416 28203 10468 28212
rect 10416 28169 10425 28203
rect 10425 28169 10459 28203
rect 10459 28169 10468 28203
rect 10416 28160 10468 28169
rect 10692 28203 10744 28212
rect 10692 28169 10701 28203
rect 10701 28169 10735 28203
rect 10735 28169 10744 28203
rect 10692 28160 10744 28169
rect 10784 28160 10836 28212
rect 11060 28160 11112 28212
rect 11244 28067 11296 28076
rect 11244 28033 11253 28067
rect 11253 28033 11287 28067
rect 11287 28033 11296 28067
rect 11244 28024 11296 28033
rect 2504 27888 2556 27940
rect 5264 27931 5316 27940
rect 5264 27897 5273 27931
rect 5273 27897 5307 27931
rect 5307 27897 5316 27931
rect 5264 27888 5316 27897
rect 5448 27931 5500 27940
rect 5448 27897 5457 27931
rect 5457 27897 5491 27931
rect 5491 27897 5500 27931
rect 5448 27888 5500 27897
rect 5632 27888 5684 27940
rect 8300 27888 8352 27940
rect 9864 27888 9916 27940
rect 1676 27863 1728 27872
rect 1676 27829 1685 27863
rect 1685 27829 1719 27863
rect 1719 27829 1728 27863
rect 1676 27820 1728 27829
rect 2412 27820 2464 27872
rect 2780 27820 2832 27872
rect 3424 27820 3476 27872
rect 5172 27820 5224 27872
rect 8484 27820 8536 27872
rect 10416 27820 10468 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4160 27548 4212 27600
rect 6736 27548 6788 27600
rect 6920 27548 6972 27600
rect 8208 27591 8260 27600
rect 8208 27557 8217 27591
rect 8217 27557 8251 27591
rect 8251 27557 8260 27591
rect 8208 27548 8260 27557
rect 5356 27523 5408 27532
rect 5356 27489 5365 27523
rect 5365 27489 5399 27523
rect 5399 27489 5408 27523
rect 5356 27480 5408 27489
rect 8300 27480 8352 27532
rect 10140 27548 10192 27600
rect 10416 27616 10468 27668
rect 11244 27616 11296 27668
rect 5632 27455 5684 27464
rect 5632 27421 5641 27455
rect 5641 27421 5675 27455
rect 5675 27421 5684 27455
rect 5632 27412 5684 27421
rect 7012 27455 7064 27464
rect 7012 27421 7021 27455
rect 7021 27421 7055 27455
rect 7055 27421 7064 27455
rect 7012 27412 7064 27421
rect 7196 27455 7248 27464
rect 7196 27421 7205 27455
rect 7205 27421 7239 27455
rect 7239 27421 7248 27455
rect 7196 27412 7248 27421
rect 8484 27412 8536 27464
rect 5540 27344 5592 27396
rect 9772 27387 9824 27396
rect 9772 27353 9781 27387
rect 9781 27353 9815 27387
rect 9815 27353 9824 27387
rect 9772 27344 9824 27353
rect 10232 27412 10284 27464
rect 2504 27319 2556 27328
rect 2504 27285 2513 27319
rect 2513 27285 2547 27319
rect 2547 27285 2556 27319
rect 2504 27276 2556 27285
rect 4528 27276 4580 27328
rect 5080 27319 5132 27328
rect 5080 27285 5089 27319
rect 5089 27285 5123 27319
rect 5123 27285 5132 27319
rect 5080 27276 5132 27285
rect 7748 27276 7800 27328
rect 10048 27276 10100 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 4160 27072 4212 27124
rect 7196 27072 7248 27124
rect 10232 27072 10284 27124
rect 10416 27115 10468 27124
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 4620 27047 4672 27056
rect 4620 27013 4629 27047
rect 4629 27013 4663 27047
rect 4663 27013 4672 27047
rect 4620 27004 4672 27013
rect 6920 27047 6972 27056
rect 6920 27013 6929 27047
rect 6929 27013 6963 27047
rect 6963 27013 6972 27047
rect 6920 27004 6972 27013
rect 10048 27047 10100 27056
rect 10048 27013 10057 27047
rect 10057 27013 10091 27047
rect 10091 27013 10100 27047
rect 10048 27004 10100 27013
rect 5080 26979 5132 26988
rect 5080 26945 5089 26979
rect 5089 26945 5123 26979
rect 5123 26945 5132 26979
rect 5080 26936 5132 26945
rect 6644 26936 6696 26988
rect 7012 26936 7064 26988
rect 7104 26936 7156 26988
rect 5264 26868 5316 26920
rect 5816 26868 5868 26920
rect 11336 26868 11388 26920
rect 11520 26868 11572 26920
rect 13820 26868 13872 26920
rect 15752 26868 15804 26920
rect 4896 26800 4948 26852
rect 7012 26800 7064 26852
rect 8208 26800 8260 26852
rect 5356 26732 5408 26784
rect 5540 26775 5592 26784
rect 5540 26741 5549 26775
rect 5549 26741 5583 26775
rect 5583 26741 5592 26775
rect 5540 26732 5592 26741
rect 7380 26775 7432 26784
rect 7380 26741 7389 26775
rect 7389 26741 7423 26775
rect 7423 26741 7432 26775
rect 7380 26732 7432 26741
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 6920 26528 6972 26580
rect 4620 26460 4672 26512
rect 4988 26460 5040 26512
rect 7564 26503 7616 26512
rect 7564 26469 7573 26503
rect 7573 26469 7607 26503
rect 7607 26469 7616 26503
rect 7564 26460 7616 26469
rect 9312 26460 9364 26512
rect 7012 26392 7064 26444
rect 9680 26392 9732 26444
rect 4804 26367 4856 26376
rect 4804 26333 4813 26367
rect 4813 26333 4847 26367
rect 4847 26333 4856 26367
rect 4804 26324 4856 26333
rect 4896 26367 4948 26376
rect 4896 26333 4905 26367
rect 4905 26333 4939 26367
rect 4939 26333 4948 26367
rect 7472 26367 7524 26376
rect 4896 26324 4948 26333
rect 7472 26333 7481 26367
rect 7481 26333 7515 26367
rect 7515 26333 7524 26367
rect 7472 26324 7524 26333
rect 7748 26324 7800 26376
rect 10140 26367 10192 26376
rect 10140 26333 10149 26367
rect 10149 26333 10183 26367
rect 10183 26333 10192 26367
rect 10140 26324 10192 26333
rect 4344 26299 4396 26308
rect 4344 26265 4353 26299
rect 4353 26265 4387 26299
rect 4387 26265 4396 26299
rect 4344 26256 4396 26265
rect 5632 26256 5684 26308
rect 6092 26256 6144 26308
rect 7104 26299 7156 26308
rect 7104 26265 7113 26299
rect 7113 26265 7147 26299
rect 7147 26265 7156 26299
rect 7104 26256 7156 26265
rect 9496 26256 9548 26308
rect 3056 26188 3108 26240
rect 7840 26188 7892 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 2228 26027 2280 26036
rect 2228 25993 2237 26027
rect 2237 25993 2271 26027
rect 2271 25993 2280 26027
rect 2228 25984 2280 25993
rect 2504 25984 2556 26036
rect 3332 25984 3384 26036
rect 4988 26027 5040 26036
rect 4988 25993 4997 26027
rect 4997 25993 5031 26027
rect 5031 25993 5040 26027
rect 4988 25984 5040 25993
rect 7380 26027 7432 26036
rect 7380 25993 7389 26027
rect 7389 25993 7423 26027
rect 7423 25993 7432 26027
rect 7380 25984 7432 25993
rect 4896 25916 4948 25968
rect 6736 25916 6788 25968
rect 7472 25916 7524 25968
rect 9128 25916 9180 25968
rect 9956 25959 10008 25968
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 7932 25848 7984 25900
rect 9956 25925 9965 25959
rect 9965 25925 9999 25959
rect 9999 25925 10008 25959
rect 9956 25916 10008 25925
rect 10600 25848 10652 25900
rect 2228 25780 2280 25832
rect 2412 25780 2464 25832
rect 9312 25780 9364 25832
rect 9680 25780 9732 25832
rect 3056 25712 3108 25764
rect 7840 25755 7892 25764
rect 2596 25687 2648 25696
rect 2596 25653 2605 25687
rect 2605 25653 2639 25687
rect 2639 25653 2648 25687
rect 2596 25644 2648 25653
rect 4804 25644 4856 25696
rect 7840 25721 7849 25755
rect 7849 25721 7883 25755
rect 7883 25721 7892 25755
rect 7840 25712 7892 25721
rect 7748 25644 7800 25696
rect 11060 25712 11112 25764
rect 8484 25644 8536 25696
rect 8576 25644 8628 25696
rect 9220 25644 9272 25696
rect 10968 25687 11020 25696
rect 10968 25653 10977 25687
rect 10977 25653 11011 25687
rect 11011 25653 11020 25687
rect 10968 25644 11020 25653
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 2964 25483 3016 25492
rect 2964 25449 2973 25483
rect 2973 25449 3007 25483
rect 3007 25449 3016 25483
rect 2964 25440 3016 25449
rect 5264 25440 5316 25492
rect 8024 25483 8076 25492
rect 8024 25449 8033 25483
rect 8033 25449 8067 25483
rect 8067 25449 8076 25483
rect 8024 25440 8076 25449
rect 4160 25372 4212 25424
rect 4896 25372 4948 25424
rect 5632 25372 5684 25424
rect 9404 25372 9456 25424
rect 10140 25440 10192 25492
rect 4712 25347 4764 25356
rect 4712 25313 4721 25347
rect 4721 25313 4755 25347
rect 4755 25313 4764 25347
rect 4712 25304 4764 25313
rect 6644 25304 6696 25356
rect 10784 25347 10836 25356
rect 10784 25313 10793 25347
rect 10793 25313 10827 25347
rect 10827 25313 10836 25347
rect 10784 25304 10836 25313
rect 11060 25347 11112 25356
rect 11060 25313 11094 25347
rect 11094 25313 11112 25347
rect 11060 25304 11112 25313
rect 2964 25279 3016 25288
rect 2964 25245 2973 25279
rect 2973 25245 3007 25279
rect 3007 25245 3016 25279
rect 2964 25236 3016 25245
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 4620 25279 4672 25288
rect 3056 25236 3108 25245
rect 4620 25245 4629 25279
rect 4629 25245 4663 25279
rect 4663 25245 4672 25279
rect 4620 25236 4672 25245
rect 2780 25168 2832 25220
rect 3056 25100 3108 25152
rect 3240 25100 3292 25152
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 11060 25100 11112 25152
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 13084 25100 13136 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 2872 24896 2924 24948
rect 4252 24896 4304 24948
rect 4620 24896 4672 24948
rect 5632 24939 5684 24948
rect 5632 24905 5641 24939
rect 5641 24905 5675 24939
rect 5675 24905 5684 24939
rect 5632 24896 5684 24905
rect 7196 24896 7248 24948
rect 7840 24896 7892 24948
rect 10784 24939 10836 24948
rect 10784 24905 10793 24939
rect 10793 24905 10827 24939
rect 10827 24905 10836 24939
rect 10784 24896 10836 24905
rect 11152 24896 11204 24948
rect 12532 24939 12584 24948
rect 12532 24905 12541 24939
rect 12541 24905 12575 24939
rect 12575 24905 12584 24939
rect 12532 24896 12584 24905
rect 2320 24760 2372 24812
rect 3332 24803 3384 24812
rect 3332 24769 3341 24803
rect 3341 24769 3375 24803
rect 3375 24769 3384 24803
rect 3332 24760 3384 24769
rect 1584 24692 1636 24744
rect 2780 24692 2832 24744
rect 3148 24692 3200 24744
rect 4160 24692 4212 24744
rect 1676 24667 1728 24676
rect 1676 24633 1685 24667
rect 1685 24633 1719 24667
rect 1719 24633 1728 24667
rect 1676 24624 1728 24633
rect 3240 24667 3292 24676
rect 3240 24633 3249 24667
rect 3249 24633 3283 24667
rect 3283 24633 3292 24667
rect 3240 24624 3292 24633
rect 5264 24692 5316 24744
rect 4344 24624 4396 24676
rect 4620 24624 4672 24676
rect 6644 24828 6696 24880
rect 7564 24760 7616 24812
rect 12072 24760 12124 24812
rect 8300 24735 8352 24744
rect 8300 24701 8309 24735
rect 8309 24701 8343 24735
rect 8343 24701 8352 24735
rect 8300 24692 8352 24701
rect 8392 24692 8444 24744
rect 11796 24735 11848 24744
rect 11796 24701 11805 24735
rect 11805 24701 11839 24735
rect 11839 24701 11848 24735
rect 11796 24692 11848 24701
rect 8576 24667 8628 24676
rect 8576 24633 8585 24667
rect 8585 24633 8619 24667
rect 8619 24633 8628 24667
rect 8576 24624 8628 24633
rect 10140 24667 10192 24676
rect 10140 24633 10149 24667
rect 10149 24633 10183 24667
rect 10183 24633 10192 24667
rect 10140 24624 10192 24633
rect 7840 24599 7892 24608
rect 7840 24565 7849 24599
rect 7849 24565 7883 24599
rect 7883 24565 7892 24599
rect 7840 24556 7892 24565
rect 8668 24556 8720 24608
rect 9864 24556 9916 24608
rect 11060 24556 11112 24608
rect 12256 24692 12308 24744
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 12348 24624 12400 24676
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 2964 24395 3016 24404
rect 2964 24361 2973 24395
rect 2973 24361 3007 24395
rect 3007 24361 3016 24395
rect 2964 24352 3016 24361
rect 4620 24395 4672 24404
rect 4620 24361 4629 24395
rect 4629 24361 4663 24395
rect 4663 24361 4672 24395
rect 4620 24352 4672 24361
rect 4712 24352 4764 24404
rect 5724 24352 5776 24404
rect 8484 24395 8536 24404
rect 8484 24361 8493 24395
rect 8493 24361 8527 24395
rect 8527 24361 8536 24395
rect 8484 24352 8536 24361
rect 11060 24352 11112 24404
rect 13084 24352 13136 24404
rect 2504 24327 2556 24336
rect 2504 24293 2513 24327
rect 2513 24293 2547 24327
rect 2547 24293 2556 24327
rect 2504 24284 2556 24293
rect 2688 24284 2740 24336
rect 3332 24327 3384 24336
rect 3332 24293 3341 24327
rect 3341 24293 3375 24327
rect 3375 24293 3384 24327
rect 3332 24284 3384 24293
rect 7196 24284 7248 24336
rect 11796 24284 11848 24336
rect 2320 24259 2372 24268
rect 2320 24225 2329 24259
rect 2329 24225 2363 24259
rect 2363 24225 2372 24259
rect 2320 24216 2372 24225
rect 6644 24216 6696 24268
rect 10232 24216 10284 24268
rect 11152 24259 11204 24268
rect 11152 24225 11161 24259
rect 11161 24225 11195 24259
rect 11195 24225 11204 24259
rect 11152 24216 11204 24225
rect 11980 24216 12032 24268
rect 12256 24216 12308 24268
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 6092 24148 6144 24200
rect 8576 24148 8628 24200
rect 10140 24148 10192 24200
rect 5264 24012 5316 24064
rect 11152 24012 11204 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 2504 23808 2556 23860
rect 4804 23851 4856 23860
rect 4804 23817 4813 23851
rect 4813 23817 4847 23851
rect 4847 23817 4856 23851
rect 4804 23808 4856 23817
rect 5908 23808 5960 23860
rect 6644 23808 6696 23860
rect 7012 23808 7064 23860
rect 7932 23851 7984 23860
rect 7932 23817 7941 23851
rect 7941 23817 7975 23851
rect 7975 23817 7984 23851
rect 7932 23808 7984 23817
rect 11796 23851 11848 23860
rect 11796 23817 11805 23851
rect 11805 23817 11839 23851
rect 11839 23817 11848 23851
rect 11796 23808 11848 23817
rect 2688 23740 2740 23792
rect 6092 23740 6144 23792
rect 7564 23740 7616 23792
rect 10600 23783 10652 23792
rect 10600 23749 10609 23783
rect 10609 23749 10643 23783
rect 10643 23749 10652 23783
rect 10600 23740 10652 23749
rect 10968 23740 11020 23792
rect 12256 23740 12308 23792
rect 2504 23672 2556 23724
rect 5356 23715 5408 23724
rect 5356 23681 5365 23715
rect 5365 23681 5399 23715
rect 5399 23681 5408 23715
rect 5356 23672 5408 23681
rect 7196 23672 7248 23724
rect 8576 23672 8628 23724
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 2688 23604 2740 23656
rect 3332 23604 3384 23656
rect 5724 23604 5776 23656
rect 7932 23604 7984 23656
rect 9404 23604 9456 23656
rect 11152 23647 11204 23656
rect 11152 23613 11161 23647
rect 11161 23613 11195 23647
rect 11195 23613 11204 23647
rect 11152 23604 11204 23613
rect 12348 23604 12400 23656
rect 12808 23647 12860 23656
rect 12808 23613 12817 23647
rect 12817 23613 12851 23647
rect 12851 23613 12860 23647
rect 12808 23604 12860 23613
rect 2412 23536 2464 23588
rect 4068 23536 4120 23588
rect 4528 23536 4580 23588
rect 5080 23579 5132 23588
rect 5080 23545 5089 23579
rect 5089 23545 5123 23579
rect 5123 23545 5132 23579
rect 5080 23536 5132 23545
rect 5264 23579 5316 23588
rect 5264 23545 5273 23579
rect 5273 23545 5307 23579
rect 5307 23545 5316 23579
rect 5264 23536 5316 23545
rect 4988 23468 5040 23520
rect 5908 23536 5960 23588
rect 7564 23468 7616 23520
rect 8116 23468 8168 23520
rect 9404 23468 9456 23520
rect 11060 23536 11112 23588
rect 10600 23468 10652 23520
rect 12532 23468 12584 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 2320 23264 2372 23316
rect 5080 23307 5132 23316
rect 5080 23273 5089 23307
rect 5089 23273 5123 23307
rect 5123 23273 5132 23307
rect 5080 23264 5132 23273
rect 6000 23264 6052 23316
rect 7196 23307 7248 23316
rect 7196 23273 7205 23307
rect 7205 23273 7239 23307
rect 7239 23273 7248 23307
rect 7196 23264 7248 23273
rect 7932 23307 7984 23316
rect 7932 23273 7941 23307
rect 7941 23273 7975 23307
rect 7975 23273 7984 23307
rect 7932 23264 7984 23273
rect 9956 23307 10008 23316
rect 9956 23273 9965 23307
rect 9965 23273 9999 23307
rect 9999 23273 10008 23307
rect 9956 23264 10008 23273
rect 11152 23264 11204 23316
rect 12440 23264 12492 23316
rect 13084 23264 13136 23316
rect 2964 23239 3016 23248
rect 2964 23205 2973 23239
rect 2973 23205 3007 23239
rect 3007 23205 3016 23239
rect 2964 23196 3016 23205
rect 2688 23128 2740 23180
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 3240 23128 3292 23180
rect 6828 23196 6880 23248
rect 8576 23239 8628 23248
rect 8576 23205 8585 23239
rect 8585 23205 8619 23239
rect 8619 23205 8628 23239
rect 8576 23196 8628 23205
rect 11612 23196 11664 23248
rect 12256 23196 12308 23248
rect 5356 23128 5408 23180
rect 8760 23128 8812 23180
rect 9496 23128 9548 23180
rect 10692 23128 10744 23180
rect 12164 23128 12216 23180
rect 3056 23103 3108 23112
rect 3056 23069 3065 23103
rect 3065 23069 3099 23103
rect 3099 23069 3108 23103
rect 3056 23060 3108 23069
rect 5908 23103 5960 23112
rect 5908 23069 5917 23103
rect 5917 23069 5951 23103
rect 5951 23069 5960 23103
rect 5908 23060 5960 23069
rect 6092 23060 6144 23112
rect 7196 23060 7248 23112
rect 9404 23060 9456 23112
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 2504 23035 2556 23044
rect 2504 23001 2513 23035
rect 2513 23001 2547 23035
rect 2547 23001 2556 23035
rect 2504 22992 2556 23001
rect 8484 22992 8536 23044
rect 9312 22992 9364 23044
rect 11980 22992 12032 23044
rect 8116 22967 8168 22976
rect 8116 22933 8125 22967
rect 8125 22933 8159 22967
rect 8159 22933 8168 22967
rect 8116 22924 8168 22933
rect 10600 22967 10652 22976
rect 10600 22933 10609 22967
rect 10609 22933 10643 22967
rect 10643 22933 10652 22967
rect 10600 22924 10652 22933
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2780 22720 2832 22772
rect 2964 22720 3016 22772
rect 5908 22720 5960 22772
rect 6092 22763 6144 22772
rect 6092 22729 6101 22763
rect 6101 22729 6135 22763
rect 6135 22729 6144 22763
rect 6092 22720 6144 22729
rect 7196 22763 7248 22772
rect 7196 22729 7205 22763
rect 7205 22729 7239 22763
rect 7239 22729 7248 22763
rect 7196 22720 7248 22729
rect 7840 22763 7892 22772
rect 7840 22729 7849 22763
rect 7849 22729 7883 22763
rect 7883 22729 7892 22763
rect 7840 22720 7892 22729
rect 8576 22720 8628 22772
rect 9864 22720 9916 22772
rect 10324 22720 10376 22772
rect 10692 22763 10744 22772
rect 10692 22729 10701 22763
rect 10701 22729 10735 22763
rect 10735 22729 10744 22763
rect 10692 22720 10744 22729
rect 11060 22720 11112 22772
rect 5632 22652 5684 22704
rect 6000 22652 6052 22704
rect 9680 22695 9732 22704
rect 9680 22661 9689 22695
rect 9689 22661 9723 22695
rect 9723 22661 9732 22695
rect 9680 22652 9732 22661
rect 11612 22584 11664 22636
rect 6920 22516 6972 22568
rect 8300 22516 8352 22568
rect 9956 22559 10008 22568
rect 9956 22525 9965 22559
rect 9965 22525 9999 22559
rect 9999 22525 10008 22559
rect 9956 22516 10008 22525
rect 8484 22448 8536 22500
rect 10140 22491 10192 22500
rect 10140 22457 10149 22491
rect 10149 22457 10183 22491
rect 10183 22457 10192 22491
rect 10140 22448 10192 22457
rect 10784 22448 10836 22500
rect 11060 22448 11112 22500
rect 3056 22380 3108 22432
rect 7840 22380 7892 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 4068 22176 4120 22228
rect 4620 22219 4672 22228
rect 4620 22185 4629 22219
rect 4629 22185 4663 22219
rect 4663 22185 4672 22219
rect 4620 22176 4672 22185
rect 8024 22176 8076 22228
rect 8484 22176 8536 22228
rect 8760 22176 8812 22228
rect 10140 22176 10192 22228
rect 10600 22176 10652 22228
rect 2780 22108 2832 22160
rect 6184 22151 6236 22160
rect 1492 22040 1544 22092
rect 2136 22040 2188 22092
rect 3148 22040 3200 22092
rect 6184 22117 6193 22151
rect 6193 22117 6227 22151
rect 6227 22117 6236 22151
rect 6184 22108 6236 22117
rect 7288 22108 7340 22160
rect 10232 22108 10284 22160
rect 10692 22108 10744 22160
rect 11152 22151 11204 22160
rect 11152 22117 11164 22151
rect 11164 22117 11204 22151
rect 11152 22108 11204 22117
rect 7564 22083 7616 22092
rect 3056 22015 3108 22024
rect 3056 21981 3065 22015
rect 3065 21981 3099 22015
rect 3099 21981 3108 22015
rect 3056 21972 3108 21981
rect 2412 21904 2464 21956
rect 7564 22049 7573 22083
rect 7573 22049 7607 22083
rect 7607 22049 7616 22083
rect 7564 22040 7616 22049
rect 10968 22040 11020 22092
rect 4712 22015 4764 22024
rect 4712 21981 4721 22015
rect 4721 21981 4755 22015
rect 4755 21981 4764 22015
rect 4712 21972 4764 21981
rect 6092 22015 6144 22024
rect 6092 21981 6101 22015
rect 6101 21981 6135 22015
rect 6135 21981 6144 22015
rect 6092 21972 6144 21981
rect 6276 22015 6328 22024
rect 6276 21981 6285 22015
rect 6285 21981 6319 22015
rect 6319 21981 6328 22015
rect 6276 21972 6328 21981
rect 7012 21972 7064 22024
rect 7380 21972 7432 22024
rect 7840 22015 7892 22024
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 5540 21904 5592 21956
rect 4712 21836 4764 21888
rect 5724 21879 5776 21888
rect 5724 21845 5733 21879
rect 5733 21845 5767 21879
rect 5767 21845 5776 21879
rect 5724 21836 5776 21845
rect 7012 21836 7064 21888
rect 10324 21836 10376 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 3056 21632 3108 21684
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 6644 21675 6696 21684
rect 6644 21641 6653 21675
rect 6653 21641 6687 21675
rect 6687 21641 6696 21675
rect 6644 21632 6696 21641
rect 7840 21632 7892 21684
rect 10968 21675 11020 21684
rect 10968 21641 10977 21675
rect 10977 21641 11011 21675
rect 11011 21641 11020 21675
rect 10968 21632 11020 21641
rect 11152 21632 11204 21684
rect 2412 21564 2464 21616
rect 3148 21564 3200 21616
rect 5908 21607 5960 21616
rect 5908 21573 5917 21607
rect 5917 21573 5951 21607
rect 5951 21573 5960 21607
rect 5908 21564 5960 21573
rect 6276 21564 6328 21616
rect 7748 21564 7800 21616
rect 9772 21607 9824 21616
rect 9772 21573 9781 21607
rect 9781 21573 9815 21607
rect 9815 21573 9824 21607
rect 9772 21564 9824 21573
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5172 21496 5224 21548
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 6828 21496 6880 21548
rect 7656 21496 7708 21548
rect 8024 21496 8076 21548
rect 4712 21428 4764 21480
rect 7104 21428 7156 21480
rect 8300 21360 8352 21412
rect 2412 21335 2464 21344
rect 2412 21301 2421 21335
rect 2421 21301 2455 21335
rect 2455 21301 2464 21335
rect 2412 21292 2464 21301
rect 3148 21292 3200 21344
rect 4068 21292 4120 21344
rect 7288 21335 7340 21344
rect 7288 21301 7297 21335
rect 7297 21301 7331 21335
rect 7331 21301 7340 21335
rect 7288 21292 7340 21301
rect 7564 21335 7616 21344
rect 7564 21301 7573 21335
rect 7573 21301 7607 21335
rect 7607 21301 7616 21335
rect 7564 21292 7616 21301
rect 10600 21496 10652 21548
rect 10324 21471 10376 21480
rect 10324 21437 10333 21471
rect 10333 21437 10367 21471
rect 10367 21437 10376 21471
rect 10324 21428 10376 21437
rect 8760 21403 8812 21412
rect 8760 21369 8769 21403
rect 8769 21369 8803 21403
rect 8803 21369 8812 21403
rect 8760 21360 8812 21369
rect 9680 21360 9732 21412
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 2688 21088 2740 21140
rect 4712 21088 4764 21140
rect 7288 21088 7340 21140
rect 7656 21088 7708 21140
rect 1676 21063 1728 21072
rect 1676 21029 1685 21063
rect 1685 21029 1719 21063
rect 1719 21029 1728 21063
rect 1676 21020 1728 21029
rect 7472 21020 7524 21072
rect 10324 21020 10376 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 4344 20995 4396 21004
rect 4344 20961 4378 20995
rect 4378 20961 4396 20995
rect 4344 20952 4396 20961
rect 6092 20952 6144 21004
rect 6920 20952 6972 21004
rect 10968 20952 11020 21004
rect 3516 20884 3568 20936
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 5540 20884 5592 20936
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 6184 20816 6236 20868
rect 6000 20791 6052 20800
rect 6000 20757 6009 20791
rect 6009 20757 6043 20791
rect 6043 20757 6052 20791
rect 6000 20748 6052 20757
rect 8300 20748 8352 20800
rect 8484 20748 8536 20800
rect 8760 20748 8812 20800
rect 9404 20748 9456 20800
rect 11060 20791 11112 20800
rect 11060 20757 11069 20791
rect 11069 20757 11103 20791
rect 11103 20757 11112 20791
rect 11060 20748 11112 20757
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 5540 20544 5592 20596
rect 7380 20544 7432 20596
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 4068 20408 4120 20460
rect 4620 20408 4672 20460
rect 4712 20408 4764 20460
rect 7012 20476 7064 20528
rect 7564 20408 7616 20460
rect 10324 20544 10376 20596
rect 10600 20476 10652 20528
rect 10968 20476 11020 20528
rect 1676 20315 1728 20324
rect 1676 20281 1685 20315
rect 1685 20281 1719 20315
rect 1719 20281 1728 20315
rect 1676 20272 1728 20281
rect 3884 20272 3936 20324
rect 4068 20272 4120 20324
rect 5448 20272 5500 20324
rect 6000 20340 6052 20392
rect 8484 20383 8536 20392
rect 4620 20247 4672 20256
rect 4620 20213 4629 20247
rect 4629 20213 4663 20247
rect 4663 20213 4672 20247
rect 4620 20204 4672 20213
rect 5264 20204 5316 20256
rect 7104 20272 7156 20324
rect 8484 20349 8518 20383
rect 8518 20349 8536 20383
rect 8484 20340 8536 20349
rect 6828 20204 6880 20256
rect 7472 20204 7524 20256
rect 9588 20247 9640 20256
rect 9588 20213 9597 20247
rect 9597 20213 9631 20247
rect 9631 20213 9640 20247
rect 9588 20204 9640 20213
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 1400 20000 1452 20052
rect 3976 20000 4028 20052
rect 4344 20043 4396 20052
rect 4344 20009 4353 20043
rect 4353 20009 4387 20043
rect 4387 20009 4396 20043
rect 4344 20000 4396 20009
rect 5908 20000 5960 20052
rect 6644 20000 6696 20052
rect 7012 20000 7064 20052
rect 9404 20043 9456 20052
rect 4712 19975 4764 19984
rect 4712 19941 4721 19975
rect 4721 19941 4755 19975
rect 4755 19941 4764 19975
rect 4712 19932 4764 19941
rect 5264 19932 5316 19984
rect 5448 19932 5500 19984
rect 7840 19975 7892 19984
rect 7840 19941 7849 19975
rect 7849 19941 7883 19975
rect 7883 19941 7892 19975
rect 7840 19932 7892 19941
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 11980 20000 12032 20052
rect 10600 19864 10652 19916
rect 10968 19907 11020 19916
rect 10968 19873 11002 19907
rect 11002 19873 11020 19907
rect 10968 19864 11020 19873
rect 4712 19796 4764 19848
rect 7932 19796 7984 19848
rect 7104 19728 7156 19780
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 6644 19499 6696 19508
rect 6644 19465 6653 19499
rect 6653 19465 6687 19499
rect 6687 19465 6696 19499
rect 6644 19456 6696 19465
rect 7932 19456 7984 19508
rect 10600 19456 10652 19508
rect 10784 19456 10836 19508
rect 4988 19320 5040 19372
rect 5816 19320 5868 19372
rect 1952 19252 2004 19304
rect 3516 19252 3568 19304
rect 4712 19252 4764 19304
rect 5540 19252 5592 19304
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 7380 19252 7432 19304
rect 7840 19252 7892 19304
rect 9864 19252 9916 19304
rect 2596 19227 2648 19236
rect 2596 19193 2630 19227
rect 2630 19193 2648 19227
rect 2596 19184 2648 19193
rect 7012 19184 7064 19236
rect 9588 19184 9640 19236
rect 9680 19227 9732 19236
rect 9680 19193 9689 19227
rect 9689 19193 9723 19227
rect 9723 19193 9732 19227
rect 9680 19184 9732 19193
rect 3976 19116 4028 19168
rect 6920 19116 6972 19168
rect 10048 19116 10100 19168
rect 10508 19116 10560 19168
rect 10968 19116 11020 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 7840 18912 7892 18964
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 9220 18912 9272 18964
rect 9680 18912 9732 18964
rect 7748 18887 7800 18896
rect 7748 18853 7757 18887
rect 7757 18853 7791 18887
rect 7791 18853 7800 18887
rect 7748 18844 7800 18853
rect 7932 18887 7984 18896
rect 7932 18853 7941 18887
rect 7941 18853 7975 18887
rect 7975 18853 7984 18887
rect 7932 18844 7984 18853
rect 10232 18887 10284 18896
rect 10232 18853 10241 18887
rect 10241 18853 10275 18887
rect 10275 18853 10284 18887
rect 10232 18844 10284 18853
rect 7012 18776 7064 18828
rect 2964 18708 3016 18760
rect 10324 18751 10376 18760
rect 7472 18683 7524 18692
rect 7472 18649 7481 18683
rect 7481 18649 7515 18683
rect 7515 18649 7524 18683
rect 7472 18640 7524 18649
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 11152 18640 11204 18692
rect 2596 18572 2648 18624
rect 9680 18572 9732 18624
rect 10600 18572 10652 18624
rect 10968 18572 11020 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 7748 18368 7800 18420
rect 10232 18368 10284 18420
rect 10968 18368 11020 18420
rect 11152 18368 11204 18420
rect 5172 18300 5224 18352
rect 7012 18300 7064 18352
rect 7472 18300 7524 18352
rect 7932 18300 7984 18352
rect 8760 18300 8812 18352
rect 9312 18300 9364 18352
rect 4804 18232 4856 18284
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 8484 18232 8536 18284
rect 9312 18164 9364 18216
rect 1952 18096 2004 18148
rect 5080 18096 5132 18148
rect 2596 18028 2648 18080
rect 8484 18096 8536 18148
rect 10140 18096 10192 18148
rect 9496 18028 9548 18080
rect 10416 18071 10468 18080
rect 10416 18037 10425 18071
rect 10425 18037 10459 18071
rect 10459 18037 10468 18071
rect 10416 18028 10468 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 5724 17824 5776 17876
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 9772 17824 9824 17876
rect 10416 17824 10468 17876
rect 10600 17824 10652 17876
rect 2872 17756 2924 17808
rect 5448 17799 5500 17808
rect 5448 17765 5457 17799
rect 5457 17765 5491 17799
rect 5491 17765 5500 17799
rect 8576 17799 8628 17808
rect 5448 17756 5500 17765
rect 8576 17765 8585 17799
rect 8585 17765 8619 17799
rect 8619 17765 8628 17799
rect 8576 17756 8628 17765
rect 1952 17688 2004 17740
rect 5080 17688 5132 17740
rect 7380 17688 7432 17740
rect 9588 17688 9640 17740
rect 9864 17688 9916 17740
rect 10324 17731 10376 17740
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 12164 17688 12216 17740
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 8668 17663 8720 17672
rect 3056 17620 3108 17629
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 2228 17552 2280 17604
rect 2596 17552 2648 17604
rect 10784 17552 10836 17604
rect 1952 17484 2004 17536
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 4988 17484 5040 17536
rect 6920 17484 6972 17536
rect 9772 17484 9824 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 1952 17280 2004 17332
rect 2964 17280 3016 17332
rect 3516 17323 3568 17332
rect 3516 17289 3525 17323
rect 3525 17289 3559 17323
rect 3559 17289 3568 17323
rect 3516 17280 3568 17289
rect 5448 17280 5500 17332
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 8576 17280 8628 17332
rect 10968 17280 11020 17332
rect 2044 17144 2096 17196
rect 2596 17144 2648 17196
rect 8668 17212 8720 17264
rect 7196 17144 7248 17196
rect 8208 17144 8260 17196
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 2504 17119 2556 17128
rect 2504 17085 2513 17119
rect 2513 17085 2547 17119
rect 2547 17085 2556 17119
rect 2504 17076 2556 17085
rect 3976 17119 4028 17128
rect 3976 17085 4010 17119
rect 4010 17085 4028 17119
rect 3976 17076 4028 17085
rect 2228 17008 2280 17060
rect 2964 17008 3016 17060
rect 5356 17008 5408 17060
rect 9404 17008 9456 17060
rect 9772 17051 9824 17060
rect 9772 17017 9781 17051
rect 9781 17017 9815 17051
rect 9815 17017 9824 17051
rect 9772 17008 9824 17017
rect 10784 17008 10836 17060
rect 11428 17051 11480 17060
rect 11428 17017 11437 17051
rect 11437 17017 11471 17051
rect 11471 17017 11480 17051
rect 11428 17008 11480 17017
rect 2688 16983 2740 16992
rect 2688 16949 2697 16983
rect 2697 16949 2731 16983
rect 2731 16949 2740 16983
rect 2688 16940 2740 16949
rect 2872 16940 2924 16992
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 2688 16736 2740 16788
rect 2136 16668 2188 16720
rect 3976 16736 4028 16788
rect 4344 16736 4396 16788
rect 5448 16779 5500 16788
rect 4620 16711 4672 16720
rect 2044 16600 2096 16652
rect 2320 16532 2372 16584
rect 4620 16677 4629 16711
rect 4629 16677 4663 16711
rect 4663 16677 4672 16711
rect 4620 16668 4672 16677
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 5080 16711 5132 16720
rect 5080 16677 5089 16711
rect 5089 16677 5123 16711
rect 5123 16677 5132 16711
rect 5080 16668 5132 16677
rect 6000 16668 6052 16720
rect 2596 16600 2648 16652
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 5540 16600 5592 16652
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 3424 16532 3476 16584
rect 9956 16532 10008 16584
rect 11428 16600 11480 16652
rect 10784 16575 10836 16584
rect 10784 16541 10793 16575
rect 10793 16541 10827 16575
rect 10827 16541 10836 16575
rect 10784 16532 10836 16541
rect 1768 16396 1820 16448
rect 3056 16396 3108 16448
rect 3516 16396 3568 16448
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 5264 16396 5316 16448
rect 7656 16439 7708 16448
rect 7656 16405 7665 16439
rect 7665 16405 7699 16439
rect 7699 16405 7708 16439
rect 7656 16396 7708 16405
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 2320 16192 2372 16244
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 2780 16192 2832 16244
rect 4252 16192 4304 16244
rect 4620 16192 4672 16244
rect 5540 16192 5592 16244
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 9404 16235 9456 16244
rect 9404 16201 9413 16235
rect 9413 16201 9447 16235
rect 9447 16201 9456 16235
rect 9404 16192 9456 16201
rect 11428 16192 11480 16244
rect 4804 16124 4856 16176
rect 7380 16167 7432 16176
rect 7380 16133 7389 16167
rect 7389 16133 7423 16167
rect 7423 16133 7432 16167
rect 7380 16124 7432 16133
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 4068 16056 4120 16108
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 7840 16099 7892 16108
rect 7840 16065 7849 16099
rect 7849 16065 7883 16099
rect 7883 16065 7892 16099
rect 7840 16056 7892 16065
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 4988 16031 5040 16040
rect 4988 15997 4997 16031
rect 4997 15997 5031 16031
rect 5031 15997 5040 16031
rect 4988 15988 5040 15997
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 8484 15988 8536 16040
rect 3516 15920 3568 15972
rect 5172 15963 5224 15972
rect 5172 15929 5181 15963
rect 5181 15929 5215 15963
rect 5215 15929 5224 15963
rect 5172 15920 5224 15929
rect 7656 15920 7708 15972
rect 10048 15920 10100 15972
rect 10232 15920 10284 15972
rect 3608 15895 3660 15904
rect 3608 15861 3617 15895
rect 3617 15861 3651 15895
rect 3651 15861 3660 15895
rect 3608 15852 3660 15861
rect 4436 15895 4488 15904
rect 4436 15861 4445 15895
rect 4445 15861 4479 15895
rect 4479 15861 4488 15895
rect 4436 15852 4488 15861
rect 8300 15852 8352 15904
rect 9404 15852 9456 15904
rect 10784 15852 10836 15904
rect 11060 15852 11112 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 4344 15691 4396 15700
rect 4344 15657 4353 15691
rect 4353 15657 4387 15691
rect 4387 15657 4396 15691
rect 4344 15648 4396 15657
rect 5172 15648 5224 15700
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 1584 15580 1636 15632
rect 3608 15580 3660 15632
rect 5264 15580 5316 15632
rect 10416 15580 10468 15632
rect 6920 15512 6972 15564
rect 8208 15512 8260 15564
rect 9956 15512 10008 15564
rect 11520 15555 11572 15564
rect 11520 15521 11554 15555
rect 11554 15521 11572 15555
rect 11520 15512 11572 15521
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 5540 15444 5592 15496
rect 5908 15444 5960 15496
rect 7012 15444 7064 15496
rect 9680 15444 9732 15496
rect 10048 15444 10100 15496
rect 11060 15444 11112 15496
rect 2136 15419 2188 15428
rect 2136 15385 2145 15419
rect 2145 15385 2179 15419
rect 2179 15385 2188 15419
rect 2136 15376 2188 15385
rect 9772 15419 9824 15428
rect 9772 15385 9781 15419
rect 9781 15385 9815 15419
rect 9815 15385 9824 15419
rect 9772 15376 9824 15385
rect 9404 15351 9456 15360
rect 9404 15317 9413 15351
rect 9413 15317 9447 15351
rect 9447 15317 9456 15351
rect 9404 15308 9456 15317
rect 12440 15308 12492 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 2228 15104 2280 15156
rect 2688 15104 2740 15156
rect 6828 15104 6880 15156
rect 7012 15104 7064 15156
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 9956 15104 10008 15156
rect 11520 15104 11572 15156
rect 2504 15036 2556 15088
rect 2780 15036 2832 15088
rect 4988 15036 5040 15088
rect 3424 15011 3476 15020
rect 3424 14977 3433 15011
rect 3433 14977 3467 15011
rect 3467 14977 3476 15011
rect 3424 14968 3476 14977
rect 5356 15036 5408 15088
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 3148 14900 3200 14952
rect 3516 14943 3568 14952
rect 3516 14909 3525 14943
rect 3525 14909 3559 14943
rect 3559 14909 3568 14943
rect 3516 14900 3568 14909
rect 4160 14900 4212 14952
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 6828 14832 6880 14884
rect 1584 14764 1636 14816
rect 3424 14807 3476 14816
rect 3424 14773 3433 14807
rect 3433 14773 3467 14807
rect 3467 14773 3476 14807
rect 3424 14764 3476 14773
rect 5816 14764 5868 14816
rect 6184 14764 6236 14816
rect 8208 14832 8260 14884
rect 8484 14832 8536 14884
rect 8760 14764 8812 14816
rect 10048 14764 10100 14816
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 11060 14764 11112 14816
rect 11520 14764 11572 14816
rect 12624 14764 12676 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 1400 14560 1452 14612
rect 2780 14560 2832 14612
rect 5632 14560 5684 14612
rect 6184 14560 6236 14612
rect 7380 14560 7432 14612
rect 8300 14560 8352 14612
rect 8852 14560 8904 14612
rect 12624 14560 12676 14612
rect 1492 14492 1544 14544
rect 3240 14535 3292 14544
rect 3240 14501 3249 14535
rect 3249 14501 3283 14535
rect 3283 14501 3292 14535
rect 3240 14492 3292 14501
rect 4804 14492 4856 14544
rect 5264 14492 5316 14544
rect 5540 14492 5592 14544
rect 8024 14492 8076 14544
rect 8576 14492 8628 14544
rect 8668 14492 8720 14544
rect 9680 14492 9732 14544
rect 10140 14492 10192 14544
rect 12348 14535 12400 14544
rect 12348 14501 12382 14535
rect 12382 14501 12400 14535
rect 12348 14492 12400 14501
rect 11060 14424 11112 14476
rect 12072 14467 12124 14476
rect 12072 14433 12081 14467
rect 12081 14433 12115 14467
rect 12115 14433 12124 14467
rect 12072 14424 12124 14433
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 5724 14288 5776 14340
rect 7656 14288 7708 14340
rect 10416 14288 10468 14340
rect 3148 14220 3200 14272
rect 4620 14263 4672 14272
rect 4620 14229 4629 14263
rect 4629 14229 4663 14263
rect 4663 14229 4672 14263
rect 4620 14220 4672 14229
rect 7472 14220 7524 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 3424 14016 3476 14068
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 8668 14016 8720 14068
rect 8760 14016 8812 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10140 14016 10192 14068
rect 11428 14016 11480 14068
rect 12348 14016 12400 14068
rect 5264 13991 5316 14000
rect 5264 13957 5273 13991
rect 5273 13957 5307 13991
rect 5307 13957 5316 13991
rect 5264 13948 5316 13957
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 2780 13880 2832 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 7012 13991 7064 14000
rect 7012 13957 7021 13991
rect 7021 13957 7055 13991
rect 7055 13957 7064 13991
rect 7012 13948 7064 13957
rect 12072 13948 12124 14000
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 7472 13880 7524 13932
rect 8300 13880 8352 13932
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 3240 13812 3292 13864
rect 3516 13812 3568 13864
rect 5172 13812 5224 13864
rect 2688 13744 2740 13796
rect 3056 13744 3108 13796
rect 3792 13787 3844 13796
rect 3792 13753 3801 13787
rect 3801 13753 3835 13787
rect 3835 13753 3844 13787
rect 3792 13744 3844 13753
rect 6184 13812 6236 13864
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 6092 13744 6144 13796
rect 6920 13744 6972 13796
rect 8024 13812 8076 13864
rect 8484 13812 8536 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 10324 13744 10376 13796
rect 2780 13719 2832 13728
rect 2780 13685 2789 13719
rect 2789 13685 2823 13719
rect 2823 13685 2832 13719
rect 2780 13676 2832 13685
rect 3240 13676 3292 13728
rect 5356 13676 5408 13728
rect 7104 13676 7156 13728
rect 7380 13676 7432 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 4804 13472 4856 13524
rect 4988 13515 5040 13524
rect 4988 13481 4997 13515
rect 4997 13481 5031 13515
rect 5031 13481 5040 13515
rect 4988 13472 5040 13481
rect 6920 13472 6972 13524
rect 10324 13515 10376 13524
rect 10324 13481 10333 13515
rect 10333 13481 10367 13515
rect 10367 13481 10376 13515
rect 10324 13472 10376 13481
rect 2228 13404 2280 13456
rect 2688 13404 2740 13456
rect 5540 13404 5592 13456
rect 5908 13404 5960 13456
rect 11520 13404 11572 13456
rect 12348 13404 12400 13456
rect 3056 13268 3108 13320
rect 2688 13200 2740 13252
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 2044 13132 2096 13184
rect 5356 13175 5408 13184
rect 5356 13141 5365 13175
rect 5365 13141 5399 13175
rect 5399 13141 5408 13175
rect 5356 13132 5408 13141
rect 6092 13132 6144 13184
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 5356 12928 5408 12980
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 10324 12928 10376 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 3056 12860 3108 12912
rect 5540 12860 5592 12912
rect 2688 12792 2740 12844
rect 6000 12860 6052 12912
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 3056 12724 3108 12733
rect 5448 12724 5500 12776
rect 5908 12724 5960 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 2136 12699 2188 12708
rect 2136 12665 2145 12699
rect 2145 12665 2179 12699
rect 2179 12665 2188 12699
rect 2136 12656 2188 12665
rect 3148 12656 3200 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 2228 12588 2280 12640
rect 9864 12724 9916 12776
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 8300 12656 8352 12708
rect 7012 12588 7064 12640
rect 7288 12588 7340 12640
rect 8208 12588 8260 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 1860 12384 1912 12436
rect 3056 12384 3108 12436
rect 5448 12384 5500 12436
rect 7012 12384 7064 12436
rect 8300 12384 8352 12436
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 2136 12316 2188 12368
rect 2412 12316 2464 12368
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 2780 12112 2832 12164
rect 4620 12316 4672 12368
rect 4988 12359 5040 12368
rect 4988 12325 4997 12359
rect 4997 12325 5031 12359
rect 5031 12325 5040 12359
rect 4988 12316 5040 12325
rect 7472 12316 7524 12368
rect 10048 12316 10100 12368
rect 4620 12180 4672 12232
rect 5264 12248 5316 12300
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 9956 12248 10008 12300
rect 4896 12180 4948 12232
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 7932 12180 7984 12189
rect 9404 12180 9456 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10600 12180 10652 12232
rect 11520 12180 11572 12232
rect 12624 12180 12676 12232
rect 7380 12155 7432 12164
rect 7380 12121 7389 12155
rect 7389 12121 7423 12155
rect 7423 12121 7432 12155
rect 7380 12112 7432 12121
rect 4528 12087 4580 12096
rect 4528 12053 4537 12087
rect 4537 12053 4571 12087
rect 4571 12053 4580 12087
rect 4528 12044 4580 12053
rect 10692 12044 10744 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 2872 11840 2924 11892
rect 4896 11883 4948 11892
rect 4896 11849 4905 11883
rect 4905 11849 4939 11883
rect 4939 11849 4948 11883
rect 4896 11840 4948 11849
rect 4988 11840 5040 11892
rect 7656 11840 7708 11892
rect 8208 11840 8260 11892
rect 8576 11840 8628 11892
rect 11060 11772 11112 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 9680 11704 9732 11756
rect 10140 11704 10192 11756
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 3056 11636 3108 11688
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 3332 11568 3384 11620
rect 7932 11568 7984 11620
rect 9680 11568 9732 11620
rect 10232 11568 10284 11620
rect 10600 11568 10652 11620
rect 2780 11500 2832 11552
rect 7472 11500 7524 11552
rect 10048 11500 10100 11552
rect 10876 11543 10928 11552
rect 10876 11509 10885 11543
rect 10885 11509 10919 11543
rect 10919 11509 10928 11543
rect 10876 11500 10928 11509
rect 12808 11500 12860 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 1400 11296 1452 11348
rect 2872 11296 2924 11348
rect 3056 11339 3108 11348
rect 3056 11305 3065 11339
rect 3065 11305 3099 11339
rect 3099 11305 3108 11339
rect 3056 11296 3108 11305
rect 4620 11296 4672 11348
rect 4896 11296 4948 11348
rect 6644 11296 6696 11348
rect 7564 11296 7616 11348
rect 7840 11296 7892 11348
rect 8392 11296 8444 11348
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 6092 11228 6144 11280
rect 10968 11271 11020 11280
rect 10968 11237 10977 11271
rect 10977 11237 11011 11271
rect 11011 11237 11020 11271
rect 10968 11228 11020 11237
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 10140 11160 10192 11212
rect 10600 11160 10652 11212
rect 13084 11296 13136 11348
rect 12348 11228 12400 11280
rect 12624 11271 12676 11280
rect 12624 11237 12633 11271
rect 12633 11237 12667 11271
rect 12667 11237 12676 11271
rect 12624 11228 12676 11237
rect 3332 11067 3384 11076
rect 3332 11033 3341 11067
rect 3341 11033 3375 11067
rect 3375 11033 3384 11067
rect 3332 11024 3384 11033
rect 7656 11024 7708 11076
rect 8484 11092 8536 11144
rect 10324 11092 10376 11144
rect 12716 11160 12768 11212
rect 12900 11160 12952 11212
rect 12624 11092 12676 11144
rect 7380 10956 7432 11008
rect 11244 10956 11296 11008
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 13084 10956 13136 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 6092 10795 6144 10804
rect 6092 10761 6101 10795
rect 6101 10761 6135 10795
rect 6135 10761 6144 10795
rect 6092 10752 6144 10761
rect 8484 10752 8536 10804
rect 10968 10752 11020 10804
rect 12348 10752 12400 10804
rect 10140 10727 10192 10736
rect 10140 10693 10149 10727
rect 10149 10693 10183 10727
rect 10183 10693 10192 10727
rect 10140 10684 10192 10693
rect 10324 10684 10376 10736
rect 11152 10684 11204 10736
rect 13360 10684 13412 10736
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 12440 10616 12492 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 4252 10548 4304 10600
rect 4528 10548 4580 10600
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 8116 10480 8168 10532
rect 11060 10480 11112 10532
rect 4988 10412 5040 10464
rect 6920 10412 6972 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 12716 10412 12768 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 1768 10208 1820 10260
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 8484 10208 8536 10260
rect 9772 10208 9824 10260
rect 11336 10208 11388 10260
rect 4252 10140 4304 10192
rect 6644 10183 6696 10192
rect 6644 10149 6678 10183
rect 6678 10149 6696 10183
rect 6644 10140 6696 10149
rect 11060 10140 11112 10192
rect 11796 10140 11848 10192
rect 12164 10140 12216 10192
rect 13084 10140 13136 10192
rect 13360 10183 13412 10192
rect 13360 10149 13369 10183
rect 13369 10149 13403 10183
rect 13403 10149 13412 10183
rect 13360 10140 13412 10149
rect 13544 10183 13596 10192
rect 13544 10149 13553 10183
rect 13553 10149 13587 10183
rect 13587 10149 13596 10183
rect 13544 10140 13596 10149
rect 4344 10072 4396 10124
rect 5540 10072 5592 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 9956 10072 10008 10124
rect 10600 10072 10652 10124
rect 12440 10072 12492 10124
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 10232 10004 10284 10056
rect 11336 10004 11388 10056
rect 4068 9936 4120 9988
rect 10876 9936 10928 9988
rect 12532 9936 12584 9988
rect 3148 9868 3200 9920
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 5172 9911 5224 9920
rect 5172 9877 5181 9911
rect 5181 9877 5215 9911
rect 5215 9877 5224 9911
rect 5172 9868 5224 9877
rect 8116 9868 8168 9920
rect 11520 9911 11572 9920
rect 11520 9877 11529 9911
rect 11529 9877 11563 9911
rect 11563 9877 11572 9911
rect 11520 9868 11572 9877
rect 12716 9868 12768 9920
rect 12808 9911 12860 9920
rect 12808 9877 12817 9911
rect 12817 9877 12851 9911
rect 12851 9877 12860 9911
rect 12808 9868 12860 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 3240 9664 3292 9716
rect 6644 9664 6696 9716
rect 8484 9707 8536 9716
rect 8484 9673 8493 9707
rect 8493 9673 8527 9707
rect 8527 9673 8536 9707
rect 8484 9664 8536 9673
rect 9772 9664 9824 9716
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 11336 9664 11388 9716
rect 11520 9664 11572 9716
rect 13544 9664 13596 9716
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 3792 9596 3844 9648
rect 6368 9639 6420 9648
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 7472 9639 7524 9648
rect 7472 9605 7481 9639
rect 7481 9605 7515 9639
rect 7515 9605 7524 9639
rect 7472 9596 7524 9605
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 3516 9571 3568 9580
rect 1768 9460 1820 9512
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 3976 9528 4028 9580
rect 4068 9528 4120 9580
rect 5080 9528 5132 9580
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 12164 9639 12216 9648
rect 12164 9605 12173 9639
rect 12173 9605 12207 9639
rect 12207 9605 12216 9639
rect 12164 9596 12216 9605
rect 12256 9596 12308 9648
rect 12440 9596 12492 9648
rect 3056 9460 3108 9512
rect 2872 9392 2924 9444
rect 3240 9435 3292 9444
rect 3240 9401 3249 9435
rect 3249 9401 3283 9435
rect 3283 9401 3292 9435
rect 3240 9392 3292 9401
rect 4988 9435 5040 9444
rect 4988 9401 4997 9435
rect 4997 9401 5031 9435
rect 5031 9401 5040 9435
rect 4988 9392 5040 9401
rect 5172 9392 5224 9444
rect 2044 9324 2096 9376
rect 3056 9324 3108 9376
rect 3148 9324 3200 9376
rect 4344 9324 4396 9376
rect 4712 9324 4764 9376
rect 5816 9324 5868 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7840 9392 7892 9444
rect 10140 9460 10192 9512
rect 13544 9367 13596 9376
rect 7196 9324 7248 9333
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 2780 9120 2832 9172
rect 4068 9120 4120 9172
rect 5172 9120 5224 9172
rect 6920 9163 6972 9172
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 11152 9120 11204 9172
rect 13452 9120 13504 9172
rect 3056 9095 3108 9104
rect 2596 8984 2648 9036
rect 2780 8984 2832 9036
rect 3056 9061 3065 9095
rect 3065 9061 3099 9095
rect 3099 9061 3108 9095
rect 3056 9052 3108 9061
rect 3516 9052 3568 9104
rect 4712 9052 4764 9104
rect 7932 9052 7984 9104
rect 10600 9052 10652 9104
rect 12348 9052 12400 9104
rect 13176 9095 13228 9104
rect 13176 9061 13185 9095
rect 13185 9061 13219 9095
rect 13219 9061 13228 9095
rect 13176 9052 13228 9061
rect 4068 8984 4120 9036
rect 4344 8984 4396 9036
rect 5540 8984 5592 9036
rect 9864 8984 9916 9036
rect 11428 8984 11480 9036
rect 12256 8984 12308 9036
rect 12900 9027 12952 9036
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 8116 8959 8168 8968
rect 2688 8848 2740 8900
rect 3148 8848 3200 8900
rect 3608 8848 3660 8900
rect 4068 8848 4120 8900
rect 7840 8848 7892 8900
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 12900 8993 12932 9027
rect 12932 8993 12952 9027
rect 12900 8984 12952 8993
rect 8208 8848 8260 8900
rect 2780 8780 2832 8832
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 3516 8576 3568 8628
rect 4988 8576 5040 8628
rect 7012 8576 7064 8628
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 6000 8508 6052 8560
rect 6276 8508 6328 8560
rect 8852 8508 8904 8560
rect 11520 8508 11572 8560
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 2044 8372 2096 8424
rect 6920 8372 6972 8424
rect 8208 8372 8260 8424
rect 6368 8304 6420 8356
rect 7380 8347 7432 8356
rect 7380 8313 7389 8347
rect 7389 8313 7423 8347
rect 7423 8313 7432 8347
rect 7380 8304 7432 8313
rect 11612 8372 11664 8424
rect 11980 8372 12032 8424
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 9496 8347 9548 8356
rect 9496 8313 9505 8347
rect 9505 8313 9539 8347
rect 9539 8313 9548 8347
rect 9496 8304 9548 8313
rect 1952 8236 2004 8288
rect 2688 8236 2740 8288
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 6092 8236 6144 8288
rect 9588 8236 9640 8288
rect 10324 8236 10376 8288
rect 10600 8279 10652 8288
rect 10600 8245 10609 8279
rect 10609 8245 10643 8279
rect 10643 8245 10652 8279
rect 10600 8236 10652 8245
rect 12348 8236 12400 8288
rect 13268 8279 13320 8288
rect 13268 8245 13277 8279
rect 13277 8245 13311 8279
rect 13311 8245 13320 8279
rect 13268 8236 13320 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 2596 8032 2648 8084
rect 2780 8032 2832 8084
rect 2044 7964 2096 8016
rect 2688 7828 2740 7880
rect 3976 8032 4028 8084
rect 4804 8032 4856 8084
rect 4988 8032 5040 8084
rect 5816 8032 5868 8084
rect 8116 8032 8168 8084
rect 5448 7964 5500 8016
rect 8392 8007 8444 8016
rect 8392 7973 8401 8007
rect 8401 7973 8435 8007
rect 8435 7973 8444 8007
rect 8392 7964 8444 7973
rect 8576 8007 8628 8016
rect 8576 7973 8585 8007
rect 8585 7973 8619 8007
rect 8619 7973 8628 8007
rect 8576 7964 8628 7973
rect 9496 8032 9548 8084
rect 11428 8075 11480 8084
rect 9864 7964 9916 8016
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 10508 7964 10560 8016
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 12348 7896 12400 7948
rect 4344 7828 4396 7880
rect 11796 7871 11848 7880
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 4804 7692 4856 7744
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 10600 7760 10652 7812
rect 5264 7692 5316 7744
rect 8300 7692 8352 7744
rect 9588 7692 9640 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 2688 7488 2740 7540
rect 2780 7488 2832 7540
rect 4252 7488 4304 7540
rect 8576 7488 8628 7540
rect 8392 7420 8444 7472
rect 9864 7420 9916 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 2504 7284 2556 7336
rect 5448 7284 5500 7336
rect 204 7216 256 7268
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 5264 7191 5316 7200
rect 2780 7148 2832 7157
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 7380 7284 7432 7336
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 10692 7284 10744 7336
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 6920 7216 6972 7268
rect 9588 7216 9640 7268
rect 11428 7216 11480 7268
rect 5264 7148 5316 7157
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8208 7148 8260 7157
rect 10324 7148 10376 7200
rect 12348 7148 12400 7200
rect 14188 7148 14240 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 5448 6987 5500 6996
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 7564 6944 7616 6996
rect 10048 6944 10100 6996
rect 2504 6876 2556 6928
rect 1676 6808 1728 6860
rect 1860 6808 1912 6860
rect 2780 6808 2832 6860
rect 10508 6876 10560 6928
rect 4344 6851 4396 6860
rect 4344 6817 4378 6851
rect 4378 6817 4396 6851
rect 4344 6808 4396 6817
rect 7656 6808 7708 6860
rect 8300 6808 8352 6860
rect 9312 6808 9364 6860
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 1492 6740 1544 6792
rect 4068 6783 4120 6792
rect 2780 6672 2832 6724
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 9864 6740 9916 6792
rect 10232 6740 10284 6792
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 2412 6604 2464 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 11244 6604 11296 6656
rect 13728 6604 13780 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2136 6400 2188 6452
rect 2320 6400 2372 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 10508 6400 10560 6452
rect 9036 6375 9088 6384
rect 9036 6341 9045 6375
rect 9045 6341 9079 6375
rect 9079 6341 9088 6375
rect 9036 6332 9088 6341
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 2228 6239 2280 6248
rect 1952 6196 2004 6205
rect 2228 6205 2262 6239
rect 2262 6205 2280 6239
rect 2228 6196 2280 6205
rect 4068 6196 4120 6248
rect 4252 6196 4304 6248
rect 6920 6196 6972 6248
rect 8392 6196 8444 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 12624 6400 12676 6452
rect 12808 6400 12860 6452
rect 2688 6060 2740 6112
rect 4344 6128 4396 6180
rect 8852 6128 8904 6180
rect 9956 6128 10008 6180
rect 10416 6128 10468 6180
rect 4252 6060 4304 6112
rect 5264 6060 5316 6112
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 7656 6060 7708 6112
rect 8760 6060 8812 6112
rect 10232 6060 10284 6112
rect 12072 6060 12124 6112
rect 12992 6060 13044 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 2228 5856 2280 5908
rect 3424 5856 3476 5908
rect 8852 5856 8904 5908
rect 9036 5856 9088 5908
rect 9864 5856 9916 5908
rect 12624 5856 12676 5908
rect 7380 5788 7432 5840
rect 8300 5831 8352 5840
rect 8300 5797 8309 5831
rect 8309 5797 8343 5831
rect 8343 5797 8352 5831
rect 8300 5788 8352 5797
rect 9772 5788 9824 5840
rect 10324 5831 10376 5840
rect 10324 5797 10333 5831
rect 10333 5797 10367 5831
rect 10367 5797 10376 5831
rect 10324 5788 10376 5797
rect 10508 5788 10560 5840
rect 12164 5788 12216 5840
rect 1952 5720 2004 5772
rect 6828 5720 6880 5772
rect 7932 5720 7984 5772
rect 1768 5652 1820 5704
rect 2688 5652 2740 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 8392 5695 8444 5704
rect 7656 5652 7708 5661
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 11428 5652 11480 5704
rect 1860 5627 1912 5636
rect 1860 5593 1869 5627
rect 1869 5593 1903 5627
rect 1903 5593 1912 5627
rect 1860 5584 1912 5593
rect 2780 5584 2832 5636
rect 10876 5584 10928 5636
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 3240 5516 3292 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 7104 5516 7156 5568
rect 8300 5516 8352 5568
rect 10416 5516 10468 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 6828 5312 6880 5364
rect 7012 5312 7064 5364
rect 4068 5176 4120 5228
rect 7380 5312 7432 5364
rect 9772 5312 9824 5364
rect 12164 5312 12216 5364
rect 7748 5287 7800 5296
rect 7748 5253 7757 5287
rect 7757 5253 7791 5287
rect 7791 5253 7800 5287
rect 7748 5244 7800 5253
rect 9956 5287 10008 5296
rect 9956 5253 9965 5287
rect 9965 5253 9999 5287
rect 9999 5253 10008 5287
rect 9956 5244 10008 5253
rect 2320 5108 2372 5160
rect 7472 5108 7524 5160
rect 3424 5040 3476 5092
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 3148 4972 3200 5024
rect 7196 5040 7248 5092
rect 10600 5176 10652 5228
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 8484 5108 8536 5160
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 8392 5040 8444 5092
rect 10416 5083 10468 5092
rect 10416 5049 10425 5083
rect 10425 5049 10459 5083
rect 10459 5049 10468 5083
rect 10416 5040 10468 5049
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 5448 4972 5500 5024
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 7012 4972 7064 5024
rect 10232 4972 10284 5024
rect 11428 4972 11480 5024
rect 12532 4972 12584 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2320 4768 2372 4820
rect 2688 4811 2740 4820
rect 2688 4777 2697 4811
rect 2697 4777 2731 4811
rect 2731 4777 2740 4811
rect 2688 4768 2740 4777
rect 4068 4768 4120 4820
rect 6644 4768 6696 4820
rect 7748 4768 7800 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 11152 4768 11204 4820
rect 4804 4700 4856 4752
rect 4988 4700 5040 4752
rect 7564 4743 7616 4752
rect 7564 4709 7573 4743
rect 7573 4709 7607 4743
rect 7607 4709 7616 4743
rect 7564 4700 7616 4709
rect 10692 4700 10744 4752
rect 4344 4632 4396 4684
rect 4896 4632 4948 4684
rect 5724 4632 5776 4684
rect 7288 4632 7340 4684
rect 7748 4632 7800 4684
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 9680 4632 9732 4684
rect 11980 4675 12032 4684
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 2228 4539 2280 4548
rect 2228 4505 2237 4539
rect 2237 4505 2271 4539
rect 2271 4505 2280 4539
rect 2228 4496 2280 4505
rect 4160 4539 4212 4548
rect 4160 4505 4169 4539
rect 4169 4505 4203 4539
rect 4203 4505 4212 4539
rect 4160 4496 4212 4505
rect 3424 4428 3476 4480
rect 7380 4564 7432 4616
rect 9404 4564 9456 4616
rect 10600 4564 10652 4616
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 12716 4632 12768 4684
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 11244 4564 11296 4616
rect 6920 4496 6972 4548
rect 8392 4539 8444 4548
rect 8392 4505 8401 4539
rect 8401 4505 8435 4539
rect 8435 4505 8444 4539
rect 8392 4496 8444 4505
rect 9588 4496 9640 4548
rect 10416 4496 10468 4548
rect 5448 4428 5500 4480
rect 7196 4428 7248 4480
rect 8668 4471 8720 4480
rect 8668 4437 8677 4471
rect 8677 4437 8711 4471
rect 8711 4437 8720 4471
rect 8668 4428 8720 4437
rect 9312 4428 9364 4480
rect 11060 4428 11112 4480
rect 12256 4428 12308 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 1952 4224 2004 4276
rect 4344 4267 4396 4276
rect 4344 4233 4353 4267
rect 4353 4233 4387 4267
rect 4387 4233 4396 4267
rect 4344 4224 4396 4233
rect 5724 4224 5776 4276
rect 6828 4224 6880 4276
rect 7104 4224 7156 4276
rect 7564 4224 7616 4276
rect 8484 4224 8536 4276
rect 4160 4088 4212 4140
rect 5172 4088 5224 4140
rect 5264 4088 5316 4140
rect 2412 3952 2464 4004
rect 5080 4020 5132 4072
rect 7380 4156 7432 4208
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 7564 4088 7616 4140
rect 8208 4088 8260 4140
rect 9312 4088 9364 4140
rect 10692 4224 10744 4276
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 13176 4267 13228 4276
rect 13176 4233 13185 4267
rect 13185 4233 13219 4267
rect 13219 4233 13228 4267
rect 13176 4224 13228 4233
rect 11060 4088 11112 4140
rect 11152 4088 11204 4140
rect 7380 4020 7432 4072
rect 9404 4020 9456 4072
rect 6920 3952 6972 4004
rect 8300 3952 8352 4004
rect 8944 3995 8996 4004
rect 8944 3961 8953 3995
rect 8953 3961 8987 3995
rect 8987 3961 8996 3995
rect 8944 3952 8996 3961
rect 9772 4020 9824 4072
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 12624 4020 12676 4072
rect 4344 3884 4396 3936
rect 4804 3884 4856 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 7012 3884 7064 3936
rect 8668 3884 8720 3936
rect 9588 3884 9640 3936
rect 9680 3884 9732 3936
rect 10048 3884 10100 3936
rect 12716 3952 12768 4004
rect 10692 3884 10744 3936
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 7564 3723 7616 3732
rect 2964 3655 3016 3664
rect 2964 3621 2973 3655
rect 2973 3621 3007 3655
rect 3007 3621 3016 3655
rect 2964 3612 3016 3621
rect 5448 3655 5500 3664
rect 5448 3621 5482 3655
rect 5482 3621 5500 3655
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 8852 3680 8904 3732
rect 7104 3655 7156 3664
rect 5448 3612 5500 3621
rect 7104 3621 7113 3655
rect 7113 3621 7147 3655
rect 7147 3621 7156 3655
rect 7104 3612 7156 3621
rect 7472 3612 7524 3664
rect 7932 3612 7984 3664
rect 8944 3612 8996 3664
rect 9404 3655 9456 3664
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 9404 3612 9456 3621
rect 10048 3655 10100 3664
rect 10048 3621 10057 3655
rect 10057 3621 10091 3655
rect 10091 3621 10100 3655
rect 10048 3612 10100 3621
rect 10416 3612 10468 3664
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 3148 3544 3200 3596
rect 3976 3544 4028 3596
rect 1768 3476 1820 3528
rect 2596 3476 2648 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 4344 3544 4396 3596
rect 6276 3544 6328 3596
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 8668 3544 8720 3596
rect 13084 3587 13136 3596
rect 13084 3553 13093 3587
rect 13093 3553 13127 3587
rect 13127 3553 13136 3587
rect 13084 3544 13136 3553
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 13360 3544 13412 3553
rect 2688 3408 2740 3460
rect 2412 3340 2464 3392
rect 4712 3476 4764 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 6920 3408 6972 3460
rect 12808 3451 12860 3460
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 12808 3408 12860 3417
rect 3424 3383 3476 3392
rect 3424 3349 3433 3383
rect 3433 3349 3467 3383
rect 3467 3349 3476 3383
rect 3424 3340 3476 3349
rect 4068 3340 4120 3392
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 2780 3136 2832 3145
rect 3148 3136 3200 3188
rect 5724 3136 5776 3188
rect 8208 3136 8260 3188
rect 9588 3136 9640 3188
rect 10416 3136 10468 3188
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 1400 3068 1452 3120
rect 6276 3111 6328 3120
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 6276 3077 6285 3111
rect 6285 3077 6319 3111
rect 6319 3077 6328 3111
rect 6276 3068 6328 3077
rect 3056 3000 3108 3052
rect 7564 3000 7616 3052
rect 10876 3068 10928 3120
rect 13084 3068 13136 3120
rect 2872 2932 2924 2984
rect 3976 2932 4028 2984
rect 4344 2932 4396 2984
rect 4988 2932 5040 2984
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 2964 2864 3016 2916
rect 3056 2864 3108 2916
rect 3240 2907 3292 2916
rect 3240 2873 3249 2907
rect 3249 2873 3283 2907
rect 3283 2873 3292 2907
rect 3240 2864 3292 2873
rect 3424 2864 3476 2916
rect 7380 2907 7432 2916
rect 7380 2873 7389 2907
rect 7389 2873 7423 2907
rect 7423 2873 7432 2907
rect 7380 2864 7432 2873
rect 2688 2796 2740 2848
rect 5448 2796 5500 2848
rect 13268 3000 13320 3052
rect 8760 2932 8812 2984
rect 9312 2932 9364 2984
rect 11336 2932 11388 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 8852 2864 8904 2916
rect 10232 2796 10284 2848
rect 11520 2796 11572 2848
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 2044 2524 2096 2576
rect 572 2320 624 2372
rect 3056 2524 3108 2576
rect 2688 2320 2740 2372
rect 4068 2524 4120 2576
rect 5448 2524 5500 2576
rect 4252 2456 4304 2508
rect 7840 2456 7892 2508
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 8300 2592 8352 2644
rect 10048 2592 10100 2644
rect 11336 2592 11388 2644
rect 8300 2456 8352 2508
rect 10876 2499 10928 2508
rect 10876 2465 10885 2499
rect 10885 2465 10919 2499
rect 10919 2465 10928 2499
rect 10876 2456 10928 2465
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 7012 2363 7064 2372
rect 7012 2329 7021 2363
rect 7021 2329 7055 2363
rect 7055 2329 7064 2363
rect 7012 2320 7064 2329
rect 8208 2320 8260 2372
rect 10600 2363 10652 2372
rect 10600 2329 10609 2363
rect 10609 2329 10643 2363
rect 10643 2329 10652 2363
rect 10600 2320 10652 2329
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 6644 1368 6696 1420
rect 8944 1368 8996 1420
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1306 39520 1362 40000
rect 1674 39520 1730 40000
rect 2134 39520 2190 40000
rect 2502 39520 2558 40000
rect 2870 39520 2926 40000
rect 3238 39520 3294 40000
rect 3698 39520 3754 40000
rect 4066 39520 4122 40000
rect 4434 39520 4490 40000
rect 4802 39520 4858 40000
rect 5262 39520 5318 40000
rect 5630 39520 5686 40000
rect 5998 39520 6054 40000
rect 6366 39520 6422 40000
rect 6826 39520 6882 40000
rect 7194 39520 7250 40000
rect 7562 39520 7618 40000
rect 7930 39520 7986 40000
rect 8390 39520 8446 40000
rect 8758 39520 8814 40000
rect 9126 39520 9182 40000
rect 9494 39520 9550 40000
rect 9954 39520 10010 40000
rect 10322 39520 10378 40000
rect 10690 39520 10746 40000
rect 11058 39520 11114 40000
rect 11518 39520 11574 40000
rect 11886 39520 11942 40000
rect 12254 39520 12310 40000
rect 12622 39520 12678 40000
rect 13082 39520 13138 40000
rect 13450 39520 13506 40000
rect 13818 39520 13874 40000
rect 14186 39520 14242 40000
rect 14646 39520 14702 40000
rect 15014 39520 15070 40000
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34785 244 39520
rect 202 34776 258 34785
rect 202 34711 258 34720
rect 584 33425 612 39520
rect 570 33416 626 33425
rect 570 33351 626 33360
rect 952 32881 980 39520
rect 938 32872 994 32881
rect 938 32807 994 32816
rect 1320 31385 1348 39520
rect 1582 36408 1638 36417
rect 1582 36343 1638 36352
rect 1596 35698 1624 36343
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1582 34096 1638 34105
rect 1582 34031 1638 34040
rect 1596 32434 1624 34031
rect 1688 33538 1716 39520
rect 1768 35624 1820 35630
rect 1768 35566 1820 35572
rect 1780 34950 1808 35566
rect 1768 34944 1820 34950
rect 1768 34886 1820 34892
rect 1780 33930 1808 34886
rect 2044 34060 2096 34066
rect 2044 34002 2096 34008
rect 1768 33924 1820 33930
rect 1768 33866 1820 33872
rect 1688 33510 1808 33538
rect 1676 33448 1728 33454
rect 1676 33390 1728 33396
rect 1688 33318 1716 33390
rect 1676 33312 1728 33318
rect 1676 33254 1728 33260
rect 1688 33114 1716 33254
rect 1780 33153 1808 33510
rect 1766 33144 1822 33153
rect 1676 33108 1728 33114
rect 1766 33079 1822 33088
rect 1676 33050 1728 33056
rect 2056 32570 2084 34002
rect 2044 32564 2096 32570
rect 2044 32506 2096 32512
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1400 32360 1452 32366
rect 1398 32328 1400 32337
rect 1452 32328 1454 32337
rect 1398 32263 1454 32272
rect 1412 32026 1440 32263
rect 2056 32026 2084 32506
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 2044 32020 2096 32026
rect 2044 31962 2096 31968
rect 2148 31906 2176 39520
rect 2228 35488 2280 35494
rect 2516 35442 2544 39520
rect 2778 38720 2834 38729
rect 2778 38655 2834 38664
rect 2228 35430 2280 35436
rect 2240 35086 2268 35430
rect 2332 35414 2544 35442
rect 2228 35080 2280 35086
rect 2228 35022 2280 35028
rect 2228 34944 2280 34950
rect 2228 34886 2280 34892
rect 2240 34202 2268 34886
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 1412 31878 2176 31906
rect 1306 31376 1362 31385
rect 1306 31311 1362 31320
rect 1412 21298 1440 31878
rect 1674 31648 1730 31657
rect 1674 31583 1730 31592
rect 1688 30870 1716 31583
rect 1676 30864 1728 30870
rect 1676 30806 1728 30812
rect 1688 30734 1716 30765
rect 1676 30728 1728 30734
rect 1674 30696 1676 30705
rect 1728 30696 1730 30705
rect 1674 30631 1730 30640
rect 1688 30394 1716 30631
rect 1676 30388 1728 30394
rect 1676 30330 1728 30336
rect 2332 29628 2360 35414
rect 2504 35216 2556 35222
rect 2504 35158 2556 35164
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 2424 32842 2452 35022
rect 2516 34746 2544 35158
rect 2504 34740 2556 34746
rect 2504 34682 2556 34688
rect 2792 34134 2820 38655
rect 2780 34128 2832 34134
rect 2780 34070 2832 34076
rect 2792 33658 2820 34070
rect 2780 33652 2832 33658
rect 2700 33612 2780 33640
rect 2700 33046 2728 33612
rect 2780 33594 2832 33600
rect 2792 33529 2820 33594
rect 2688 33040 2740 33046
rect 2688 32982 2740 32988
rect 2780 33040 2832 33046
rect 2780 32982 2832 32988
rect 2792 32881 2820 32982
rect 2778 32872 2834 32881
rect 2412 32836 2464 32842
rect 2778 32807 2834 32816
rect 2412 32778 2464 32784
rect 2792 32366 2820 32807
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2884 31822 2912 39520
rect 3252 35714 3280 39520
rect 3712 37210 3740 39520
rect 3068 35686 3280 35714
rect 3344 37182 3740 37210
rect 2964 35080 3016 35086
rect 2964 35022 3016 35028
rect 2976 33998 3004 35022
rect 2964 33992 3016 33998
rect 2964 33934 3016 33940
rect 2976 33386 3004 33934
rect 2964 33380 3016 33386
rect 2964 33322 3016 33328
rect 2976 32230 3004 33322
rect 2964 32224 3016 32230
rect 2964 32166 3016 32172
rect 2976 32026 3004 32166
rect 2964 32020 3016 32026
rect 2964 31962 3016 31968
rect 2872 31816 2924 31822
rect 2872 31758 2924 31764
rect 3068 30161 3096 35686
rect 3240 34944 3292 34950
rect 3240 34886 3292 34892
rect 3252 34746 3280 34886
rect 3240 34740 3292 34746
rect 3240 34682 3292 34688
rect 3146 34640 3202 34649
rect 3146 34575 3148 34584
rect 3200 34575 3202 34584
rect 3148 34546 3200 34552
rect 3252 34406 3280 34682
rect 3240 34400 3292 34406
rect 3240 34342 3292 34348
rect 3238 33008 3294 33017
rect 3148 32972 3200 32978
rect 3238 32943 3294 32952
rect 3148 32914 3200 32920
rect 3160 31958 3188 32914
rect 3252 32910 3280 32943
rect 3240 32904 3292 32910
rect 3240 32846 3292 32852
rect 3252 32502 3280 32846
rect 3240 32496 3292 32502
rect 3240 32438 3292 32444
rect 3148 31952 3200 31958
rect 3148 31894 3200 31900
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 3054 30152 3110 30161
rect 3054 30087 3110 30096
rect 1504 29600 2360 29628
rect 1504 22098 1532 29600
rect 1674 29336 1730 29345
rect 1674 29271 1730 29280
rect 1688 28694 1716 29271
rect 1676 28688 1728 28694
rect 1676 28630 1728 28636
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1688 27878 1716 28494
rect 2504 27940 2556 27946
rect 2504 27882 2556 27888
rect 1676 27872 1728 27878
rect 1674 27840 1676 27849
rect 2412 27872 2464 27878
rect 1728 27840 1730 27849
rect 2412 27814 2464 27820
rect 1674 27775 1730 27784
rect 1582 27024 1638 27033
rect 1582 26959 1638 26968
rect 1596 25906 1624 26959
rect 2226 26344 2282 26353
rect 2226 26279 2282 26288
rect 2240 26042 2268 26279
rect 2228 26036 2280 26042
rect 2228 25978 2280 25984
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 2240 25838 2268 25978
rect 2424 25838 2452 27814
rect 2516 27334 2544 27882
rect 2780 27872 2832 27878
rect 2700 27832 2780 27860
rect 2504 27328 2556 27334
rect 2504 27270 2556 27276
rect 2516 26042 2544 27270
rect 2504 26036 2556 26042
rect 2504 25978 2556 25984
rect 2228 25832 2280 25838
rect 2228 25774 2280 25780
rect 2412 25832 2464 25838
rect 2412 25774 2464 25780
rect 2596 25696 2648 25702
rect 2594 25664 2596 25673
rect 2648 25664 2650 25673
rect 2594 25599 2650 25608
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1596 24410 1624 24686
rect 1676 24676 1728 24682
rect 1676 24618 1728 24624
rect 1688 24585 1716 24618
rect 1674 24576 1730 24585
rect 1674 24511 1730 24520
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 2332 24274 2360 24754
rect 2700 24342 2728 27832
rect 2780 27814 2832 27820
rect 3056 26240 3108 26246
rect 3056 26182 3108 26188
rect 2962 25800 3018 25809
rect 3068 25770 3096 26182
rect 2962 25735 3018 25744
rect 3056 25764 3108 25770
rect 2976 25498 3004 25735
rect 3056 25706 3108 25712
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 2976 25378 3004 25434
rect 2884 25350 3004 25378
rect 2780 25220 2832 25226
rect 2780 25162 2832 25168
rect 2792 24750 2820 25162
rect 2884 24954 2912 25350
rect 3068 25294 3096 25706
rect 2964 25288 3016 25294
rect 2964 25230 3016 25236
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2504 24336 2556 24342
rect 2504 24278 2556 24284
rect 2688 24336 2740 24342
rect 2688 24278 2740 24284
rect 2320 24268 2372 24274
rect 2320 24210 2372 24216
rect 2332 23322 2360 24210
rect 2516 23866 2544 24278
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2700 23798 2728 24278
rect 2688 23792 2740 23798
rect 2688 23734 2740 23740
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2320 23316 2372 23322
rect 2320 23258 2372 23264
rect 1674 22264 1730 22273
rect 1674 22199 1730 22208
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1412 21270 1624 21298
rect 1398 21040 1454 21049
rect 1596 21026 1624 21270
rect 1688 21078 1716 22199
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 1398 20975 1400 20984
rect 1452 20975 1454 20984
rect 1504 20998 1624 21026
rect 1676 21072 1728 21078
rect 1676 21014 1728 21020
rect 1400 20946 1452 20952
rect 1412 20058 1440 20946
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1398 16144 1454 16153
rect 1398 16079 1454 16088
rect 1412 16046 1440 16079
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 14618 1440 15982
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1504 14550 1532 20998
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 1688 19961 1716 20266
rect 1674 19952 1730 19961
rect 1674 19887 1730 19896
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18426 1992 19246
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1964 17746 1992 18090
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 1582 17640 1638 17649
rect 1582 17575 1638 17584
rect 1596 16114 1624 17575
rect 1964 17542 1992 17682
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17338 1992 17478
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16658 2084 17138
rect 2148 16969 2176 22034
rect 2424 21962 2452 23530
rect 2516 23050 2544 23666
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 2700 23186 2728 23598
rect 2688 23180 2740 23186
rect 2688 23122 2740 23128
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2504 23044 2556 23050
rect 2504 22986 2556 22992
rect 2792 22778 2820 23122
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 2412 21956 2464 21962
rect 2412 21898 2464 21904
rect 2412 21616 2464 21622
rect 2412 21558 2464 21564
rect 2424 21350 2452 21558
rect 2412 21344 2464 21350
rect 2412 21286 2464 21292
rect 2226 20496 2282 20505
rect 2226 20431 2228 20440
rect 2280 20431 2282 20440
rect 2228 20402 2280 20408
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2240 17066 2268 17546
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 2134 16960 2190 16969
rect 2134 16895 2190 16904
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1584 15632 1636 15638
rect 1584 15574 1636 15580
rect 1596 14822 1624 15574
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1492 14544 1544 14550
rect 1492 14486 1544 14492
rect 1596 12986 1624 14758
rect 1688 13870 1716 15127
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1398 11792 1454 11801
rect 1596 11762 1624 12815
rect 1398 11727 1454 11736
rect 1584 11756 1636 11762
rect 1412 11694 1440 11727
rect 1584 11698 1636 11704
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11354 1440 11630
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1596 9586 1624 10503
rect 1780 10266 1808 16390
rect 2148 15434 2176 16662
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2240 15162 2268 17002
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2332 16250 2360 16526
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2226 13968 2282 13977
rect 2226 13903 2228 13912
rect 2280 13903 2282 13912
rect 2228 13874 2280 13880
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1872 12442 1900 12650
rect 2056 12646 2084 13126
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 2148 12374 2176 12650
rect 2240 12646 2268 13398
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2136 12368 2188 12374
rect 2136 12310 2188 12316
rect 2240 12186 2268 12582
rect 2424 12374 2452 21286
rect 2792 21162 2820 22102
rect 2700 21146 2820 21162
rect 2688 21140 2820 21146
rect 2740 21134 2820 21140
rect 2688 21082 2740 21088
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2608 18630 2636 19178
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2608 18086 2636 18566
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2608 17610 2636 18022
rect 2884 17814 2912 24890
rect 2976 24410 3004 25230
rect 3068 25158 3096 25230
rect 3056 25152 3108 25158
rect 3056 25094 3108 25100
rect 2964 24404 3016 24410
rect 2964 24346 3016 24352
rect 2964 23248 3016 23254
rect 2964 23190 3016 23196
rect 2976 23089 3004 23190
rect 3068 23118 3096 25094
rect 3160 24750 3188 31758
rect 3344 26194 3372 37182
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3976 35760 4028 35766
rect 3976 35702 4028 35708
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3422 34776 3478 34785
rect 3622 34768 3918 34788
rect 3422 34711 3478 34720
rect 3436 34610 3464 34711
rect 3424 34604 3476 34610
rect 3424 34546 3476 34552
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3516 32836 3568 32842
rect 3516 32778 3568 32784
rect 3528 32298 3556 32778
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3988 32434 4016 35702
rect 3976 32428 4028 32434
rect 3976 32370 4028 32376
rect 3516 32292 3568 32298
rect 3516 32234 3568 32240
rect 3988 32026 4016 32370
rect 3976 32020 4028 32026
rect 3976 31962 4028 31968
rect 4080 31906 4108 39520
rect 4344 36032 4396 36038
rect 4344 35974 4396 35980
rect 4356 34542 4384 35974
rect 4448 35601 4476 39520
rect 4620 36032 4672 36038
rect 4620 35974 4672 35980
rect 4632 35698 4660 35974
rect 4528 35692 4580 35698
rect 4528 35634 4580 35640
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 4434 35592 4490 35601
rect 4434 35527 4490 35536
rect 4540 34610 4568 35634
rect 4816 35494 4844 39520
rect 5276 35714 5304 39520
rect 5540 37732 5592 37738
rect 5540 37674 5592 37680
rect 5184 35686 5304 35714
rect 4804 35488 4856 35494
rect 4804 35430 4856 35436
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 4896 35080 4948 35086
rect 4896 35022 4948 35028
rect 4620 34944 4672 34950
rect 4620 34886 4672 34892
rect 4528 34604 4580 34610
rect 4528 34546 4580 34552
rect 4632 34542 4660 34886
rect 4802 34776 4858 34785
rect 4802 34711 4858 34720
rect 4344 34536 4396 34542
rect 4344 34478 4396 34484
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 4160 34060 4212 34066
rect 4160 34002 4212 34008
rect 4172 33454 4200 34002
rect 4356 33862 4384 34478
rect 4632 34134 4660 34478
rect 4816 34406 4844 34711
rect 4908 34406 4936 35022
rect 4804 34400 4856 34406
rect 4804 34342 4856 34348
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 4620 34128 4672 34134
rect 4620 34070 4672 34076
rect 4344 33856 4396 33862
rect 4344 33798 4396 33804
rect 4356 33454 4384 33798
rect 4632 33640 4660 34070
rect 4632 33612 4752 33640
rect 4160 33448 4212 33454
rect 4160 33390 4212 33396
rect 4344 33448 4396 33454
rect 4344 33390 4396 33396
rect 4356 32978 4384 33390
rect 4618 33144 4674 33153
rect 4724 33114 4752 33612
rect 4618 33079 4620 33088
rect 4672 33079 4674 33088
rect 4712 33108 4764 33114
rect 4620 33050 4672 33056
rect 4712 33050 4764 33056
rect 4344 32972 4396 32978
rect 4344 32914 4396 32920
rect 4632 32570 4660 33050
rect 4344 32564 4396 32570
rect 4344 32506 4396 32512
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4160 32360 4212 32366
rect 4160 32302 4212 32308
rect 3988 31878 4108 31906
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3424 30048 3476 30054
rect 3424 29990 3476 29996
rect 3436 29510 3464 29990
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 3436 27878 3464 29446
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3424 27872 3476 27878
rect 3424 27814 3476 27820
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3344 26166 3464 26194
rect 3332 26036 3384 26042
rect 3332 25978 3384 25984
rect 3240 25152 3292 25158
rect 3240 25094 3292 25100
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3252 24682 3280 25094
rect 3344 24818 3372 25978
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 3240 24676 3292 24682
rect 3240 24618 3292 24624
rect 3344 24342 3372 24754
rect 3436 24721 3464 26166
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3422 24712 3478 24721
rect 3422 24647 3478 24656
rect 3332 24336 3384 24342
rect 3332 24278 3384 24284
rect 3146 23760 3202 23769
rect 3146 23695 3202 23704
rect 3056 23112 3108 23118
rect 2962 23080 3018 23089
rect 3056 23054 3108 23060
rect 2962 23015 3018 23024
rect 2976 22778 3004 23015
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 3068 22438 3096 23054
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 3068 22030 3096 22374
rect 3160 22098 3188 23695
rect 3344 23662 3372 24278
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3068 21690 3096 21966
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 3160 21622 3188 22034
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2516 17134 2544 17478
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2516 16250 2544 17070
rect 2608 16658 2636 17138
rect 2884 16998 2912 17750
rect 2976 17678 3004 18702
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2976 17338 3004 17614
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2700 16794 2728 16934
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2700 16674 2728 16730
rect 2596 16652 2648 16658
rect 2700 16646 2820 16674
rect 2596 16594 2648 16600
rect 2792 16250 2820 16646
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2884 15960 2912 16934
rect 2608 15932 2912 15960
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 15094 2544 15438
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2148 12158 2268 12186
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1780 9518 1808 10202
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9178 2084 9318
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 8430 2084 9114
rect 2148 8537 2176 12158
rect 2502 10568 2558 10577
rect 2502 10503 2558 10512
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 2134 8528 2190 8537
rect 2134 8463 2190 8472
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1582 8120 1638 8129
rect 1582 8055 1638 8064
rect 1596 7410 1624 8055
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 204 7268 256 7274
rect 204 7210 256 7216
rect 216 480 244 7210
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 572 2372 624 2378
rect 572 2314 624 2320
rect 584 480 612 2314
rect 952 480 980 3567
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 1412 480 1440 3062
rect 1504 1193 1532 6734
rect 1688 5574 1716 6802
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 1596 3058 1624 3431
rect 1688 3369 1716 5510
rect 1780 5370 1808 5646
rect 1872 5642 1900 6802
rect 1964 6254 1992 8230
rect 2056 8022 2084 8366
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2148 6610 2176 8463
rect 2332 7449 2360 9415
rect 2516 7970 2544 10503
rect 2608 9761 2636 15932
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2700 15162 2728 15438
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2792 14618 2820 15030
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2700 13462 2728 13738
rect 2792 13734 2820 13874
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2792 13274 2820 13670
rect 2700 13258 2820 13274
rect 2688 13252 2820 13258
rect 2740 13246 2820 13252
rect 2688 13194 2740 13200
rect 2700 12850 2728 13194
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2700 12356 2728 12786
rect 2700 12328 2912 12356
rect 2884 12238 2912 12328
rect 2688 12232 2740 12238
rect 2686 12200 2688 12209
rect 2872 12232 2924 12238
rect 2740 12200 2742 12209
rect 2872 12174 2924 12180
rect 2686 12135 2742 12144
rect 2780 12164 2832 12170
rect 2700 11898 2728 12135
rect 2780 12106 2832 12112
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2792 11558 2820 12106
rect 2884 11898 2912 12174
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2594 9752 2650 9761
rect 2594 9687 2650 9696
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8090 2636 8978
rect 2700 8906 2728 9551
rect 2792 9330 2820 11494
rect 2884 11354 2912 11834
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2976 9738 3004 17002
rect 3068 16454 3096 17614
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3160 16266 3188 21286
rect 3252 19417 3280 23122
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3528 20942 3556 21422
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3882 20360 3938 20369
rect 3882 20295 3884 20304
rect 3936 20295 3938 20304
rect 3988 20346 4016 31878
rect 4068 28688 4120 28694
rect 4068 28630 4120 28636
rect 4080 23594 4108 28630
rect 4172 27606 4200 32302
rect 4252 30184 4304 30190
rect 4252 30126 4304 30132
rect 4264 29714 4292 30126
rect 4252 29708 4304 29714
rect 4252 29650 4304 29656
rect 4264 29170 4292 29650
rect 4252 29164 4304 29170
rect 4252 29106 4304 29112
rect 4160 27600 4212 27606
rect 4160 27542 4212 27548
rect 4172 27130 4200 27542
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4356 26874 4384 32506
rect 4436 30048 4488 30054
rect 4436 29990 4488 29996
rect 4448 29034 4476 29990
rect 4436 29028 4488 29034
rect 4620 29028 4672 29034
rect 4436 28970 4488 28976
rect 4540 28988 4620 29016
rect 4448 28626 4476 28970
rect 4540 28694 4568 28988
rect 4620 28970 4672 28976
rect 4816 28694 4844 34342
rect 4908 34066 4936 34342
rect 4896 34060 4948 34066
rect 4896 34002 4948 34008
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 4908 32502 4936 32846
rect 4896 32496 4948 32502
rect 4894 32464 4896 32473
rect 4948 32464 4950 32473
rect 4894 32399 4950 32408
rect 4908 32373 4936 32399
rect 5000 29034 5028 35430
rect 5080 34672 5132 34678
rect 5080 34614 5132 34620
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 4528 28688 4580 28694
rect 4528 28630 4580 28636
rect 4804 28688 4856 28694
rect 4804 28630 4856 28636
rect 4436 28620 4488 28626
rect 4436 28562 4488 28568
rect 5092 28558 5120 34614
rect 5184 29209 5212 35686
rect 5448 35216 5500 35222
rect 5448 35158 5500 35164
rect 5460 34542 5488 35158
rect 5448 34536 5500 34542
rect 5448 34478 5500 34484
rect 5460 34202 5488 34478
rect 5448 34196 5500 34202
rect 5448 34138 5500 34144
rect 5264 32496 5316 32502
rect 5264 32438 5316 32444
rect 5276 32337 5304 32438
rect 5460 32366 5488 34138
rect 5448 32360 5500 32366
rect 5262 32328 5318 32337
rect 5448 32302 5500 32308
rect 5262 32263 5318 32272
rect 5264 32224 5316 32230
rect 5264 32166 5316 32172
rect 5276 32026 5304 32166
rect 5264 32020 5316 32026
rect 5264 31962 5316 31968
rect 5170 29200 5226 29209
rect 5170 29135 5226 29144
rect 5552 29034 5580 37674
rect 5644 35193 5672 39520
rect 6012 37890 6040 39520
rect 5828 37862 6040 37890
rect 5630 35184 5686 35193
rect 5630 35119 5686 35128
rect 5724 33108 5776 33114
rect 5724 33050 5776 33056
rect 5736 32434 5764 33050
rect 5724 32428 5776 32434
rect 5724 32370 5776 32376
rect 5828 31793 5856 37862
rect 6380 37738 6408 39520
rect 6368 37732 6420 37738
rect 6368 37674 6420 37680
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6736 34672 6788 34678
rect 6642 34640 6698 34649
rect 6736 34614 6788 34620
rect 6642 34575 6698 34584
rect 6092 34400 6144 34406
rect 6092 34342 6144 34348
rect 6104 33998 6132 34342
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6092 33992 6144 33998
rect 6092 33934 6144 33940
rect 6104 33318 6132 33934
rect 6092 33312 6144 33318
rect 6012 33260 6092 33266
rect 6012 33254 6144 33260
rect 6012 33238 6132 33254
rect 6012 32366 6040 33238
rect 6104 33189 6132 33238
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6656 33046 6684 34575
rect 6748 33114 6776 34614
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6644 33040 6696 33046
rect 6644 32982 6696 32988
rect 6184 32972 6236 32978
rect 6184 32914 6236 32920
rect 6092 32768 6144 32774
rect 6092 32710 6144 32716
rect 6000 32360 6052 32366
rect 6000 32302 6052 32308
rect 6012 32042 6040 32302
rect 6104 32230 6132 32710
rect 6092 32224 6144 32230
rect 6092 32166 6144 32172
rect 6012 32014 6132 32042
rect 6196 32026 6224 32914
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6656 32026 6684 32982
rect 6736 32836 6788 32842
rect 6736 32778 6788 32784
rect 6748 32026 6776 32778
rect 5814 31784 5870 31793
rect 5814 31719 5870 31728
rect 5722 30152 5778 30161
rect 5722 30087 5778 30096
rect 5632 29776 5684 29782
rect 5632 29718 5684 29724
rect 5540 29028 5592 29034
rect 5540 28970 5592 28976
rect 5644 28966 5672 29718
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 5172 28688 5224 28694
rect 5172 28630 5224 28636
rect 4528 28552 4580 28558
rect 4528 28494 4580 28500
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 4540 27334 4568 28494
rect 4896 28144 4948 28150
rect 4896 28086 4948 28092
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4540 27033 4568 27270
rect 4620 27056 4672 27062
rect 4526 27024 4582 27033
rect 4620 26998 4672 27004
rect 4526 26959 4582 26968
rect 4356 26846 4476 26874
rect 4342 26344 4398 26353
rect 4342 26279 4344 26288
rect 4396 26279 4398 26288
rect 4344 26250 4396 26256
rect 4342 25664 4398 25673
rect 4342 25599 4398 25608
rect 4160 25424 4212 25430
rect 4160 25366 4212 25372
rect 4172 24750 4200 25366
rect 4252 24948 4304 24954
rect 4252 24890 4304 24896
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4172 23633 4200 24686
rect 4158 23624 4214 23633
rect 4068 23588 4120 23594
rect 4158 23559 4214 23568
rect 4068 23530 4120 23536
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 4080 21350 4108 22170
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4080 20466 4108 20878
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 4264 20346 4292 24890
rect 4356 24682 4384 25599
rect 4344 24676 4396 24682
rect 4344 24618 4396 24624
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 3988 20330 4108 20346
rect 3988 20324 4120 20330
rect 3988 20318 4068 20324
rect 3884 20266 3936 20272
rect 3988 20058 4016 20318
rect 4068 20266 4120 20272
rect 4172 20318 4292 20346
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3988 19417 4016 19994
rect 3238 19408 3294 19417
rect 3238 19343 3294 19352
rect 3974 19408 4030 19417
rect 3974 19343 4030 19352
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 17338 3556 19246
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3988 17134 4016 19110
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3988 16794 4016 17070
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3424 16584 3476 16590
rect 4172 16538 4200 20318
rect 4356 20058 4384 20946
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4448 19281 4476 26846
rect 4540 23746 4568 26959
rect 4632 26518 4660 26998
rect 4908 26858 4936 28086
rect 5184 27878 5212 28630
rect 5644 28422 5672 28902
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5262 28112 5318 28121
rect 5262 28047 5318 28056
rect 5276 27946 5304 28047
rect 5460 27946 5488 28358
rect 5644 27946 5672 28358
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5448 27940 5500 27946
rect 5448 27882 5500 27888
rect 5632 27940 5684 27946
rect 5632 27882 5684 27888
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 5538 27840 5594 27849
rect 5080 27328 5132 27334
rect 5080 27270 5132 27276
rect 5092 26994 5120 27270
rect 5080 26988 5132 26994
rect 5080 26930 5132 26936
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4620 26512 4672 26518
rect 4620 26454 4672 26460
rect 4988 26512 5040 26518
rect 4988 26454 5040 26460
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4816 25702 4844 26318
rect 4908 25974 4936 26318
rect 5000 26042 5028 26454
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 4896 25968 4948 25974
rect 4896 25910 4948 25916
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4712 25356 4764 25362
rect 4712 25298 4764 25304
rect 4620 25288 4672 25294
rect 4618 25256 4620 25265
rect 4672 25256 4674 25265
rect 4618 25191 4674 25200
rect 4632 24954 4660 25191
rect 4620 24948 4672 24954
rect 4620 24890 4672 24896
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4632 24410 4660 24618
rect 4724 24410 4752 25298
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4816 23866 4844 25638
rect 4908 25430 4936 25910
rect 4896 25424 4948 25430
rect 4896 25366 4948 25372
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4540 23718 4844 23746
rect 4528 23588 4580 23594
rect 4528 23530 4580 23536
rect 4434 19272 4490 19281
rect 4434 19207 4490 19216
rect 4540 17785 4568 23530
rect 4618 22536 4674 22545
rect 4618 22471 4674 22480
rect 4632 22234 4660 22471
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4724 21894 4752 21966
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21486 4752 21830
rect 4712 21480 4764 21486
rect 4712 21422 4764 21428
rect 4724 21146 4752 21422
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4632 20262 4660 20402
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4632 19802 4660 20198
rect 4724 19990 4752 20402
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4712 19848 4764 19854
rect 4632 19796 4712 19802
rect 4632 19790 4764 19796
rect 4632 19774 4752 19790
rect 4724 19310 4752 19774
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4816 18970 4844 23718
rect 4894 23624 4950 23633
rect 4894 23559 4950 23568
rect 5080 23588 5132 23594
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4816 18290 4844 18906
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4526 17776 4582 17785
rect 4526 17711 4582 17720
rect 4618 17232 4674 17241
rect 4908 17218 4936 23559
rect 5080 23530 5132 23536
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 5000 19378 5028 23462
rect 5092 23322 5120 23530
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 5184 23202 5212 27814
rect 5538 27775 5594 27784
rect 5354 27568 5410 27577
rect 5354 27503 5356 27512
rect 5408 27503 5410 27512
rect 5356 27474 5408 27480
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 5276 25498 5304 26862
rect 5368 26790 5396 27474
rect 5552 27402 5580 27775
rect 5644 27470 5672 27882
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5540 27396 5592 27402
rect 5540 27338 5592 27344
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5276 24750 5304 25434
rect 5264 24744 5316 24750
rect 5316 24692 5396 24698
rect 5264 24686 5396 24692
rect 5276 24670 5396 24686
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5276 23594 5304 24006
rect 5368 23730 5396 24670
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5092 23174 5212 23202
rect 5368 23186 5396 23666
rect 5356 23180 5408 23186
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5092 18154 5120 23174
rect 5356 23122 5408 23128
rect 5552 22080 5580 26726
rect 5644 26314 5672 27406
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5632 25424 5684 25430
rect 5632 25366 5684 25372
rect 5644 24954 5672 25366
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5736 24410 5764 30087
rect 6104 29782 6132 32014
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6736 32020 6788 32026
rect 6736 31962 6788 31968
rect 6840 31906 6868 39520
rect 7208 35057 7236 39520
rect 7194 35048 7250 35057
rect 7194 34983 7250 34992
rect 7012 34944 7064 34950
rect 7012 34886 7064 34892
rect 7024 34474 7052 34886
rect 7104 34536 7156 34542
rect 7104 34478 7156 34484
rect 7012 34468 7064 34474
rect 7012 34410 7064 34416
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6932 34134 6960 34342
rect 6920 34128 6972 34134
rect 6920 34070 6972 34076
rect 6932 33454 6960 34070
rect 7116 33658 7144 34478
rect 7288 34468 7340 34474
rect 7288 34410 7340 34416
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 6920 33448 6972 33454
rect 6920 33390 6972 33396
rect 6932 32978 6960 33390
rect 7104 33380 7156 33386
rect 7104 33322 7156 33328
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 7116 32774 7144 33322
rect 7300 32842 7328 34410
rect 7576 33386 7604 39520
rect 7944 35290 7972 39520
rect 8404 35850 8432 39520
rect 8220 35834 8432 35850
rect 8208 35828 8432 35834
rect 8260 35822 8432 35828
rect 8208 35770 8260 35776
rect 8392 35624 8444 35630
rect 8114 35592 8170 35601
rect 8392 35566 8444 35572
rect 8576 35624 8628 35630
rect 8576 35566 8628 35572
rect 8114 35527 8170 35536
rect 7932 35284 7984 35290
rect 7932 35226 7984 35232
rect 7930 35184 7986 35193
rect 7840 35148 7892 35154
rect 7930 35119 7986 35128
rect 7840 35090 7892 35096
rect 7852 34785 7880 35090
rect 7838 34776 7894 34785
rect 7838 34711 7840 34720
rect 7892 34711 7894 34720
rect 7840 34682 7892 34688
rect 7564 33380 7616 33386
rect 7564 33322 7616 33328
rect 7656 33380 7708 33386
rect 7656 33322 7708 33328
rect 7576 33289 7604 33322
rect 7562 33280 7618 33289
rect 7562 33215 7618 33224
rect 7668 33114 7696 33322
rect 7656 33108 7708 33114
rect 7656 33050 7708 33056
rect 7288 32836 7340 32842
rect 7288 32778 7340 32784
rect 7104 32768 7156 32774
rect 7104 32710 7156 32716
rect 7116 32026 7144 32710
rect 7668 32366 7696 33050
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7194 32056 7250 32065
rect 7104 32020 7156 32026
rect 7194 31991 7250 32000
rect 7104 31962 7156 31968
rect 7208 31958 7236 31991
rect 7668 31958 7696 32302
rect 6564 31878 6868 31906
rect 7196 31952 7248 31958
rect 7196 31894 7248 31900
rect 7380 31952 7432 31958
rect 7380 31894 7432 31900
rect 7656 31952 7708 31958
rect 7656 31894 7708 31900
rect 6564 31226 6592 31878
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6826 31784 6882 31793
rect 6656 31482 6684 31758
rect 6826 31719 6882 31728
rect 6644 31476 6696 31482
rect 6644 31418 6696 31424
rect 6564 31198 6684 31226
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29782 6684 31198
rect 6092 29776 6144 29782
rect 6092 29718 6144 29724
rect 6644 29776 6696 29782
rect 6644 29718 6696 29724
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 5816 29504 5868 29510
rect 5816 29446 5868 29452
rect 5828 26926 5856 29446
rect 6288 29034 6316 29650
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 6276 29028 6328 29034
rect 6276 28970 6328 28976
rect 5908 28552 5960 28558
rect 5908 28494 5960 28500
rect 5920 28218 5948 28494
rect 5908 28212 5960 28218
rect 5908 28154 5960 28160
rect 5816 26920 5868 26926
rect 5816 26862 5868 26868
rect 5724 24404 5776 24410
rect 5724 24346 5776 24352
rect 5736 23662 5764 24346
rect 5906 24304 5962 24313
rect 5906 24239 5962 24248
rect 5920 24206 5948 24239
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5920 23866 5948 24142
rect 5908 23860 5960 23866
rect 5828 23820 5908 23848
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5460 22052 5580 22080
rect 5460 22012 5488 22052
rect 5368 21984 5488 22012
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5184 18442 5212 21490
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19990 5304 20198
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5276 19514 5304 19926
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5184 18414 5304 18442
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 4618 17167 4674 17176
rect 4724 17190 4936 17218
rect 4434 16960 4490 16969
rect 4434 16895 4490 16904
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 3424 16526 3476 16532
rect 3068 16238 3188 16266
rect 3068 13802 3096 16238
rect 3436 15706 3464 16526
rect 4080 16510 4200 16538
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 15978 3556 16390
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 4080 16114 4108 16510
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 16017 4108 16050
rect 4066 16008 4122 16017
rect 3516 15972 3568 15978
rect 4066 15943 4122 15952
rect 3516 15914 3568 15920
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3148 14952 3200 14958
rect 3436 14929 3464 14962
rect 3528 14958 3556 15914
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3620 15638 3648 15846
rect 3608 15632 3660 15638
rect 3606 15600 3608 15609
rect 3660 15600 3662 15609
rect 3606 15535 3662 15544
rect 3620 15509 3648 15535
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 4172 14958 4200 16390
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 3516 14952 3568 14958
rect 3148 14894 3200 14900
rect 3422 14920 3478 14929
rect 3160 14278 3188 14894
rect 4160 14952 4212 14958
rect 3516 14894 3568 14900
rect 3606 14920 3662 14929
rect 3422 14855 3478 14864
rect 4160 14894 4212 14900
rect 3606 14855 3662 14864
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12918 3096 13262
rect 3056 12912 3108 12918
rect 3054 12880 3056 12889
rect 3108 12880 3110 12889
rect 3054 12815 3110 12824
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3068 12442 3096 12718
rect 3160 12714 3188 14214
rect 3252 13870 3280 14486
rect 3436 14074 3464 14758
rect 3620 14362 3648 14855
rect 3528 14334 3648 14362
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3528 13954 3556 14334
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3436 13926 3556 13954
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3068 11694 3096 12378
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3068 11354 3096 11630
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3146 10024 3202 10033
rect 3146 9959 3202 9968
rect 3160 9926 3188 9959
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 2884 9710 3004 9738
rect 2884 9450 2912 9710
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2792 9302 2912 9330
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2792 9042 2820 9114
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2884 8786 2912 9302
rect 2976 8974 3004 9590
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 9382 3096 9454
rect 3160 9382 3188 9862
rect 3252 9722 3280 13670
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3344 11082 3372 11562
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3068 9110 3096 9318
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2516 7942 2636 7970
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2318 7440 2374 7449
rect 2318 7375 2374 7384
rect 2056 6582 2176 6610
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1964 5370 1992 5714
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1964 4282 1992 4762
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1964 3738 1992 4218
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1674 3360 1730 3369
rect 1674 3295 1730 3304
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1490 1184 1546 1193
rect 1490 1119 1546 1128
rect 1780 480 1808 3470
rect 2056 2582 2084 6582
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 2148 480 2176 6394
rect 2240 6254 2268 6598
rect 2332 6458 2360 7375
rect 2516 7342 2544 7686
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2516 6934 2544 7278
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 6066 2268 6190
rect 2240 6038 2360 6066
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2240 4554 2268 5850
rect 2332 5166 2360 6038
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2332 4826 2360 5102
rect 2424 5030 2452 6598
rect 2412 5024 2464 5030
rect 2410 4992 2412 5001
rect 2464 4992 2466 5001
rect 2410 4927 2466 4936
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2502 4584 2558 4593
rect 2228 4548 2280 4554
rect 2502 4519 2558 4528
rect 2228 4490 2280 4496
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2424 3398 2452 3946
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2516 3346 2544 4519
rect 2608 3534 2636 7942
rect 2700 7886 2728 8230
rect 2792 8090 2820 8774
rect 2884 8758 3096 8786
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 7546 2728 7822
rect 2792 7546 2820 8026
rect 3068 7993 3096 8758
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6866 2820 7142
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5710 2728 6054
rect 2792 5817 2820 6666
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2962 5672 3018 5681
rect 2780 5636 2832 5642
rect 2962 5607 3018 5616
rect 2780 5578 2832 5584
rect 2792 4842 2820 5578
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2700 4826 2820 4842
rect 2688 4820 2820 4826
rect 2740 4814 2820 4820
rect 2688 4762 2740 4768
rect 2686 4720 2742 4729
rect 2686 4655 2742 4664
rect 2700 4622 2728 4655
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2700 3466 2728 4558
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2516 3318 2636 3346
rect 2608 480 2636 3318
rect 2792 3194 2820 4814
rect 2884 4049 2912 4966
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2884 2990 2912 3975
rect 2976 3670 3004 5607
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2964 3528 3016 3534
rect 2962 3496 2964 3505
rect 3016 3496 3018 3505
rect 2962 3431 3018 3440
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2976 2922 3004 3431
rect 3068 3058 3096 7919
rect 3160 5030 3188 8842
rect 3252 7528 3280 9386
rect 3344 8294 3372 11018
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3252 7500 3372 7528
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3194 3188 3538
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3252 2922 3280 5510
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2700 2378 2728 2790
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 2976 480 3004 2858
rect 3068 2582 3096 2858
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3344 480 3372 7500
rect 3436 6746 3464 13926
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3790 13832 3846 13841
rect 3528 9704 3556 13806
rect 3790 13767 3792 13776
rect 3844 13767 3846 13776
rect 3792 13738 3844 13744
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 4264 10606 4292 16186
rect 4356 15706 4384 16730
rect 4448 16658 4476 16895
rect 4632 16726 4660 17167
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4448 15910 4476 16594
rect 4632 16250 4660 16662
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4342 10704 4398 10713
rect 4342 10639 4398 10648
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3528 9676 3648 9704
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3528 9110 3556 9522
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3528 8634 3556 9046
rect 3620 8906 3648 9676
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 9489 3832 9590
rect 4080 9586 4108 9930
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3988 8090 4016 9522
rect 4172 9194 4200 9862
rect 4080 9178 4200 9194
rect 4068 9172 4200 9178
rect 4120 9166 4200 9172
rect 4068 9114 4120 9120
rect 4068 9036 4120 9042
rect 4264 9024 4292 10134
rect 4356 10130 4384 10639
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4356 9382 4384 10066
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 9217 4384 9318
rect 4342 9208 4398 9217
rect 4342 9143 4398 9152
rect 4120 8996 4292 9024
rect 4068 8978 4120 8984
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4080 7857 4108 8842
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 4264 7546 4292 8996
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8294 4384 8978
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 7886 4384 8230
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4068 6792 4120 6798
rect 3436 6718 3556 6746
rect 4068 6734 4120 6740
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5914 3464 6598
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 5098 3464 5510
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 4486 3464 5034
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 3398 3464 4422
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 2922 3464 3334
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3436 2825 3464 2858
rect 3528 2836 3556 6718
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 4080 6254 4108 6734
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 6118 4292 6190
rect 4356 6186 4384 6802
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 4080 5234 4108 5646
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4080 4826 4108 5170
rect 4158 4992 4214 5001
rect 4158 4927 4214 4936
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4172 4554 4200 4927
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3988 2990 4016 3538
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3422 2816 3478 2825
rect 3528 2808 3648 2836
rect 3422 2751 3478 2760
rect 3620 2360 3648 2808
rect 4080 2582 4108 3334
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 3528 2332 3648 2360
rect 3528 1986 3556 2332
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3528 1958 3832 1986
rect 3804 480 3832 1958
rect 4172 480 4200 4082
rect 4264 3924 4292 6054
rect 4448 5273 4476 15846
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4632 12374 4660 14214
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11801 4568 12038
rect 4526 11792 4582 11801
rect 4526 11727 4582 11736
rect 4632 11354 4660 12174
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4540 5409 4568 10542
rect 4724 10146 4752 17190
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4816 14550 4844 16118
rect 5000 16046 5028 17478
rect 5092 17105 5120 17682
rect 5078 17096 5134 17105
rect 5078 17031 5134 17040
rect 5092 16726 5120 17031
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 5078 16008 5134 16017
rect 5184 15978 5212 18294
rect 5276 16572 5304 18414
rect 5368 17066 5396 21984
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5552 21554 5580 21898
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5552 20602 5580 20878
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5460 19990 5488 20266
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5460 17814 5488 18158
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5460 17338 5488 17750
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5460 16794 5488 17274
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5552 16658 5580 19246
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5276 16544 5488 16572
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 16114 5304 16390
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5078 15943 5134 15952
rect 5172 15972 5224 15978
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4816 13530 4844 14486
rect 5000 14414 5028 15030
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5000 13530 5028 14350
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 11898 4936 12174
rect 5000 11898 5028 12310
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4908 11354 4936 11834
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5092 10554 5120 15943
rect 5172 15914 5224 15920
rect 5184 15706 5212 15914
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5276 15638 5304 16050
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5276 15026 5304 15574
rect 5354 15192 5410 15201
rect 5354 15127 5410 15136
rect 5368 15094 5396 15127
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5276 14550 5304 14962
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 13870 5212 14350
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5276 12306 5304 13942
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5368 13190 5396 13670
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12986 5396 13126
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5354 12880 5410 12889
rect 5460 12866 5488 16544
rect 5552 16250 5580 16594
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5552 15502 5580 16186
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5644 14618 5672 22646
rect 5828 22522 5856 23820
rect 5908 23802 5960 23808
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 5920 23118 5948 23530
rect 6012 23322 6040 28970
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6736 27600 6788 27606
rect 6736 27542 6788 27548
rect 6748 27441 6776 27542
rect 6734 27432 6790 27441
rect 6734 27367 6790 27376
rect 6644 26988 6696 26994
rect 6644 26930 6696 26936
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6092 26308 6144 26314
rect 6092 26250 6144 26256
rect 6104 24206 6132 26250
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6656 25362 6684 26930
rect 6736 25968 6788 25974
rect 6736 25910 6788 25916
rect 6644 25356 6696 25362
rect 6644 25298 6696 25304
rect 6656 24886 6684 25298
rect 6644 24880 6696 24886
rect 6644 24822 6696 24828
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6656 24274 6684 24822
rect 6644 24268 6696 24274
rect 6644 24210 6696 24216
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6104 23798 6132 24142
rect 6656 23866 6684 24210
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6092 23792 6144 23798
rect 6092 23734 6144 23740
rect 6000 23316 6052 23322
rect 6000 23258 6052 23264
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5920 22778 5948 23054
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 6012 22710 6040 23258
rect 6104 23118 6132 23734
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6104 22778 6132 23054
rect 6092 22772 6144 22778
rect 6092 22714 6144 22720
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 5828 22494 6040 22522
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5736 21049 5764 21830
rect 5908 21616 5960 21622
rect 5908 21558 5960 21564
rect 5722 21040 5778 21049
rect 5722 20975 5778 20984
rect 5920 20058 5948 21558
rect 6012 20890 6040 22494
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6104 21010 6132 21966
rect 6196 21690 6224 22102
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6012 20862 6132 20890
rect 6196 20874 6224 21626
rect 6288 21622 6316 21966
rect 6644 21684 6696 21690
rect 6644 21626 6696 21632
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 6012 20398 6040 20742
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5736 16998 5764 17818
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16697 5764 16934
rect 5722 16688 5778 16697
rect 5722 16623 5778 16632
rect 5722 15192 5778 15201
rect 5722 15127 5778 15136
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5540 14544 5592 14550
rect 5736 14498 5764 15127
rect 5828 15065 5856 19314
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 16250 6040 16662
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5814 15056 5870 15065
rect 5814 14991 5870 15000
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5540 14486 5592 14492
rect 5552 13462 5580 14486
rect 5644 14470 5764 14498
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 12918 5580 13398
rect 5410 12838 5488 12866
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5354 12815 5410 12824
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 4908 10526 5120 10554
rect 4724 10118 4844 10146
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 9382 4752 9998
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9110 4752 9318
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4710 8664 4766 8673
rect 4710 8599 4766 8608
rect 4618 6896 4674 6905
rect 4618 6831 4674 6840
rect 4526 5400 4582 5409
rect 4526 5335 4582 5344
rect 4434 5264 4490 5273
rect 4434 5199 4490 5208
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4729 4476 4966
rect 4434 4720 4490 4729
rect 4344 4684 4396 4690
rect 4434 4655 4490 4664
rect 4344 4626 4396 4632
rect 4356 4282 4384 4626
rect 4540 4593 4568 5335
rect 4526 4584 4582 4593
rect 4526 4519 4582 4528
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4344 3936 4396 3942
rect 4264 3896 4344 3924
rect 4344 3878 4396 3884
rect 4356 3602 4384 3878
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 3097 4292 3334
rect 4250 3088 4306 3097
rect 4250 3023 4306 3032
rect 4356 2990 4384 3538
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4252 2508 4304 2514
rect 4356 2496 4384 2926
rect 4304 2468 4384 2496
rect 4252 2450 4304 2456
rect 4632 626 4660 6831
rect 4724 3534 4752 8599
rect 4816 8090 4844 10118
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7410 4844 7686
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4816 7313 4844 7346
rect 4802 7304 4858 7313
rect 4802 7239 4858 7248
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4816 3942 4844 4694
rect 4908 4690 4936 10526
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 9450 5028 10406
rect 5262 10160 5318 10169
rect 5262 10095 5318 10104
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5000 8634 5028 9386
rect 5092 9081 5120 9522
rect 5184 9450 5212 9862
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5184 9178 5212 9386
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5078 9072 5134 9081
rect 5276 9058 5304 10095
rect 5078 9007 5134 9016
rect 5184 9030 5304 9058
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5000 4758 5028 8026
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4804 3936 4856 3942
rect 4908 3913 4936 4626
rect 5184 4146 5212 9030
rect 5368 8673 5396 12815
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 12442 5488 12718
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5460 11218 5488 12378
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10826 5488 11154
rect 5644 11121 5672 14470
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 5736 13938 5764 14282
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5722 13696 5778 13705
rect 5722 13631 5778 13640
rect 5630 11112 5686 11121
rect 5630 11047 5686 11056
rect 5460 10810 5580 10826
rect 5460 10804 5592 10810
rect 5460 10798 5540 10804
rect 5540 10746 5592 10752
rect 5552 10130 5580 10746
rect 5644 10169 5672 11047
rect 5630 10160 5686 10169
rect 5540 10124 5592 10130
rect 5630 10095 5686 10104
rect 5540 10066 5592 10072
rect 5552 9042 5580 10066
rect 5630 10024 5686 10033
rect 5630 9959 5686 9968
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5354 8664 5410 8673
rect 5354 8599 5410 8608
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 7206 5304 7686
rect 5460 7342 5488 7958
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6118 5304 7142
rect 5460 7002 5488 7278
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5354 5536 5410 5545
rect 5354 5471 5410 5480
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5080 4072 5132 4078
rect 5276 4049 5304 4082
rect 5080 4014 5132 4020
rect 5262 4040 5318 4049
rect 4988 3936 5040 3942
rect 4804 3878 4856 3884
rect 4894 3904 4950 3913
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4816 3233 4844 3878
rect 4988 3878 5040 3884
rect 4894 3839 4950 3848
rect 5000 3398 5028 3878
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4802 3224 4858 3233
rect 4802 3159 4858 3168
rect 5000 2990 5028 3334
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5092 2836 5120 4014
rect 5262 3975 5318 3984
rect 4540 598 4660 626
rect 5000 2808 5120 2836
rect 4540 480 4568 598
rect 5000 480 5028 2808
rect 5368 480 5396 5471
rect 5644 5114 5672 9959
rect 5736 8294 5764 13631
rect 5828 12628 5856 14758
rect 5920 13462 5948 15438
rect 6104 14906 6132 20862
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6182 20360 6238 20369
rect 6182 20295 6238 20304
rect 6012 14878 6132 14906
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5920 12782 5948 13398
rect 6012 12918 6040 14878
rect 6196 14822 6224 20295
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6656 20058 6684 21626
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6656 15201 6684 19450
rect 6642 15192 6698 15201
rect 6642 15127 6698 15136
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6196 14074 6224 14554
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6656 13870 6684 14350
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6104 13190 6132 13738
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5828 12600 5948 12628
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 8498 5856 9318
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5828 8090 5856 8434
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5644 5086 5764 5114
rect 5448 5024 5500 5030
rect 5632 5024 5684 5030
rect 5500 4984 5580 5012
rect 5448 4966 5500 4972
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 3670 5488 4422
rect 5552 3924 5580 4984
rect 5632 4966 5684 4972
rect 5644 4146 5672 4966
rect 5736 4690 5764 5086
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5736 4282 5764 4626
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5724 3936 5776 3942
rect 5552 3896 5724 3924
rect 5724 3878 5776 3884
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5736 3194 5764 3878
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5920 3074 5948 12600
rect 6012 10169 6040 12854
rect 6104 11286 6132 13126
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6104 10810 6132 11222
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5998 10160 6054 10169
rect 5998 10095 6054 10104
rect 6012 8566 6040 10095
rect 6196 9058 6224 13806
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6656 10198 6684 11290
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9654 6408 10066
rect 6656 9722 6684 10134
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6196 9030 6408 9058
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6092 8288 6144 8294
rect 6288 8276 6316 8502
rect 6380 8362 6408 9030
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6092 8230 6144 8236
rect 6196 8248 6316 8276
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 5736 3046 5948 3074
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2582 5488 2790
rect 5538 2680 5594 2689
rect 5538 2615 5540 2624
rect 5592 2615 5594 2624
rect 5540 2586 5592 2592
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5736 480 5764 3046
rect 6012 1442 6040 3839
rect 6104 2553 6132 8230
rect 6090 2544 6146 2553
rect 6090 2479 6146 2488
rect 6196 1578 6224 8248
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6748 5545 6776 25910
rect 6840 25809 6868 31719
rect 7208 31482 7236 31894
rect 7196 31476 7248 31482
rect 7116 31436 7196 31464
rect 7012 30320 7064 30326
rect 7012 30262 7064 30268
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6932 27062 6960 27542
rect 7024 27470 7052 30262
rect 7116 29073 7144 31436
rect 7196 31418 7248 31424
rect 7392 31414 7420 31894
rect 7380 31408 7432 31414
rect 7378 31376 7380 31385
rect 7432 31376 7434 31385
rect 7378 31311 7434 31320
rect 7392 31285 7420 31311
rect 7944 30841 7972 35119
rect 8128 33046 8156 35527
rect 8208 33448 8260 33454
rect 8208 33390 8260 33396
rect 8116 33040 8168 33046
rect 8036 33000 8116 33028
rect 8036 31890 8064 33000
rect 8116 32982 8168 32988
rect 8116 32904 8168 32910
rect 8114 32872 8116 32881
rect 8168 32872 8170 32881
rect 8114 32807 8170 32816
rect 8220 32824 8248 33390
rect 8128 31958 8156 32807
rect 8220 32796 8340 32824
rect 8312 32570 8340 32796
rect 8404 32570 8432 35566
rect 8484 34672 8536 34678
rect 8482 34640 8484 34649
rect 8536 34640 8538 34649
rect 8482 34575 8538 34584
rect 8588 34542 8616 35566
rect 8772 34746 8800 39520
rect 9140 37346 9168 39520
rect 9140 37318 9352 37346
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9324 35834 9352 37318
rect 9312 35828 9364 35834
rect 9312 35770 9364 35776
rect 9508 35290 9536 39520
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9496 35284 9548 35290
rect 9496 35226 9548 35232
rect 9772 35148 9824 35154
rect 9772 35090 9824 35096
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 8760 34740 8812 34746
rect 8760 34682 8812 34688
rect 8864 34610 8892 34886
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8852 34604 8904 34610
rect 8772 34564 8852 34592
rect 8576 34536 8628 34542
rect 8576 34478 8628 34484
rect 8484 33448 8536 33454
rect 8484 33390 8536 33396
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8392 32564 8444 32570
rect 8392 32506 8444 32512
rect 8496 32298 8524 33390
rect 8484 32292 8536 32298
rect 8484 32234 8536 32240
rect 8116 31952 8168 31958
rect 8116 31894 8168 31900
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 7930 30832 7986 30841
rect 7930 30767 7986 30776
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 7392 30122 7420 30534
rect 7196 30116 7248 30122
rect 7196 30058 7248 30064
rect 7380 30116 7432 30122
rect 7380 30058 7432 30064
rect 7208 29578 7236 30058
rect 7288 29708 7340 29714
rect 7288 29650 7340 29656
rect 7196 29572 7248 29578
rect 7196 29514 7248 29520
rect 7300 29510 7328 29650
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 7102 29064 7158 29073
rect 7300 29034 7328 29446
rect 7392 29306 7420 30058
rect 7472 29504 7524 29510
rect 7472 29446 7524 29452
rect 7380 29300 7432 29306
rect 7380 29242 7432 29248
rect 7378 29200 7434 29209
rect 7378 29135 7434 29144
rect 7102 28999 7158 29008
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 7392 28966 7420 29135
rect 7104 28960 7156 28966
rect 7104 28902 7156 28908
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7116 28558 7144 28902
rect 7392 28762 7420 28902
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7392 28665 7420 28698
rect 7378 28656 7434 28665
rect 7378 28591 7434 28600
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7116 27146 7144 28494
rect 7484 28082 7512 29446
rect 7562 29200 7618 29209
rect 7562 29135 7564 29144
rect 7616 29135 7618 29144
rect 7564 29106 7616 29112
rect 7562 29064 7618 29073
rect 7562 28999 7618 29008
rect 7748 29028 7800 29034
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7196 27464 7248 27470
rect 7196 27406 7248 27412
rect 7286 27432 7342 27441
rect 7024 27118 7144 27146
rect 7208 27130 7236 27406
rect 7286 27367 7342 27376
rect 7196 27124 7248 27130
rect 6920 27056 6972 27062
rect 6920 26998 6972 27004
rect 6932 26586 6960 26998
rect 7024 26994 7052 27118
rect 7196 27066 7248 27072
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 7012 26852 7064 26858
rect 7012 26794 7064 26800
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 7024 26450 7052 26794
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 7116 26314 7144 26930
rect 7104 26308 7156 26314
rect 7104 26250 7156 26256
rect 7300 26194 7328 27367
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7116 26166 7328 26194
rect 6826 25800 6882 25809
rect 6826 25735 6882 25744
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 6826 23488 6882 23497
rect 6826 23423 6882 23432
rect 6840 23254 6868 23423
rect 6828 23248 6880 23254
rect 6828 23190 6880 23196
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 6932 21570 6960 22510
rect 7024 22030 7052 23802
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6840 21554 6960 21570
rect 6828 21548 6960 21554
rect 6880 21542 6960 21548
rect 6828 21490 6880 21496
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6828 20256 6880 20262
rect 6932 20210 6960 20946
rect 7024 20534 7052 21830
rect 7116 21486 7144 26166
rect 7392 26042 7420 26726
rect 7576 26625 7604 28999
rect 7748 28970 7800 28976
rect 7760 28626 7788 28970
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7748 28620 7800 28626
rect 7748 28562 7800 28568
rect 7654 28112 7710 28121
rect 7654 28047 7710 28056
rect 7562 26616 7618 26625
rect 7562 26551 7618 26560
rect 7564 26512 7616 26518
rect 7564 26454 7616 26460
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7380 26036 7432 26042
rect 7380 25978 7432 25984
rect 7484 25974 7512 26318
rect 7472 25968 7524 25974
rect 7470 25936 7472 25945
rect 7524 25936 7526 25945
rect 7470 25871 7526 25880
rect 7484 25845 7512 25871
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7208 24954 7236 25094
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 7208 24342 7236 24890
rect 7576 24818 7604 26454
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7196 24336 7248 24342
rect 7196 24278 7248 24284
rect 7208 23730 7236 24278
rect 7564 23792 7616 23798
rect 7562 23760 7564 23769
rect 7616 23760 7618 23769
rect 7196 23724 7248 23730
rect 7562 23695 7618 23704
rect 7196 23666 7248 23672
rect 7208 23322 7236 23666
rect 7576 23526 7604 23695
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7208 22778 7236 23054
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7288 22160 7340 22166
rect 7288 22102 7340 22108
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7300 21350 7328 22102
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 21146 7328 21286
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7012 20528 7064 20534
rect 7012 20470 7064 20476
rect 7116 20330 7144 20878
rect 7392 20602 7420 21966
rect 7576 21350 7604 22034
rect 7668 21554 7696 28047
rect 7760 27334 7788 28562
rect 7852 28422 7880 28902
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7852 28218 7880 28358
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 7760 26382 7788 27270
rect 7944 26602 7972 30767
rect 8036 26761 8064 31350
rect 8208 30184 8260 30190
rect 8208 30126 8260 30132
rect 8116 29776 8168 29782
rect 8116 29718 8168 29724
rect 8128 29034 8156 29718
rect 8116 29028 8168 29034
rect 8116 28970 8168 28976
rect 8022 26752 8078 26761
rect 8128 26738 8156 28970
rect 8220 28778 8248 30126
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8496 29034 8524 29446
rect 8484 29028 8536 29034
rect 8484 28970 8536 28976
rect 8220 28762 8340 28778
rect 8220 28756 8352 28762
rect 8220 28750 8300 28756
rect 8300 28698 8352 28704
rect 8312 27946 8340 28698
rect 8300 27940 8352 27946
rect 8220 27900 8300 27928
rect 8220 27606 8248 27900
rect 8300 27882 8352 27888
rect 8496 27878 8524 28970
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8208 27600 8260 27606
rect 8208 27542 8260 27548
rect 8298 27568 8354 27577
rect 8220 26858 8248 27542
rect 8298 27503 8300 27512
rect 8352 27503 8354 27512
rect 8300 27474 8352 27480
rect 8496 27470 8524 27814
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8208 26852 8260 26858
rect 8208 26794 8260 26800
rect 8128 26710 8248 26738
rect 8022 26687 8078 26696
rect 7944 26574 8156 26602
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7760 25702 7788 26318
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7852 25770 7880 26182
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7840 25764 7892 25770
rect 7840 25706 7892 25712
rect 7748 25696 7800 25702
rect 7748 25638 7800 25644
rect 7852 24954 7880 25706
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7852 22778 7880 24550
rect 7944 23866 7972 25842
rect 8022 25528 8078 25537
rect 8022 25463 8024 25472
rect 8076 25463 8078 25472
rect 8024 25434 8076 25440
rect 8128 25378 8156 26574
rect 8036 25350 8156 25378
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7944 23322 7972 23598
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7944 23089 7972 23258
rect 7930 23080 7986 23089
rect 7930 23015 7986 23024
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7852 22545 7880 22714
rect 7838 22536 7894 22545
rect 7838 22471 7894 22480
rect 7852 22438 7880 22471
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 8036 22234 8064 25350
rect 8114 24848 8170 24857
rect 8114 24783 8170 24792
rect 8128 23526 8156 24783
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8128 22545 8156 22918
rect 8114 22536 8170 22545
rect 8114 22471 8170 22480
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 21690 7880 21966
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 6880 20204 6960 20210
rect 6828 20198 6960 20204
rect 6840 20182 6960 20198
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 18970 6868 19246
rect 6932 19174 6960 20182
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7024 19242 7052 19994
rect 7116 19786 7144 20266
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7102 19408 7158 19417
rect 7102 19343 7158 19352
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 7024 18834 7052 19178
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7024 18358 7052 18770
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 16153 6960 17478
rect 6918 16144 6974 16153
rect 6918 16079 6974 16088
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15156 6880 15162
rect 6932 15144 6960 15506
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7024 15162 7052 15438
rect 6880 15116 6960 15144
rect 7012 15156 7064 15162
rect 6828 15098 6880 15104
rect 7012 15098 7064 15104
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6840 5778 6868 14826
rect 7012 14000 7064 14006
rect 7010 13968 7012 13977
rect 7064 13968 7066 13977
rect 7010 13903 7066 13912
rect 7116 13818 7144 19343
rect 7392 19310 7420 20538
rect 7484 20262 7512 21014
rect 7576 20466 7604 21286
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7562 20224 7618 20233
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7484 18698 7512 20198
rect 7562 20159 7618 20168
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7484 17882 7512 18294
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7392 17338 7420 17682
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 7024 13790 7144 13818
rect 6932 13530 6960 13738
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7024 12646 7052 13790
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12442 7052 12582
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 9178 6960 10406
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6932 8430 6960 9114
rect 7010 9072 7066 9081
rect 7010 9007 7066 9016
rect 7024 8634 7052 9007
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6920 7268 6972 7274
rect 7116 7256 7144 13670
rect 7208 9489 7236 17138
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7392 14618 7420 16118
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7392 13938 7420 14554
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13938 7512 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7392 13190 7420 13670
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 9625 7328 12582
rect 7392 12170 7420 13126
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7484 11558 7512 12310
rect 7472 11552 7524 11558
rect 7378 11520 7434 11529
rect 7576 11529 7604 20159
rect 7668 18306 7696 21082
rect 7760 18902 7788 21558
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7930 19952 7986 19961
rect 7852 19310 7880 19926
rect 7930 19887 7986 19896
rect 7944 19854 7972 19887
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7944 19514 7972 19790
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7852 18970 7880 19246
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7760 18426 7788 18838
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7944 18358 7972 18838
rect 7932 18352 7984 18358
rect 7668 18278 7788 18306
rect 7932 18294 7984 18300
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7668 15978 7696 16390
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7668 14346 7696 15914
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7668 11898 7696 12242
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7472 11494 7524 11500
rect 7562 11520 7618 11529
rect 7378 11455 7434 11464
rect 7392 11014 7420 11455
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10470 7420 10950
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7286 9616 7342 9625
rect 7286 9551 7342 9560
rect 7194 9480 7250 9489
rect 7194 9415 7250 9424
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 7993 7236 9318
rect 7392 9024 7420 10406
rect 7484 9654 7512 11494
rect 7562 11455 7618 11464
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7576 10674 7604 11290
rect 7668 11082 7696 11834
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7392 8996 7512 9024
rect 7484 8945 7512 8996
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7378 8392 7434 8401
rect 7378 8327 7380 8336
rect 7432 8327 7434 8336
rect 7380 8298 7432 8304
rect 7194 7984 7250 7993
rect 7194 7919 7250 7928
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7116 7228 7328 7256
rect 6920 7210 6972 7216
rect 6932 7002 6960 7210
rect 7194 7168 7250 7177
rect 7194 7103 7250 7112
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6734 5536 6790 5545
rect 6734 5471 6790 5480
rect 6840 5370 6868 5714
rect 6932 5681 6960 6190
rect 7116 6118 7144 6734
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6918 5672 6974 5681
rect 6918 5607 6974 5616
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7010 5400 7066 5409
rect 6828 5364 6880 5370
rect 7010 5335 7012 5344
rect 6828 5306 6880 5312
rect 7064 5335 7066 5344
rect 7012 5306 7064 5312
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6288 3126 6316 3538
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6196 1550 6592 1578
rect 6012 1414 6224 1442
rect 6196 480 6224 1414
rect 6564 480 6592 1550
rect 6656 1426 6684 4762
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6840 3777 6868 4218
rect 6932 4010 6960 4490
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6826 3768 6882 3777
rect 6826 3703 6882 3712
rect 6932 3466 6960 3946
rect 7024 3942 7052 4966
rect 7116 4593 7144 5510
rect 7208 5098 7236 7103
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7300 4690 7328 7228
rect 7392 5846 7420 7278
rect 7484 6905 7512 8871
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7470 6896 7526 6905
rect 7470 6831 7526 6840
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7392 5370 7420 5782
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7380 4616 7432 4622
rect 7102 4584 7158 4593
rect 7380 4558 7432 4564
rect 7102 4519 7158 4528
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 7024 2378 7052 3878
rect 7116 3670 7144 4218
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7208 2990 7236 4422
rect 7392 4214 7420 4558
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7392 2922 7420 4014
rect 7484 3670 7512 5102
rect 7576 4758 7604 6938
rect 7760 6905 7788 18278
rect 8036 16697 8064 21490
rect 8220 17202 8248 26710
rect 8588 25702 8616 34478
rect 8772 33046 8800 34564
rect 8852 34546 8904 34552
rect 9784 34406 9812 35090
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 9772 34400 9824 34406
rect 9772 34342 9824 34348
rect 8864 33862 8892 34342
rect 8852 33856 8904 33862
rect 8852 33798 8904 33804
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9402 33416 9458 33425
rect 8852 33380 8904 33386
rect 9402 33351 9458 33360
rect 8852 33322 8904 33328
rect 8864 33114 8892 33322
rect 9310 33280 9366 33289
rect 9310 33215 9366 33224
rect 8852 33108 8904 33114
rect 8852 33050 8904 33056
rect 8760 33040 8812 33046
rect 8760 32982 8812 32988
rect 8668 32564 8720 32570
rect 8668 32506 8720 32512
rect 8484 25696 8536 25702
rect 8484 25638 8536 25644
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8298 25528 8354 25537
rect 8298 25463 8354 25472
rect 8312 24750 8340 25463
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8312 22574 8340 24686
rect 8404 23633 8432 24686
rect 8496 24410 8524 25638
rect 8588 24857 8616 25638
rect 8574 24848 8630 24857
rect 8574 24783 8630 24792
rect 8576 24676 8628 24682
rect 8576 24618 8628 24624
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8588 24206 8616 24618
rect 8680 24614 8708 32506
rect 8772 32502 8800 32982
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8760 32496 8812 32502
rect 8760 32438 8812 32444
rect 8852 31884 8904 31890
rect 8852 31826 8904 31832
rect 8760 31680 8812 31686
rect 8760 31622 8812 31628
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 23730 8616 24142
rect 8772 23769 8800 31622
rect 8758 23760 8814 23769
rect 8576 23724 8628 23730
rect 8758 23695 8814 23704
rect 8576 23666 8628 23672
rect 8390 23624 8446 23633
rect 8390 23559 8446 23568
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 8390 23080 8446 23089
rect 8390 23015 8446 23024
rect 8484 23044 8536 23050
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8312 20806 8340 21354
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8312 17105 8340 20742
rect 8298 17096 8354 17105
rect 8298 17031 8354 17040
rect 8022 16688 8078 16697
rect 8022 16623 8078 16632
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7852 15162 7880 16050
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7944 12986 7972 15982
rect 8128 14958 8156 16594
rect 8312 15910 8340 17031
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8220 14890 8248 15506
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 8036 14074 8064 14486
rect 8312 14074 8340 14554
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8036 13870 8064 14010
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8022 13696 8078 13705
rect 8022 13631 8078 13640
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7944 12238 7972 12922
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11354 7880 11698
rect 7944 11626 7972 12174
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7852 8906 7880 9386
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7838 8528 7894 8537
rect 7944 8514 7972 9046
rect 7894 8486 7972 8514
rect 7838 8463 7840 8472
rect 7892 8463 7894 8472
rect 7840 8434 7892 8440
rect 8036 7562 8064 13631
rect 8312 12714 8340 13874
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 11898 8248 12582
rect 8312 12442 8340 12650
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8404 12209 8432 23015
rect 8484 22986 8536 22992
rect 8496 22506 8524 22986
rect 8588 22778 8616 23190
rect 8760 23180 8812 23186
rect 8760 23122 8812 23128
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8496 22234 8524 22442
rect 8772 22234 8800 23122
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8760 21412 8812 21418
rect 8760 21354 8812 21360
rect 8772 20806 8800 21354
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8496 20398 8524 20742
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8496 18970 8524 20334
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8496 18290 8524 18906
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8496 16130 8524 18090
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8588 17338 8616 17750
rect 8668 17672 8720 17678
rect 8666 17640 8668 17649
rect 8720 17640 8722 17649
rect 8666 17575 8722 17584
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8680 17270 8708 17575
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8496 16102 8708 16130
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8496 15706 8524 15982
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8574 15056 8630 15065
rect 8574 14991 8630 15000
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8496 14414 8524 14826
rect 8588 14550 8616 14991
rect 8680 14550 8708 16102
rect 8772 14822 8800 18294
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8864 14618 8892 31826
rect 9324 31686 9352 33215
rect 9416 32298 9444 33351
rect 9508 32570 9536 33798
rect 9680 33312 9732 33318
rect 9680 33254 9732 33260
rect 9586 33144 9642 33153
rect 9586 33079 9642 33088
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 9600 32473 9628 33079
rect 9692 33046 9720 33254
rect 9680 33040 9732 33046
rect 9784 33017 9812 34342
rect 9680 32982 9732 32988
rect 9770 33008 9826 33017
rect 9770 32943 9826 32952
rect 9586 32464 9642 32473
rect 9586 32399 9642 32408
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 9416 32026 9444 32234
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9312 31680 9364 31686
rect 9312 31622 9364 31628
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9312 31136 9364 31142
rect 9312 31078 9364 31084
rect 9324 30598 9352 31078
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 9324 30394 9352 30534
rect 9312 30388 9364 30394
rect 9312 30330 9364 30336
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9324 26024 9352 26454
rect 9232 25996 9352 26024
rect 9128 25968 9180 25974
rect 9126 25936 9128 25945
rect 9180 25936 9182 25945
rect 9126 25871 9182 25880
rect 9232 25702 9260 25996
rect 9312 25832 9364 25838
rect 9312 25774 9364 25780
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9324 23050 9352 25774
rect 9416 25537 9444 31962
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9402 25528 9458 25537
rect 9402 25463 9458 25472
rect 9404 25424 9456 25430
rect 9404 25366 9456 25372
rect 9416 23662 9444 25366
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 9416 23118 9444 23462
rect 9508 23186 9536 26250
rect 9600 23905 9628 32399
rect 9876 31822 9904 35430
rect 9968 35290 9996 39520
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 10336 34746 10364 39520
rect 10704 35834 10732 39520
rect 10966 36680 11022 36689
rect 10966 36615 11022 36624
rect 10980 36378 11008 36615
rect 10968 36372 11020 36378
rect 10968 36314 11020 36320
rect 10784 36236 10836 36242
rect 10784 36178 10836 36184
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 10796 35578 10824 36178
rect 11072 35834 11100 39520
rect 11336 36712 11388 36718
rect 11336 36654 11388 36660
rect 11060 35828 11112 35834
rect 11060 35770 11112 35776
rect 10704 35550 10824 35578
rect 11152 35624 11204 35630
rect 11152 35566 11204 35572
rect 10704 35494 10732 35550
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10138 34640 10194 34649
rect 10138 34575 10194 34584
rect 10152 34542 10180 34575
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 9968 33046 9996 34002
rect 10048 33108 10100 33114
rect 10048 33050 10100 33056
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 9968 32314 9996 32982
rect 10060 32434 10088 33050
rect 10048 32428 10100 32434
rect 10048 32370 10100 32376
rect 9968 32286 10088 32314
rect 9956 31952 10008 31958
rect 9956 31894 10008 31900
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9680 31748 9732 31754
rect 9680 31690 9732 31696
rect 9692 26602 9720 31690
rect 9772 31680 9824 31686
rect 9772 31622 9824 31628
rect 9784 30705 9812 31622
rect 9968 31414 9996 31894
rect 10060 31890 10088 32286
rect 10048 31884 10100 31890
rect 10048 31826 10100 31832
rect 10060 31482 10088 31826
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 9956 31408 10008 31414
rect 9956 31350 10008 31356
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9770 30696 9826 30705
rect 9770 30631 9826 30640
rect 9772 30116 9824 30122
rect 9772 30058 9824 30064
rect 9784 27402 9812 30058
rect 9876 29050 9904 31078
rect 9968 30938 9996 31350
rect 10048 31340 10100 31346
rect 10048 31282 10100 31288
rect 9956 30932 10008 30938
rect 9956 30874 10008 30880
rect 9954 30152 10010 30161
rect 9954 30087 10010 30096
rect 9968 29170 9996 30087
rect 10060 29578 10088 31282
rect 10152 30258 10180 34478
rect 10416 34400 10468 34406
rect 10416 34342 10468 34348
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 10244 33454 10272 34070
rect 10232 33448 10284 33454
rect 10232 33390 10284 33396
rect 10244 33318 10272 33390
rect 10232 33312 10284 33318
rect 10232 33254 10284 33260
rect 10244 32978 10272 33254
rect 10322 33008 10378 33017
rect 10232 32972 10284 32978
rect 10322 32943 10378 32952
rect 10232 32914 10284 32920
rect 10244 32570 10272 32914
rect 10232 32564 10284 32570
rect 10232 32506 10284 32512
rect 10232 31816 10284 31822
rect 10336 31770 10364 32943
rect 10232 31758 10284 31764
rect 10244 31385 10272 31758
rect 10326 31742 10364 31770
rect 10326 31668 10354 31742
rect 10326 31640 10364 31668
rect 10336 31482 10364 31640
rect 10324 31476 10376 31482
rect 10324 31418 10376 31424
rect 10230 31376 10286 31385
rect 10230 31311 10286 31320
rect 10244 30938 10272 31311
rect 10428 31260 10456 34342
rect 10508 31476 10560 31482
rect 10508 31418 10560 31424
rect 10336 31232 10456 31260
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 10140 30116 10192 30122
rect 10140 30058 10192 30064
rect 10048 29572 10100 29578
rect 10048 29514 10100 29520
rect 10152 29510 10180 30058
rect 10140 29504 10192 29510
rect 10140 29446 10192 29452
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10140 29232 10192 29238
rect 10140 29174 10192 29180
rect 9956 29164 10008 29170
rect 9956 29106 10008 29112
rect 9876 29022 10088 29050
rect 9864 28416 9916 28422
rect 9864 28358 9916 28364
rect 9876 27946 9904 28358
rect 9864 27940 9916 27946
rect 9864 27882 9916 27888
rect 9876 27441 9904 27882
rect 10060 27452 10088 29022
rect 10152 27606 10180 29174
rect 10244 28762 10272 29242
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10244 28218 10272 28698
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10140 27600 10192 27606
rect 10140 27542 10192 27548
rect 10232 27464 10284 27470
rect 9862 27432 9918 27441
rect 9772 27396 9824 27402
rect 10060 27424 10180 27452
rect 9862 27367 9918 27376
rect 9772 27338 9824 27344
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 10060 27062 10088 27270
rect 10048 27056 10100 27062
rect 10046 27024 10048 27033
rect 10100 27024 10102 27033
rect 10046 26959 10102 26968
rect 10152 26897 10180 27424
rect 10232 27406 10284 27412
rect 10244 27130 10272 27406
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10138 26888 10194 26897
rect 10138 26823 10194 26832
rect 10138 26752 10194 26761
rect 10138 26687 10194 26696
rect 9692 26574 9904 26602
rect 9680 26444 9732 26450
rect 9680 26386 9732 26392
rect 9692 25838 9720 26386
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9876 24614 9904 26574
rect 10152 26382 10180 26687
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9586 23896 9642 23905
rect 9586 23831 9642 23840
rect 9586 23760 9642 23769
rect 9586 23695 9642 23704
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9600 22930 9628 23695
rect 9876 23497 9904 24550
rect 9862 23488 9918 23497
rect 9862 23423 9918 23432
rect 9968 23322 9996 25910
rect 10152 25498 10180 26318
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10244 24800 10272 27066
rect 10060 24772 10272 24800
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9324 22902 9628 22930
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9218 19272 9274 19281
rect 9218 19207 9274 19216
rect 9232 18970 9260 19207
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9324 18358 9352 22902
rect 9494 22808 9550 22817
rect 9494 22743 9550 22752
rect 9864 22772 9916 22778
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9416 20097 9444 20742
rect 9402 20088 9458 20097
rect 9402 20023 9404 20032
rect 9456 20023 9458 20032
rect 9404 19994 9456 20000
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9324 16794 9352 18158
rect 9508 18086 9536 22743
rect 9864 22714 9916 22720
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9692 21418 9720 22646
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9784 20505 9812 21558
rect 9770 20496 9826 20505
rect 9770 20431 9826 20440
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9600 19242 9628 20198
rect 9876 19394 9904 22714
rect 9968 22574 9996 23258
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 10060 21706 10088 24772
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 10152 24206 10180 24618
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10138 22536 10194 22545
rect 10138 22471 10140 22480
rect 10192 22471 10194 22480
rect 10140 22442 10192 22448
rect 10152 22234 10180 22442
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10244 22166 10272 24210
rect 10336 22778 10364 31232
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10428 28218 10456 30194
rect 10416 28212 10468 28218
rect 10416 28154 10468 28160
rect 10428 28121 10456 28154
rect 10414 28112 10470 28121
rect 10414 28047 10470 28056
rect 10428 27878 10456 28047
rect 10416 27872 10468 27878
rect 10416 27814 10468 27820
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10428 27130 10456 27610
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10060 21678 10180 21706
rect 9954 20088 10010 20097
rect 9954 20023 10010 20032
rect 9784 19366 9904 19394
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9692 18970 9720 19178
rect 9784 19156 9812 19366
rect 9864 19304 9916 19310
rect 9968 19292 9996 20023
rect 9916 19264 9996 19292
rect 9864 19246 9916 19252
rect 10048 19168 10100 19174
rect 9784 19128 9996 19156
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9692 18714 9720 18906
rect 9692 18686 9812 18714
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9416 16250 9444 17002
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 15366 9444 15846
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 13870 8524 14350
rect 8680 14226 8708 14486
rect 8680 14198 8800 14226
rect 8772 14074 8800 14198
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8390 12200 8446 12209
rect 8390 12135 8446 12144
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8404 11354 8432 12135
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 9926 8156 10474
rect 8404 10266 8432 11290
rect 8496 11150 8524 13806
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8588 11898 8616 12378
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 10810 8524 11086
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8496 10266 8524 10746
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8128 8974 8156 9862
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8090 8156 8910
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8673 8248 8842
rect 8206 8664 8262 8673
rect 8206 8599 8208 8608
rect 8260 8599 8262 8608
rect 8208 8570 8260 8576
rect 8220 8430 8248 8570
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8404 8022 8432 10202
rect 8496 9722 8524 10202
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8392 8016 8444 8022
rect 8576 8016 8628 8022
rect 8392 7958 8444 7964
rect 8574 7984 8576 7993
rect 8628 7984 8630 7993
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 7852 7534 8064 7562
rect 7746 6896 7802 6905
rect 7656 6860 7708 6866
rect 7746 6831 7802 6840
rect 7656 6802 7708 6808
rect 7668 6118 7696 6802
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 5710 7696 6054
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7760 4826 7788 5238
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7576 4282 7604 4694
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7576 3738 7604 4082
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7576 3058 7604 3674
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7470 2680 7526 2689
rect 7470 2615 7472 2624
rect 7524 2615 7526 2624
rect 7472 2586 7524 2592
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6918 1456 6974 1465
rect 6644 1420 6696 1426
rect 6918 1391 6974 1400
rect 6644 1362 6696 1368
rect 6932 480 6960 1391
rect 7392 480 7420 2382
rect 7760 480 7788 4626
rect 7852 2514 7880 7534
rect 7930 7304 7986 7313
rect 7930 7239 7986 7248
rect 7944 7041 7972 7239
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 7930 7032 7986 7041
rect 7930 6967 7986 6976
rect 7944 5778 7972 6967
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7944 4826 7972 5714
rect 8022 5264 8078 5273
rect 8022 5199 8078 5208
rect 8036 5166 8064 5199
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7932 4820 7984 4826
rect 7984 4780 8156 4808
rect 7932 4762 7984 4768
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7944 2650 7972 3606
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7840 2508 7892 2514
rect 8128 2496 8156 4780
rect 8220 4146 8248 7142
rect 8312 6866 8340 7686
rect 8404 7478 8432 7958
rect 8574 7919 8630 7928
rect 8588 7546 8616 7919
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8404 6458 8432 7414
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8404 6254 8432 6394
rect 8392 6248 8444 6254
rect 8298 6216 8354 6225
rect 8392 6190 8444 6196
rect 8298 6151 8354 6160
rect 8312 5846 8340 6151
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8206 4040 8262 4049
rect 8312 4010 8340 5510
rect 8404 5098 8432 5646
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8404 4554 8432 5034
rect 8496 4690 8524 5102
rect 8680 4865 8708 14010
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9416 12238 9444 15302
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8864 6186 8892 8502
rect 9508 8480 9536 18022
rect 9692 17762 9720 18566
rect 9784 17882 9812 18686
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9600 17746 9720 17762
rect 9588 17740 9720 17746
rect 9640 17734 9720 17740
rect 9864 17740 9916 17746
rect 9588 17682 9640 17688
rect 9864 17682 9916 17688
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9784 17066 9812 17478
rect 9876 17202 9904 17682
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9692 15502 9720 16623
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9784 15434 9812 17002
rect 9968 16674 9996 19128
rect 10048 19110 10100 19116
rect 9876 16646 9996 16674
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9692 11762 9720 14486
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11506 9720 11562
rect 9600 11478 9720 11506
rect 9600 10033 9628 11478
rect 9784 10266 9812 14010
rect 9876 13954 9904 16646
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 16114 9996 16526
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9968 15570 9996 16050
rect 10060 15978 10088 19110
rect 10152 18154 10180 21678
rect 10336 21486 10364 21830
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10336 21078 10364 21422
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10336 20602 10364 21014
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10520 19174 10548 31418
rect 10598 30152 10654 30161
rect 10598 30087 10654 30096
rect 10612 29782 10640 30087
rect 10600 29776 10652 29782
rect 10600 29718 10652 29724
rect 10704 29594 10732 35430
rect 11164 35290 11192 35566
rect 11152 35284 11204 35290
rect 11072 35244 11152 35272
rect 10784 35148 10836 35154
rect 10784 35090 10836 35096
rect 10796 34406 10824 35090
rect 10784 34400 10836 34406
rect 10784 34342 10836 34348
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10980 33114 11008 33798
rect 10968 33108 11020 33114
rect 10968 33050 11020 33056
rect 10784 32972 10836 32978
rect 10784 32914 10836 32920
rect 10796 32570 10824 32914
rect 10784 32564 10836 32570
rect 10784 32506 10836 32512
rect 10796 31657 10824 32506
rect 10968 32360 11020 32366
rect 10968 32302 11020 32308
rect 10980 32065 11008 32302
rect 10966 32056 11022 32065
rect 10966 31991 11022 32000
rect 10782 31648 10838 31657
rect 10782 31583 10838 31592
rect 10796 31278 10824 31583
rect 11072 31278 11100 35244
rect 11152 35226 11204 35232
rect 11150 35048 11206 35057
rect 11150 34983 11206 34992
rect 11164 31958 11192 34983
rect 11244 34468 11296 34474
rect 11244 34410 11296 34416
rect 11152 31952 11204 31958
rect 11152 31894 11204 31900
rect 11256 31278 11284 34410
rect 11348 33153 11376 36654
rect 11532 35290 11560 39520
rect 11900 37754 11928 39520
rect 11900 37726 12020 37754
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11520 35284 11572 35290
rect 11520 35226 11572 35232
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 11428 33312 11480 33318
rect 11428 33254 11480 33260
rect 11334 33144 11390 33153
rect 11334 33079 11390 33088
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 11244 31272 11296 31278
rect 11244 31214 11296 31220
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 10784 30864 10836 30870
rect 10782 30832 10784 30841
rect 10836 30832 10838 30841
rect 10782 30767 10838 30776
rect 10888 29782 10916 31214
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11256 30870 11284 31078
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 10966 30288 11022 30297
rect 10966 30223 11022 30232
rect 10876 29776 10928 29782
rect 10612 29566 10732 29594
rect 10796 29736 10876 29764
rect 10612 25906 10640 29566
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10704 28218 10732 29446
rect 10796 29238 10824 29736
rect 10876 29718 10928 29724
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10888 29306 10916 29582
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10784 29232 10836 29238
rect 10784 29174 10836 29180
rect 10874 29200 10930 29209
rect 10980 29186 11008 30223
rect 11256 30190 11284 30534
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 10930 29158 11008 29186
rect 10874 29135 10930 29144
rect 10692 28212 10744 28218
rect 10692 28154 10744 28160
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10796 25362 10824 28154
rect 10784 25356 10836 25362
rect 10784 25298 10836 25304
rect 10796 24954 10824 25298
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 10782 24712 10838 24721
rect 10782 24647 10838 24656
rect 10600 23792 10652 23798
rect 10598 23760 10600 23769
rect 10652 23760 10654 23769
rect 10598 23695 10654 23704
rect 10612 23526 10640 23695
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 22234 10640 22918
rect 10704 22778 10732 23122
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10612 21554 10640 22170
rect 10704 22166 10732 22714
rect 10796 22506 10824 24647
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10692 22160 10744 22166
rect 10692 22102 10744 22108
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10612 19922 10640 20470
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19514 10640 19858
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10244 18426 10272 18838
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15162 9996 15506
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10060 14822 10088 15438
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9876 13926 9996 13954
rect 9864 13864 9916 13870
rect 9968 13841 9996 13926
rect 9864 13806 9916 13812
rect 9954 13832 10010 13841
rect 9876 13190 9904 13806
rect 9954 13767 10010 13776
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 12782 9904 13126
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 10060 12374 10088 14758
rect 10152 14550 10180 18090
rect 10336 17746 10364 18702
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10428 17882 10456 18022
rect 10612 17882 10640 18566
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10428 17513 10456 17818
rect 10612 17649 10640 17818
rect 10690 17776 10746 17785
rect 10690 17711 10746 17720
rect 10598 17640 10654 17649
rect 10598 17575 10654 17584
rect 10414 17504 10470 17513
rect 10414 17439 10470 17448
rect 10704 16998 10732 17711
rect 10796 17610 10824 19450
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10796 17066 10824 17546
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10152 14074 10180 14486
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10244 12866 10272 15914
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10428 14822 10456 15574
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10336 13802 10364 14350
rect 10428 14346 10456 14758
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10336 13530 10364 13738
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10336 12986 10364 13466
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10244 12838 10456 12866
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 11354 9996 12242
rect 10060 11558 10088 12310
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10152 11506 10180 11698
rect 10244 11626 10272 12174
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9586 10024 9642 10033
rect 9586 9959 9642 9968
rect 9784 9722 9812 10202
rect 9968 10130 9996 11290
rect 10060 10713 10088 11494
rect 10152 11478 10272 11506
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10742 10180 11154
rect 10140 10736 10192 10742
rect 10046 10704 10102 10713
rect 10140 10678 10192 10684
rect 10046 10639 10102 10648
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10244 10062 10272 11478
rect 10336 11150 10364 11181
rect 10324 11144 10376 11150
rect 10322 11112 10324 11121
rect 10376 11112 10378 11121
rect 10322 11047 10378 11056
rect 10336 10742 10364 11047
rect 10324 10736 10376 10742
rect 10428 10713 10456 12838
rect 10704 12356 10732 16934
rect 10796 16590 10824 17002
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10796 15910 10824 16526
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10888 14498 10916 29135
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11072 28778 11100 28902
rect 11256 28778 11284 30126
rect 11072 28750 11284 28778
rect 11072 28626 11100 28750
rect 11244 28688 11296 28694
rect 11244 28630 11296 28636
rect 11060 28620 11112 28626
rect 11060 28562 11112 28568
rect 11072 28218 11100 28562
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11256 28082 11284 28630
rect 11244 28076 11296 28082
rect 11244 28018 11296 28024
rect 11256 27674 11284 28018
rect 11244 27668 11296 27674
rect 11244 27610 11296 27616
rect 11348 27554 11376 31214
rect 11256 27526 11376 27554
rect 11060 25764 11112 25770
rect 11060 25706 11112 25712
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10980 25401 11008 25638
rect 10966 25392 11022 25401
rect 11072 25362 11100 25706
rect 10966 25327 11022 25336
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 11072 25158 11100 25298
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11072 24614 11100 25094
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11072 24410 11100 24550
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 10980 23338 11008 23734
rect 11072 23594 11100 24346
rect 11164 24274 11192 24890
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11164 23662 11192 24006
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10980 23310 11100 23338
rect 11164 23322 11192 23598
rect 11072 23118 11100 23310
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22778 11100 23054
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10980 21690 11008 22034
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 10980 21010 11008 21626
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10980 20534 11008 20946
rect 11072 20890 11100 22442
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 11164 21690 11192 22102
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11072 20862 11192 20890
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 11072 20097 11100 20742
rect 11058 20088 11114 20097
rect 11058 20023 11114 20032
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10980 19174 11008 19858
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 18630 11008 19110
rect 11164 18850 11192 20862
rect 11256 19224 11284 27526
rect 11336 26920 11388 26926
rect 11336 26862 11388 26868
rect 11348 19292 11376 26862
rect 11440 19961 11468 33254
rect 11532 26926 11560 34478
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11992 33658 12020 37726
rect 12268 36394 12296 39520
rect 12636 36938 12664 39520
rect 12360 36922 12664 36938
rect 12348 36916 12664 36922
rect 12400 36910 12664 36916
rect 12348 36858 12400 36864
rect 13096 36689 13124 39520
rect 13082 36680 13138 36689
rect 13082 36615 13138 36624
rect 12176 36366 12296 36394
rect 13464 36378 13492 39520
rect 13452 36372 13504 36378
rect 12072 35148 12124 35154
rect 12072 35090 12124 35096
rect 12084 34542 12112 35090
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11796 31952 11848 31958
rect 11796 31894 11848 31900
rect 11888 31952 11940 31958
rect 11888 31894 11940 31900
rect 11808 31278 11836 31894
rect 11900 31346 11928 31894
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11980 29708 12032 29714
rect 11980 29650 12032 29656
rect 11992 29034 12020 29650
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11992 26466 12020 28970
rect 11532 26438 12020 26466
rect 11532 20369 11560 26438
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 12084 24818 12112 34478
rect 12176 32570 12204 36366
rect 13452 36314 13504 36320
rect 12256 36236 12308 36242
rect 12256 36178 12308 36184
rect 12268 35494 12296 36178
rect 13832 35850 13860 39520
rect 13740 35834 13860 35850
rect 13728 35828 13860 35834
rect 13780 35822 13860 35828
rect 13728 35770 13780 35776
rect 12256 35488 12308 35494
rect 12256 35430 12308 35436
rect 13268 35488 13320 35494
rect 13268 35430 13320 35436
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 12164 31748 12216 31754
rect 12164 31690 12216 31696
rect 12176 31142 12204 31690
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 12176 30258 12204 31078
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12164 30116 12216 30122
rect 12164 30058 12216 30064
rect 12176 30025 12204 30058
rect 12162 30016 12218 30025
rect 12162 29951 12218 29960
rect 12268 29714 12296 35430
rect 13176 35148 13228 35154
rect 13176 35090 13228 35096
rect 13188 34542 13216 35090
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 12716 34060 12768 34066
rect 12716 34002 12768 34008
rect 12728 33318 12756 34002
rect 12716 33312 12768 33318
rect 12716 33254 12768 33260
rect 12440 31884 12492 31890
rect 12440 31826 12492 31832
rect 12452 31736 12480 31826
rect 12452 31708 12572 31736
rect 12438 31648 12494 31657
rect 12438 31583 12494 31592
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12360 30802 12388 31282
rect 12452 31278 12480 31583
rect 12544 31498 12572 31708
rect 12624 31680 12676 31686
rect 12622 31648 12624 31657
rect 12676 31648 12678 31657
rect 12622 31583 12678 31592
rect 12544 31482 12664 31498
rect 12544 31476 12676 31482
rect 12544 31470 12624 31476
rect 12624 31418 12676 31424
rect 12532 31408 12584 31414
rect 12530 31376 12532 31385
rect 12584 31376 12586 31385
rect 12530 31311 12586 31320
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12452 30938 12480 31214
rect 12440 30932 12492 30938
rect 12440 30874 12492 30880
rect 12348 30796 12400 30802
rect 12348 30738 12400 30744
rect 12360 30054 12388 30738
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12360 29646 12388 29990
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12360 28966 12388 29582
rect 12636 29306 12664 29786
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 12348 28960 12400 28966
rect 12348 28902 12400 28908
rect 12360 28762 12388 28902
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12438 28656 12494 28665
rect 12438 28591 12494 28600
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11796 24744 11848 24750
rect 11794 24712 11796 24721
rect 11848 24712 11850 24721
rect 11794 24647 11850 24656
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11796 24336 11848 24342
rect 11796 24278 11848 24284
rect 11808 23866 11836 24278
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11612 23248 11664 23254
rect 11612 23190 11664 23196
rect 11624 22642 11652 23190
rect 11992 23050 12020 24210
rect 11980 23044 12032 23050
rect 11980 22986 12032 22992
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11518 20360 11574 20369
rect 11518 20295 11574 20304
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11992 20058 12020 22986
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11348 19264 11560 19292
rect 11256 19196 11468 19224
rect 11072 18822 11192 18850
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10980 17338 11008 18362
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11072 16402 11100 18822
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11164 18426 11192 18634
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11440 17524 11468 19196
rect 11348 17496 11468 17524
rect 11072 16374 11192 16402
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15502 11100 15846
rect 11164 15609 11192 16374
rect 11150 15600 11206 15609
rect 11150 15535 11206 15544
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14822 11100 15438
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10520 12328 10732 12356
rect 10796 14470 10916 14498
rect 11072 14482 11100 14758
rect 11060 14476 11112 14482
rect 10324 10678 10376 10684
rect 10414 10704 10470 10713
rect 10414 10639 10470 10648
rect 10520 10588 10548 12328
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10612 11626 10640 12174
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11694 10732 12038
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10612 11218 10640 11562
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10336 10560 10548 10588
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9722 10272 9998
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9784 8922 9812 9658
rect 10152 9518 10180 9549
rect 10140 9512 10192 9518
rect 10138 9480 10140 9489
rect 10192 9480 10194 9489
rect 10138 9415 10194 9424
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 8945 9904 8978
rect 9416 8452 9536 8480
rect 9692 8894 9812 8922
rect 9862 8936 9918 8945
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8666 4856 8722 4865
rect 8666 4791 8722 4800
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8496 4282 8524 4626
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8680 4185 8708 4422
rect 8666 4176 8722 4185
rect 8666 4111 8722 4120
rect 8206 3975 8262 3984
rect 8300 4004 8352 4010
rect 8220 3738 8248 3975
rect 8300 3946 8352 3952
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8220 3194 8248 3674
rect 8680 3602 8708 3878
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8312 2650 8340 3538
rect 8574 3088 8630 3097
rect 8574 3023 8630 3032
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8300 2508 8352 2514
rect 8128 2468 8300 2496
rect 7840 2450 7892 2456
rect 8300 2450 8352 2456
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8220 480 8248 2314
rect 8588 480 8616 3023
rect 8772 2990 8800 6054
rect 8864 5914 8892 6122
rect 9048 5914 9076 6326
rect 9324 6254 9352 6802
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9416 4622 9444 8452
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 8090 9536 8298
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9600 7750 9628 8230
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7274 9628 7686
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9600 6254 9628 7210
rect 9588 6248 9640 6254
rect 9692 6225 9720 8894
rect 9862 8871 9918 8880
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9588 6190 9640 6196
rect 9678 6216 9734 6225
rect 9600 6100 9628 6190
rect 9678 6151 9734 6160
rect 9600 6072 9720 6100
rect 9692 4690 9720 6072
rect 9784 5846 9812 8774
rect 9876 8634 9904 8871
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9876 7478 9904 7958
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10060 7857 10088 7890
rect 10046 7848 10102 7857
rect 10046 7783 10102 7792
rect 9864 7472 9916 7478
rect 9862 7440 9864 7449
rect 9916 7440 9918 7449
rect 9862 7375 9918 7384
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 6798 9904 7278
rect 10060 7002 10088 7783
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9784 5370 9812 5782
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9876 4826 9904 5850
rect 9968 5692 9996 6122
rect 10060 5817 10088 6938
rect 10046 5808 10102 5817
rect 10046 5743 10102 5752
rect 9968 5664 10088 5692
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9324 4146 9352 4422
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8864 2922 8892 3674
rect 8956 3670 8984 3946
rect 9416 3670 9444 4014
rect 9600 3942 9628 4490
rect 9968 4321 9996 5238
rect 9954 4312 10010 4321
rect 9954 4247 10010 4256
rect 10060 4196 10088 5664
rect 9968 4168 10088 4196
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 9600 3194 9628 3878
rect 9692 3641 9720 3878
rect 9678 3632 9734 3641
rect 9678 3567 9734 3576
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 9324 2666 9352 2926
rect 9324 2638 9444 2666
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8944 1420 8996 1426
rect 8944 1362 8996 1368
rect 8956 480 8984 1362
rect 9416 480 9444 2638
rect 9784 480 9812 4014
rect 9968 2689 9996 4168
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3777 10088 3878
rect 10046 3768 10102 3777
rect 10046 3703 10102 3712
rect 10060 3670 10088 3703
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10152 3516 10180 9415
rect 10244 7041 10272 9658
rect 10336 9602 10364 10560
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10612 9722 10640 10066
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10336 9574 10456 9602
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8294 10364 8910
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10230 7032 10286 7041
rect 10230 6967 10286 6976
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6118 10272 6734
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5030 10272 6054
rect 10336 5846 10364 7142
rect 10428 6186 10456 9574
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10612 8294 10640 9046
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10520 6934 10548 7958
rect 10612 7818 10640 8230
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7342 10732 7686
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10520 6458 10548 6870
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 5098 10456 5510
rect 10520 5166 10548 5782
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10244 3534 10272 4966
rect 10428 4554 10456 5034
rect 10416 4548 10468 4554
rect 10416 4490 10468 4496
rect 10520 4264 10548 5102
rect 10612 4622 10640 5170
rect 10796 5080 10824 14470
rect 11060 14418 11112 14424
rect 11072 13326 11100 14418
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12782 11100 13262
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 9994 10916 11494
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10980 10810 11008 11222
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11072 10538 11100 11766
rect 11164 11098 11192 15535
rect 11348 12084 11376 17496
rect 11532 17241 11560 19264
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11518 17232 11574 17241
rect 11518 17167 11574 17176
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11440 16658 11468 17002
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 16250 11468 16594
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11440 14074 11468 16186
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15162 11560 15506
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11532 14822 11560 15098
rect 12084 14929 12112 24754
rect 12176 23186 12204 25094
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12346 24712 12402 24721
rect 12268 24274 12296 24686
rect 12346 24647 12348 24656
rect 12400 24647 12402 24656
rect 12348 24618 12400 24624
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12268 23254 12296 23734
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 16794 12204 17682
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12360 15065 12388 23598
rect 12452 23508 12480 28591
rect 12530 25392 12586 25401
rect 12530 25327 12586 25336
rect 12544 24954 12572 25327
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12728 24313 12756 33254
rect 12806 32872 12862 32881
rect 12806 32807 12862 32816
rect 12714 24304 12770 24313
rect 12714 24239 12770 24248
rect 12820 23662 12848 32807
rect 12900 31680 12952 31686
rect 12900 31622 12952 31628
rect 12912 31210 12940 31622
rect 12900 31204 12952 31210
rect 12900 31146 12952 31152
rect 13188 30297 13216 34478
rect 13174 30288 13230 30297
rect 13174 30223 13230 30232
rect 13280 25265 13308 35430
rect 13358 35320 13414 35329
rect 13358 35255 13360 35264
rect 13412 35255 13414 35264
rect 13360 35226 13412 35232
rect 13634 35048 13690 35057
rect 13634 34983 13690 34992
rect 13648 34746 13676 34983
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 14200 34202 14228 39520
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14660 35329 14688 39520
rect 14646 35320 14702 35329
rect 14646 35255 14702 35264
rect 15028 35057 15056 39520
rect 15014 35048 15070 35057
rect 15014 34983 15070 34992
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14188 34196 14240 34202
rect 14188 34138 14240 34144
rect 15396 33969 15424 39520
rect 13634 33960 13690 33969
rect 13634 33895 13690 33904
rect 15382 33960 15438 33969
rect 15382 33895 15438 33904
rect 13648 33658 13676 33895
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13452 33448 13504 33454
rect 13452 33390 13504 33396
rect 13464 32881 13492 33390
rect 13450 32872 13506 32881
rect 13450 32807 13506 32816
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 15764 26926 15792 39520
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 15752 26920 15804 26926
rect 15752 26862 15804 26868
rect 13266 25256 13322 25265
rect 13266 25191 13322 25200
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 24750 13124 25094
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13096 23730 13124 24346
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12532 23520 12584 23526
rect 12452 23480 12532 23508
rect 12452 23322 12480 23480
rect 12532 23462 12584 23468
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12346 15056 12402 15065
rect 12346 14991 12402 15000
rect 12070 14920 12126 14929
rect 12070 14855 12126 14864
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 12346 14648 12402 14657
rect 12346 14583 12402 14592
rect 12360 14550 12388 14583
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 12084 14006 12112 14418
rect 12360 14074 12388 14486
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 12452 13546 12480 15302
rect 12360 13518 12480 13546
rect 12360 13462 12388 13518
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 11532 12986 11560 13398
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11532 12238 11560 12922
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11348 12056 11560 12084
rect 11164 11070 11468 11098
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10198 11100 10474
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10876 9988 10928 9994
rect 10876 9930 10928 9936
rect 11164 9178 11192 10678
rect 11256 10674 11284 10950
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11348 10266 11376 10610
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11334 10160 11390 10169
rect 11334 10095 11390 10104
rect 11348 10062 11376 10095
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9722 11376 9998
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11440 9194 11468 11070
rect 11532 10248 11560 12056
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 10810 12388 11222
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12360 10577 12388 10746
rect 12452 10674 12480 13126
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12346 10568 12402 10577
rect 12346 10503 12402 10512
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11532 10220 11652 10248
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11532 9722 11560 9862
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11624 9466 11652 10220
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 11808 9654 11836 10134
rect 12176 9654 12204 10134
rect 12452 10130 12480 10610
rect 12544 10146 12572 23462
rect 13096 23322 13124 23666
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12714 17504 12770 17513
rect 12714 17439 12770 17448
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 14618 12664 14758
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12636 12238 12664 14554
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 11286 12664 12174
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12636 11150 12664 11222
rect 12728 11218 12756 17439
rect 13832 14657 13860 26862
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 13818 14648 13874 14657
rect 13818 14583 13874 14592
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12820 10606 12848 11494
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12716 10464 12768 10470
rect 12912 10418 12940 11154
rect 13096 11014 13124 11290
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10674 13124 10950
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12716 10406 12768 10412
rect 12440 10124 12492 10130
rect 12544 10118 12664 10146
rect 12440 10066 12492 10072
rect 12452 9654 12480 10066
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 11796 9648 11848 9654
rect 11794 9616 11796 9625
rect 12164 9648 12216 9654
rect 11848 9616 11850 9625
rect 12164 9590 12216 9596
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 11794 9551 11850 9560
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11348 9166 11468 9194
rect 11532 9438 11652 9466
rect 11164 8634 11192 9114
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10704 5052 10824 5080
rect 10704 4758 10732 5052
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10428 4236 10548 4264
rect 10428 3670 10456 4236
rect 10506 4176 10562 4185
rect 10506 4111 10562 4120
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10060 3488 10180 3516
rect 10232 3528 10284 3534
rect 9954 2680 10010 2689
rect 10060 2650 10088 3488
rect 10232 3470 10284 3476
rect 10138 3224 10194 3233
rect 10138 3159 10194 3168
rect 9954 2615 10010 2624
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10152 480 10180 3159
rect 10244 2854 10272 3470
rect 10428 3194 10456 3606
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10520 1442 10548 4111
rect 10612 2378 10640 4558
rect 10704 4282 10732 4694
rect 10692 4276 10744 4282
rect 10744 4236 10824 4264
rect 10692 4218 10744 4224
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10704 3641 10732 3878
rect 10690 3632 10746 3641
rect 10690 3567 10746 3576
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10796 1465 10824 4236
rect 10888 3126 10916 5578
rect 11150 5128 11206 5137
rect 11150 5063 11206 5072
rect 10966 4856 11022 4865
rect 11164 4826 11192 5063
rect 10966 4791 10968 4800
rect 11020 4791 11022 4800
rect 11152 4820 11204 4826
rect 10968 4762 11020 4768
rect 11152 4762 11204 4768
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4146 11100 4422
rect 11164 4146 11192 4762
rect 11256 4622 11284 6598
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10966 2952 11022 2961
rect 10966 2887 11022 2896
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10888 2417 10916 2450
rect 10874 2408 10930 2417
rect 10874 2343 10930 2352
rect 10782 1456 10838 1465
rect 10520 1414 10640 1442
rect 10612 480 10640 1414
rect 10782 1391 10838 1400
rect 10980 480 11008 2887
rect 11256 2836 11284 4558
rect 11348 2990 11376 9166
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8090 11468 8978
rect 11532 8650 11560 9438
rect 12268 9330 12296 9590
rect 12176 9302 12296 9330
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11532 8622 11652 8650
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11440 7177 11468 7210
rect 11426 7168 11482 7177
rect 11426 7103 11482 7112
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11440 5030 11468 5646
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11532 3641 11560 8502
rect 11624 8430 11652 8622
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7342 11836 7822
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11992 4808 12020 8366
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11900 4780 12020 4808
rect 11900 4049 11928 4780
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11992 4282 12020 4626
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11518 3632 11574 3641
rect 11518 3567 11574 3576
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11520 2848 11572 2854
rect 11256 2808 11376 2836
rect 11348 2650 11376 2808
rect 12084 2825 12112 6054
rect 12176 5846 12204 9302
rect 12544 9194 12572 9930
rect 12268 9166 12572 9194
rect 12268 9042 12296 9166
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12360 8294 12388 9046
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12360 7954 12388 8230
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12360 7206 12388 7890
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12360 6882 12388 7142
rect 12360 6854 12480 6882
rect 12452 6338 12480 6854
rect 12636 6458 12664 10118
rect 12728 9926 12756 10406
rect 12820 10390 12940 10418
rect 12820 9926 12848 10390
rect 13096 10198 13124 10610
rect 13372 10198 13400 10678
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13360 10192 13412 10198
rect 13544 10192 13596 10198
rect 13412 10152 13492 10180
rect 13360 10134 13412 10140
rect 13174 10024 13230 10033
rect 13174 9959 13230 9968
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12728 8401 12756 9862
rect 12714 8392 12770 8401
rect 12714 8327 12770 8336
rect 12820 7188 12848 9862
rect 12990 9480 13046 9489
rect 12990 9415 13046 9424
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8634 12940 8978
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12728 7160 12848 7188
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12452 6310 12664 6338
rect 12636 5914 12664 6310
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12622 5808 12678 5817
rect 12176 5370 12204 5782
rect 12622 5743 12678 5752
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12440 5160 12492 5166
rect 12438 5128 12440 5137
rect 12492 5128 12494 5137
rect 12438 5063 12494 5072
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 11520 2790 11572 2796
rect 12070 2816 12126 2825
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11334 1456 11390 1465
rect 11532 1442 11560 2790
rect 11622 2748 11918 2768
rect 12070 2751 12126 2760
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11532 1414 11836 1442
rect 11334 1391 11390 1400
rect 11348 480 11376 1391
rect 11808 480 11836 1414
rect 12268 626 12296 4422
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12452 3534 12480 4014
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12438 3088 12494 3097
rect 12438 3023 12494 3032
rect 12452 2990 12480 3023
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12176 598 12296 626
rect 12176 480 12204 598
rect 12544 480 12572 4966
rect 12636 4078 12664 5743
rect 12728 4690 12756 7160
rect 12806 6896 12862 6905
rect 12806 6831 12808 6840
rect 12860 6831 12862 6840
rect 12808 6802 12860 6808
rect 12820 6458 12848 6802
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 13004 6202 13032 9415
rect 13188 9110 13216 9959
rect 13464 9178 13492 10152
rect 13544 10134 13596 10140
rect 13556 9722 13584 10134
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13084 8424 13136 8430
rect 13082 8392 13084 8401
rect 13136 8392 13138 8401
rect 13082 8327 13138 8336
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13004 6174 13124 6202
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3233 12664 3878
rect 12622 3224 12678 3233
rect 12622 3159 12678 3168
rect 12622 2952 12678 2961
rect 12622 2887 12678 2896
rect 12636 2854 12664 2887
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12622 2544 12678 2553
rect 12622 2479 12624 2488
rect 12676 2479 12678 2488
rect 12624 2450 12676 2456
rect 12728 2417 12756 3946
rect 12806 3496 12862 3505
rect 12806 3431 12808 3440
rect 12860 3431 12862 3440
rect 12808 3402 12860 3408
rect 12714 2408 12770 2417
rect 12714 2343 12770 2352
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 1465 12848 2246
rect 12806 1456 12862 1465
rect 12806 1391 12862 1400
rect 13004 480 13032 6054
rect 13096 4690 13124 6174
rect 13084 4684 13136 4690
rect 13136 4644 13216 4672
rect 13084 4626 13136 4632
rect 13082 4312 13138 4321
rect 13188 4282 13216 4644
rect 13082 4247 13138 4256
rect 13176 4276 13228 4282
rect 13096 3602 13124 4247
rect 13176 4218 13228 4224
rect 13280 3913 13308 8230
rect 13556 4049 13584 9318
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13542 4040 13598 4049
rect 13542 3975 13598 3984
rect 13266 3904 13322 3913
rect 13266 3839 13322 3848
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13096 3126 13124 3538
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13280 3058 13308 3606
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13372 3194 13400 3538
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13358 2816 13414 2825
rect 13358 2751 13414 2760
rect 13372 480 13400 2751
rect 13740 480 13768 6598
rect 14200 480 14228 7142
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 15750 4584 15806 4593
rect 15750 4519 15806 4528
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14922 4040 14978 4049
rect 14922 3975 14978 3984
rect 14646 3904 14702 3913
rect 14646 3839 14702 3848
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 3839
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 3975
rect 15382 3632 15438 3641
rect 15382 3567 15438 3576
rect 15396 480 15424 3567
rect 15764 480 15792 4519
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 202 34720 258 34776
rect 570 33360 626 33416
rect 938 32816 994 32872
rect 1582 36352 1638 36408
rect 1582 34040 1638 34096
rect 1766 33088 1822 33144
rect 1398 32308 1400 32328
rect 1400 32308 1452 32328
rect 1452 32308 1454 32328
rect 1398 32272 1454 32308
rect 2778 38664 2834 38720
rect 1306 31320 1362 31376
rect 1674 31592 1730 31648
rect 1674 30676 1676 30696
rect 1676 30676 1728 30696
rect 1728 30676 1730 30696
rect 1674 30640 1730 30676
rect 2778 32816 2834 32872
rect 3146 34604 3202 34640
rect 3146 34584 3148 34604
rect 3148 34584 3200 34604
rect 3200 34584 3202 34604
rect 3238 32952 3294 33008
rect 3054 30096 3110 30152
rect 1674 29280 1730 29336
rect 1674 27820 1676 27840
rect 1676 27820 1728 27840
rect 1728 27820 1730 27840
rect 1674 27784 1730 27820
rect 1582 26968 1638 27024
rect 2226 26288 2282 26344
rect 2594 25644 2596 25664
rect 2596 25644 2648 25664
rect 2648 25644 2650 25664
rect 2594 25608 2650 25644
rect 1674 24520 1730 24576
rect 2962 25744 3018 25800
rect 1674 22208 1730 22264
rect 1398 21004 1454 21040
rect 1398 20984 1400 21004
rect 1400 20984 1452 21004
rect 1452 20984 1454 21004
rect 1398 16088 1454 16144
rect 1674 19896 1730 19952
rect 1582 17584 1638 17640
rect 2226 20460 2282 20496
rect 2226 20440 2228 20460
rect 2228 20440 2280 20460
rect 2280 20440 2282 20460
rect 2134 16904 2190 16960
rect 1674 15136 1730 15192
rect 1582 12824 1638 12880
rect 1398 11736 1454 11792
rect 1582 10512 1638 10568
rect 2226 13932 2282 13968
rect 2226 13912 2228 13932
rect 2228 13912 2280 13932
rect 2280 13912 2282 13932
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3422 34720 3478 34776
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 4434 35536 4490 35592
rect 4802 34720 4858 34776
rect 4618 33108 4674 33144
rect 4618 33088 4620 33108
rect 4620 33088 4672 33108
rect 4672 33088 4674 33108
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3422 24656 3478 24712
rect 3146 23704 3202 23760
rect 2962 23024 3018 23080
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 2502 10512 2558 10568
rect 2318 9424 2374 9480
rect 2134 8472 2190 8528
rect 1582 8064 1638 8120
rect 938 3576 994 3632
rect 1582 3440 1638 3496
rect 2686 12180 2688 12200
rect 2688 12180 2740 12200
rect 2740 12180 2742 12200
rect 2686 12144 2742 12180
rect 2594 9696 2650 9752
rect 2686 9560 2742 9616
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3882 20324 3938 20360
rect 3882 20304 3884 20324
rect 3884 20304 3936 20324
rect 3936 20304 3938 20324
rect 4894 32444 4896 32464
rect 4896 32444 4948 32464
rect 4948 32444 4950 32464
rect 4894 32408 4950 32444
rect 5262 32272 5318 32328
rect 5170 29144 5226 29200
rect 5630 35128 5686 35184
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6642 34584 6698 34640
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 5814 31728 5870 31784
rect 5722 30096 5778 30152
rect 4526 26968 4582 27024
rect 4342 26308 4398 26344
rect 4342 26288 4344 26308
rect 4344 26288 4396 26308
rect 4396 26288 4398 26308
rect 4342 25608 4398 25664
rect 4158 23568 4214 23624
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3238 19352 3294 19408
rect 3974 19352 4030 19408
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 5262 28056 5318 28112
rect 4618 25236 4620 25256
rect 4620 25236 4672 25256
rect 4672 25236 4674 25256
rect 4618 25200 4674 25236
rect 4434 19216 4490 19272
rect 4618 22480 4674 22536
rect 4894 23568 4950 23624
rect 4526 17720 4582 17776
rect 4618 17176 4674 17232
rect 5538 27784 5594 27840
rect 5354 27532 5410 27568
rect 5354 27512 5356 27532
rect 5356 27512 5408 27532
rect 5408 27512 5410 27532
rect 7194 34992 7250 35048
rect 8114 35536 8170 35592
rect 7930 35128 7986 35184
rect 7838 34740 7894 34776
rect 7838 34720 7840 34740
rect 7840 34720 7892 34740
rect 7892 34720 7894 34740
rect 7562 33224 7618 33280
rect 7194 32000 7250 32056
rect 6826 31728 6882 31784
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 5906 24248 5962 24304
rect 4434 16904 4490 16960
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 4066 15952 4122 16008
rect 3606 15580 3608 15600
rect 3608 15580 3660 15600
rect 3660 15580 3662 15600
rect 3606 15544 3662 15580
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3422 14864 3478 14920
rect 3606 14864 3662 14920
rect 3054 12860 3056 12880
rect 3056 12860 3108 12880
rect 3108 12860 3110 12880
rect 3054 12824 3110 12860
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3146 9968 3202 10024
rect 2318 7384 2374 7440
rect 1674 3304 1730 3360
rect 1490 1128 1546 1184
rect 2410 4972 2412 4992
rect 2412 4972 2464 4992
rect 2464 4972 2466 4992
rect 2410 4936 2466 4972
rect 2502 4528 2558 4584
rect 3054 7928 3110 7984
rect 2778 5752 2834 5808
rect 2962 5616 3018 5672
rect 2686 4664 2742 4720
rect 2870 3984 2926 4040
rect 2962 3476 2964 3496
rect 2964 3476 3016 3496
rect 3016 3476 3018 3496
rect 2962 3440 3018 3476
rect 3790 13796 3846 13832
rect 3790 13776 3792 13796
rect 3792 13776 3844 13796
rect 3844 13776 3846 13796
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 4342 10648 4398 10704
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3790 9424 3846 9480
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 4342 9152 4398 9208
rect 4066 7792 4122 7848
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 4158 4936 4214 4992
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3422 2760 3478 2816
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 4526 11736 4582 11792
rect 5078 17040 5134 17096
rect 5078 15952 5134 16008
rect 5354 15136 5410 15192
rect 5354 12824 5410 12880
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6734 27376 6790 27432
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 5722 20984 5778 21040
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 5722 16632 5778 16688
rect 5722 15136 5778 15192
rect 5814 15000 5870 15056
rect 4710 8608 4766 8664
rect 4618 6840 4674 6896
rect 4526 5344 4582 5400
rect 4434 5208 4490 5264
rect 4434 4664 4490 4720
rect 4526 4528 4582 4584
rect 4250 3032 4306 3088
rect 4802 7248 4858 7304
rect 5262 10104 5318 10160
rect 5078 9016 5134 9072
rect 5722 13640 5778 13696
rect 5630 11056 5686 11112
rect 5630 10104 5686 10160
rect 5630 9968 5686 10024
rect 5354 8608 5410 8664
rect 5354 5480 5410 5536
rect 4894 3848 4950 3904
rect 4802 3168 4858 3224
rect 5262 3984 5318 4040
rect 6182 20304 6238 20360
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6642 15136 6698 15192
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 5998 10104 6054 10160
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 5998 3848 6054 3904
rect 5538 2644 5594 2680
rect 5538 2624 5540 2644
rect 5540 2624 5592 2644
rect 5592 2624 5594 2644
rect 6090 2488 6146 2544
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 7378 31356 7380 31376
rect 7380 31356 7432 31376
rect 7432 31356 7434 31376
rect 7378 31320 7434 31356
rect 8114 32852 8116 32872
rect 8116 32852 8168 32872
rect 8168 32852 8170 32872
rect 8114 32816 8170 32852
rect 8482 34620 8484 34640
rect 8484 34620 8536 34640
rect 8536 34620 8538 34640
rect 8482 34584 8538 34620
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 7930 30776 7986 30832
rect 7102 29008 7158 29064
rect 7378 29144 7434 29200
rect 7378 28600 7434 28656
rect 7562 29164 7618 29200
rect 7562 29144 7564 29164
rect 7564 29144 7616 29164
rect 7616 29144 7618 29164
rect 7562 29008 7618 29064
rect 7286 27376 7342 27432
rect 6826 25744 6882 25800
rect 6826 23432 6882 23488
rect 7654 28056 7710 28112
rect 7562 26560 7618 26616
rect 7470 25916 7472 25936
rect 7472 25916 7524 25936
rect 7524 25916 7526 25936
rect 7470 25880 7526 25916
rect 7562 23740 7564 23760
rect 7564 23740 7616 23760
rect 7616 23740 7618 23760
rect 7562 23704 7618 23740
rect 8022 26696 8078 26752
rect 8298 27532 8354 27568
rect 8298 27512 8300 27532
rect 8300 27512 8352 27532
rect 8352 27512 8354 27532
rect 8022 25492 8078 25528
rect 8022 25472 8024 25492
rect 8024 25472 8076 25492
rect 8076 25472 8078 25492
rect 7930 23024 7986 23080
rect 7838 22480 7894 22536
rect 8114 24792 8170 24848
rect 8114 22480 8170 22536
rect 7102 19352 7158 19408
rect 6918 16088 6974 16144
rect 7010 13948 7012 13968
rect 7012 13948 7064 13968
rect 7064 13948 7066 13968
rect 7010 13912 7066 13948
rect 7562 20168 7618 20224
rect 7010 9016 7066 9072
rect 7378 11464 7434 11520
rect 7930 19896 7986 19952
rect 7286 9560 7342 9616
rect 7194 9424 7250 9480
rect 7562 11464 7618 11520
rect 7470 8880 7526 8936
rect 7378 8356 7434 8392
rect 7378 8336 7380 8356
rect 7380 8336 7432 8356
rect 7432 8336 7434 8356
rect 7194 7928 7250 7984
rect 7194 7112 7250 7168
rect 6734 5480 6790 5536
rect 6918 5616 6974 5672
rect 7010 5364 7066 5400
rect 7010 5344 7012 5364
rect 7012 5344 7064 5364
rect 7064 5344 7066 5364
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6826 3712 6882 3768
rect 7470 6840 7526 6896
rect 7102 4528 7158 4584
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9402 33360 9458 33416
rect 9310 33224 9366 33280
rect 8298 25472 8354 25528
rect 8574 24792 8630 24848
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8758 23704 8814 23760
rect 8390 23568 8446 23624
rect 8390 23024 8446 23080
rect 8298 17040 8354 17096
rect 8022 16632 8078 16688
rect 8022 13640 8078 13696
rect 7838 8492 7894 8528
rect 7838 8472 7840 8492
rect 7840 8472 7892 8492
rect 7892 8472 7894 8492
rect 8666 17620 8668 17640
rect 8668 17620 8720 17640
rect 8720 17620 8722 17640
rect 8666 17584 8722 17620
rect 8574 15000 8630 15056
rect 9586 33088 9642 33144
rect 9770 32952 9826 33008
rect 9586 32408 9642 32464
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 9126 25916 9128 25936
rect 9128 25916 9180 25936
rect 9180 25916 9182 25936
rect 9126 25880 9182 25916
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 9402 25472 9458 25528
rect 10966 36624 11022 36680
rect 10138 34584 10194 34640
rect 9770 30640 9826 30696
rect 9954 30096 10010 30152
rect 10322 32952 10378 33008
rect 10230 31320 10286 31376
rect 9862 27376 9918 27432
rect 10046 27004 10048 27024
rect 10048 27004 10100 27024
rect 10100 27004 10102 27024
rect 10046 26968 10102 27004
rect 10138 26832 10194 26888
rect 10138 26696 10194 26752
rect 9586 23840 9642 23896
rect 9586 23704 9642 23760
rect 9862 23432 9918 23488
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 9218 19216 9274 19272
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 9494 22752 9550 22808
rect 9402 20052 9458 20088
rect 9402 20032 9404 20052
rect 9404 20032 9456 20052
rect 9456 20032 9458 20052
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 9770 20440 9826 20496
rect 10138 22500 10194 22536
rect 10138 22480 10140 22500
rect 10140 22480 10192 22500
rect 10192 22480 10194 22500
rect 10414 28056 10470 28112
rect 9954 20032 10010 20088
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8390 12144 8446 12200
rect 8206 8628 8262 8664
rect 8206 8608 8208 8628
rect 8208 8608 8260 8628
rect 8260 8608 8262 8628
rect 8574 7964 8576 7984
rect 8576 7964 8628 7984
rect 8628 7964 8630 7984
rect 7746 6840 7802 6896
rect 7470 2644 7526 2680
rect 7470 2624 7472 2644
rect 7472 2624 7524 2644
rect 7524 2624 7526 2644
rect 6918 1400 6974 1456
rect 7930 7248 7986 7304
rect 7930 6976 7986 7032
rect 8022 5208 8078 5264
rect 8574 7928 8630 7964
rect 8298 6160 8354 6216
rect 8206 3984 8262 4040
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 9678 16632 9734 16688
rect 10598 30096 10654 30152
rect 10966 32000 11022 32056
rect 10782 31592 10838 31648
rect 11150 34992 11206 35048
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11334 33088 11390 33144
rect 10782 30812 10784 30832
rect 10784 30812 10836 30832
rect 10836 30812 10838 30832
rect 10782 30776 10838 30812
rect 10966 30232 11022 30288
rect 10874 29144 10930 29200
rect 10782 24656 10838 24712
rect 10598 23740 10600 23760
rect 10600 23740 10652 23760
rect 10652 23740 10654 23760
rect 10598 23704 10654 23740
rect 9954 13776 10010 13832
rect 10690 17720 10746 17776
rect 10598 17584 10654 17640
rect 10414 17448 10470 17504
rect 9586 9968 9642 10024
rect 10046 10648 10102 10704
rect 10322 11092 10324 11112
rect 10324 11092 10376 11112
rect 10376 11092 10378 11112
rect 10322 11056 10378 11092
rect 10966 25336 11022 25392
rect 11058 20032 11114 20088
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 13082 36624 13138 36680
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 12162 29960 12218 30016
rect 12438 31592 12494 31648
rect 12622 31628 12624 31648
rect 12624 31628 12676 31648
rect 12676 31628 12678 31648
rect 12622 31592 12678 31628
rect 12530 31356 12532 31376
rect 12532 31356 12584 31376
rect 12584 31356 12586 31376
rect 12530 31320 12586 31356
rect 12438 28600 12494 28656
rect 11794 24692 11796 24712
rect 11796 24692 11848 24712
rect 11848 24692 11850 24712
rect 11794 24656 11850 24692
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11518 20304 11574 20360
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11426 19896 11482 19952
rect 11150 15544 11206 15600
rect 10414 10648 10470 10704
rect 10138 9460 10140 9480
rect 10140 9460 10192 9480
rect 10192 9460 10194 9480
rect 10138 9424 10194 9460
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8666 4800 8722 4856
rect 8666 4120 8722 4176
rect 8574 3032 8630 3088
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 9862 8880 9918 8936
rect 9678 6160 9734 6216
rect 10046 7792 10102 7848
rect 9862 7420 9864 7440
rect 9864 7420 9916 7440
rect 9916 7420 9918 7440
rect 9862 7384 9918 7420
rect 10046 5752 10102 5808
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 9954 4256 10010 4312
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9678 3576 9734 3632
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10046 3712 10102 3768
rect 10230 6976 10286 7032
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11518 17176 11574 17232
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 12346 24676 12402 24712
rect 12346 24656 12348 24676
rect 12348 24656 12400 24676
rect 12400 24656 12402 24676
rect 12530 25336 12586 25392
rect 12806 32816 12862 32872
rect 12714 24248 12770 24304
rect 13174 30232 13230 30288
rect 13358 35284 13414 35320
rect 13358 35264 13360 35284
rect 13360 35264 13412 35284
rect 13412 35264 13414 35284
rect 13634 34992 13690 35048
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14646 35264 14702 35320
rect 15014 34992 15070 35048
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 13634 33904 13690 33960
rect 15382 33904 15438 33960
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 13450 32816 13506 32872
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 13266 25200 13322 25256
rect 12346 15000 12402 15056
rect 12070 14864 12126 14920
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 12346 14592 12402 14648
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11334 10104 11390 10160
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 12346 10512 12402 10568
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 12714 17448 12770 17504
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 13818 14592 13874 14648
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 11794 9596 11796 9616
rect 11796 9596 11848 9616
rect 11848 9596 11850 9616
rect 11794 9560 11850 9596
rect 10506 4120 10562 4176
rect 9954 2624 10010 2680
rect 10138 3168 10194 3224
rect 10690 3576 10746 3632
rect 11150 5072 11206 5128
rect 10966 4820 11022 4856
rect 10966 4800 10968 4820
rect 10968 4800 11020 4820
rect 11020 4800 11022 4820
rect 10966 2896 11022 2952
rect 10874 2352 10930 2408
rect 10782 1400 10838 1456
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11426 7112 11482 7168
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11886 3984 11942 4040
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11518 3576 11574 3632
rect 13174 9968 13230 10024
rect 12714 8336 12770 8392
rect 12990 9424 13046 9480
rect 12622 5752 12678 5808
rect 12438 5108 12440 5128
rect 12440 5108 12492 5128
rect 12492 5108 12494 5128
rect 12438 5072 12494 5108
rect 11334 1400 11390 1456
rect 12070 2760 12126 2816
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12438 3032 12494 3088
rect 12806 6860 12862 6896
rect 12806 6840 12808 6860
rect 12808 6840 12860 6860
rect 12860 6840 12862 6860
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 13082 8372 13084 8392
rect 13084 8372 13136 8392
rect 13136 8372 13138 8392
rect 13082 8336 13138 8372
rect 12622 3168 12678 3224
rect 12622 2896 12678 2952
rect 12622 2508 12678 2544
rect 12622 2488 12624 2508
rect 12624 2488 12676 2508
rect 12676 2488 12678 2508
rect 12806 3460 12862 3496
rect 12806 3440 12808 3460
rect 12808 3440 12860 3460
rect 12860 3440 12862 3460
rect 12714 2352 12770 2408
rect 12806 1400 12862 1456
rect 13082 4256 13138 4312
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 13542 3984 13598 4040
rect 13266 3848 13322 3904
rect 13358 2760 13414 2816
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 15750 4528 15806 4584
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14922 3984 14978 4040
rect 14646 3848 14702 3904
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 15382 3576 15438 3632
<< metal3 >>
rect 0 38722 480 38752
rect 2773 38722 2839 38725
rect 0 38720 2839 38722
rect 0 38664 2778 38720
rect 2834 38664 2839 38720
rect 0 38662 2839 38664
rect 0 38632 480 38662
rect 2773 38659 2839 38662
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 10961 36682 11027 36685
rect 13077 36682 13143 36685
rect 10961 36680 13143 36682
rect 10961 36624 10966 36680
rect 11022 36624 13082 36680
rect 13138 36624 13143 36680
rect 10961 36622 13143 36624
rect 10961 36619 11027 36622
rect 13077 36619 13143 36622
rect 6277 36480 6597 36481
rect 0 36410 480 36440
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 1577 36410 1643 36413
rect 0 36408 1643 36410
rect 0 36352 1582 36408
rect 1638 36352 1643 36408
rect 0 36350 1643 36352
rect 0 36320 480 36350
rect 1577 36347 1643 36350
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 4429 35594 4495 35597
rect 8109 35594 8175 35597
rect 4429 35592 8175 35594
rect 4429 35536 4434 35592
rect 4490 35536 8114 35592
rect 8170 35536 8175 35592
rect 4429 35534 8175 35536
rect 4429 35531 4495 35534
rect 8109 35531 8175 35534
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 13353 35322 13419 35325
rect 14641 35322 14707 35325
rect 13353 35320 14707 35322
rect 13353 35264 13358 35320
rect 13414 35264 14646 35320
rect 14702 35264 14707 35320
rect 13353 35262 14707 35264
rect 13353 35259 13419 35262
rect 14641 35259 14707 35262
rect 5625 35186 5691 35189
rect 7925 35186 7991 35189
rect 5625 35184 7991 35186
rect 5625 35128 5630 35184
rect 5686 35128 7930 35184
rect 7986 35128 7991 35184
rect 5625 35126 7991 35128
rect 5625 35123 5691 35126
rect 7925 35123 7991 35126
rect 7189 35050 7255 35053
rect 11145 35050 11211 35053
rect 7189 35048 11211 35050
rect 7189 34992 7194 35048
rect 7250 34992 11150 35048
rect 11206 34992 11211 35048
rect 7189 34990 11211 34992
rect 7189 34987 7255 34990
rect 11145 34987 11211 34990
rect 13629 35050 13695 35053
rect 15009 35050 15075 35053
rect 13629 35048 15075 35050
rect 13629 34992 13634 35048
rect 13690 34992 15014 35048
rect 15070 34992 15075 35048
rect 13629 34990 15075 34992
rect 13629 34987 13695 34990
rect 15009 34987 15075 34990
rect 4110 34854 8770 34914
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 197 34778 263 34781
rect 3417 34778 3483 34781
rect 197 34776 3483 34778
rect 197 34720 202 34776
rect 258 34720 3422 34776
rect 3478 34720 3483 34776
rect 197 34718 3483 34720
rect 197 34715 263 34718
rect 3417 34715 3483 34718
rect 3141 34642 3207 34645
rect 4110 34642 4170 34854
rect 4797 34778 4863 34781
rect 7833 34778 7899 34781
rect 4797 34776 7899 34778
rect 4797 34720 4802 34776
rect 4858 34720 7838 34776
rect 7894 34720 7899 34776
rect 4797 34718 7899 34720
rect 4797 34715 4863 34718
rect 7833 34715 7899 34718
rect 3141 34640 4170 34642
rect 3141 34584 3146 34640
rect 3202 34584 4170 34640
rect 3141 34582 4170 34584
rect 6637 34642 6703 34645
rect 8477 34642 8543 34645
rect 6637 34640 8543 34642
rect 6637 34584 6642 34640
rect 6698 34584 8482 34640
rect 8538 34584 8543 34640
rect 6637 34582 8543 34584
rect 8710 34642 8770 34854
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 10133 34642 10199 34645
rect 8710 34640 10199 34642
rect 8710 34584 10138 34640
rect 10194 34584 10199 34640
rect 8710 34582 10199 34584
rect 3141 34579 3207 34582
rect 6637 34579 6703 34582
rect 8477 34579 8543 34582
rect 10133 34579 10199 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 0 34098 480 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 480 34038
rect 1577 34035 1643 34038
rect 13629 33962 13695 33965
rect 15377 33962 15443 33965
rect 13629 33960 15443 33962
rect 13629 33904 13634 33960
rect 13690 33904 15382 33960
rect 15438 33904 15443 33960
rect 13629 33902 15443 33904
rect 13629 33899 13695 33902
rect 15377 33899 15443 33902
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 565 33418 631 33421
rect 9397 33418 9463 33421
rect 565 33416 9463 33418
rect 565 33360 570 33416
rect 626 33360 9402 33416
rect 9458 33360 9463 33416
rect 565 33358 9463 33360
rect 565 33355 631 33358
rect 9397 33355 9463 33358
rect 7557 33282 7623 33285
rect 9305 33282 9371 33285
rect 7557 33280 9371 33282
rect 7557 33224 7562 33280
rect 7618 33224 9310 33280
rect 9366 33224 9371 33280
rect 7557 33222 9371 33224
rect 7557 33219 7623 33222
rect 9305 33219 9371 33222
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 1761 33146 1827 33149
rect 4613 33146 4679 33149
rect 1761 33144 4679 33146
rect 1761 33088 1766 33144
rect 1822 33088 4618 33144
rect 4674 33088 4679 33144
rect 1761 33086 4679 33088
rect 1761 33083 1827 33086
rect 4613 33083 4679 33086
rect 9581 33146 9647 33149
rect 11329 33146 11395 33149
rect 9581 33144 11395 33146
rect 9581 33088 9586 33144
rect 9642 33088 11334 33144
rect 11390 33088 11395 33144
rect 9581 33086 11395 33088
rect 9581 33083 9647 33086
rect 11329 33083 11395 33086
rect 3233 33010 3299 33013
rect 9765 33010 9831 33013
rect 10317 33010 10383 33013
rect 3233 33008 10383 33010
rect 3233 32952 3238 33008
rect 3294 32952 9770 33008
rect 9826 32952 10322 33008
rect 10378 32952 10383 33008
rect 3233 32950 10383 32952
rect 3233 32947 3299 32950
rect 9765 32947 9831 32950
rect 10317 32947 10383 32950
rect 933 32874 999 32877
rect 2773 32874 2839 32877
rect 933 32872 2839 32874
rect 933 32816 938 32872
rect 994 32816 2778 32872
rect 2834 32816 2839 32872
rect 933 32814 2839 32816
rect 933 32811 999 32814
rect 2773 32811 2839 32814
rect 8109 32874 8175 32877
rect 12801 32874 12867 32877
rect 13445 32874 13511 32877
rect 8109 32872 13511 32874
rect 8109 32816 8114 32872
rect 8170 32816 12806 32872
rect 12862 32816 13450 32872
rect 13506 32816 13511 32872
rect 8109 32814 13511 32816
rect 8109 32811 8175 32814
rect 12801 32811 12867 32814
rect 13445 32811 13511 32814
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 4889 32466 4955 32469
rect 9581 32466 9647 32469
rect 4889 32464 9647 32466
rect 4889 32408 4894 32464
rect 4950 32408 9586 32464
rect 9642 32408 9647 32464
rect 4889 32406 9647 32408
rect 4889 32403 4955 32406
rect 9581 32403 9647 32406
rect 1393 32330 1459 32333
rect 5257 32330 5323 32333
rect 1393 32328 5323 32330
rect 1393 32272 1398 32328
rect 1454 32272 5262 32328
rect 5318 32272 5323 32328
rect 1393 32270 5323 32272
rect 1393 32267 1459 32270
rect 5257 32267 5323 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 7189 32058 7255 32061
rect 10961 32058 11027 32061
rect 7189 32056 11027 32058
rect 7189 32000 7194 32056
rect 7250 32000 10966 32056
rect 11022 32000 11027 32056
rect 7189 31998 11027 32000
rect 7189 31995 7255 31998
rect 10961 31995 11027 31998
rect 5809 31786 5875 31789
rect 6821 31786 6887 31789
rect 5809 31784 6887 31786
rect 5809 31728 5814 31784
rect 5870 31728 6826 31784
rect 6882 31728 6887 31784
rect 5809 31726 6887 31728
rect 5809 31723 5875 31726
rect 6821 31723 6887 31726
rect 0 31650 480 31680
rect 1669 31650 1735 31653
rect 0 31648 1735 31650
rect 0 31592 1674 31648
rect 1730 31592 1735 31648
rect 0 31590 1735 31592
rect 0 31560 480 31590
rect 1669 31587 1735 31590
rect 10777 31650 10843 31653
rect 12433 31650 12499 31653
rect 12617 31650 12683 31653
rect 10777 31648 12683 31650
rect 10777 31592 10782 31648
rect 10838 31592 12438 31648
rect 12494 31592 12622 31648
rect 12678 31592 12683 31648
rect 10777 31590 12683 31592
rect 10777 31587 10843 31590
rect 12433 31587 12499 31590
rect 12617 31587 12683 31590
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 1301 31378 1367 31381
rect 7373 31378 7439 31381
rect 1301 31376 7439 31378
rect 1301 31320 1306 31376
rect 1362 31320 7378 31376
rect 7434 31320 7439 31376
rect 1301 31318 7439 31320
rect 1301 31315 1367 31318
rect 7373 31315 7439 31318
rect 10225 31378 10291 31381
rect 12525 31378 12591 31381
rect 10225 31376 12591 31378
rect 10225 31320 10230 31376
rect 10286 31320 12530 31376
rect 12586 31320 12591 31376
rect 10225 31318 12591 31320
rect 10225 31315 10291 31318
rect 12525 31315 12591 31318
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 7925 30834 7991 30837
rect 10777 30834 10843 30837
rect 7925 30832 10843 30834
rect 7925 30776 7930 30832
rect 7986 30776 10782 30832
rect 10838 30776 10843 30832
rect 7925 30774 10843 30776
rect 7925 30771 7991 30774
rect 10777 30771 10843 30774
rect 1669 30698 1735 30701
rect 9765 30698 9831 30701
rect 1669 30696 9831 30698
rect 1669 30640 1674 30696
rect 1730 30640 9770 30696
rect 9826 30640 9831 30696
rect 1669 30638 9831 30640
rect 1669 30635 1735 30638
rect 9765 30635 9831 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 10961 30290 11027 30293
rect 13169 30290 13235 30293
rect 10961 30288 13235 30290
rect 10961 30232 10966 30288
rect 11022 30232 13174 30288
rect 13230 30232 13235 30288
rect 10961 30230 13235 30232
rect 10961 30227 11027 30230
rect 13169 30227 13235 30230
rect 3049 30154 3115 30157
rect 5717 30154 5783 30157
rect 9949 30154 10015 30157
rect 10593 30154 10659 30157
rect 3049 30152 10659 30154
rect 3049 30096 3054 30152
rect 3110 30096 5722 30152
rect 5778 30096 9954 30152
rect 10010 30096 10598 30152
rect 10654 30096 10659 30152
rect 3049 30094 10659 30096
rect 3049 30091 3115 30094
rect 5717 30091 5783 30094
rect 9949 30091 10015 30094
rect 10593 30091 10659 30094
rect 12157 30018 12223 30021
rect 15520 30018 16000 30048
rect 12157 30016 16000 30018
rect 12157 29960 12162 30016
rect 12218 29960 16000 30016
rect 12157 29958 16000 29960
rect 12157 29955 12223 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 0 29338 480 29368
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 1669 29338 1735 29341
rect 0 29336 1735 29338
rect 0 29280 1674 29336
rect 1730 29280 1735 29336
rect 0 29278 1735 29280
rect 0 29248 480 29278
rect 1669 29275 1735 29278
rect 5165 29202 5231 29205
rect 7373 29202 7439 29205
rect 5165 29200 7439 29202
rect 5165 29144 5170 29200
rect 5226 29144 7378 29200
rect 7434 29144 7439 29200
rect 5165 29142 7439 29144
rect 5165 29139 5231 29142
rect 7373 29139 7439 29142
rect 7557 29202 7623 29205
rect 10869 29202 10935 29205
rect 7557 29200 10935 29202
rect 7557 29144 7562 29200
rect 7618 29144 10874 29200
rect 10930 29144 10935 29200
rect 7557 29142 10935 29144
rect 7557 29139 7623 29142
rect 10869 29139 10935 29142
rect 7097 29066 7163 29069
rect 7557 29066 7623 29069
rect 7097 29064 7623 29066
rect 7097 29008 7102 29064
rect 7158 29008 7562 29064
rect 7618 29008 7623 29064
rect 7097 29006 7623 29008
rect 7097 29003 7163 29006
rect 7557 29003 7623 29006
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 7373 28658 7439 28661
rect 12433 28658 12499 28661
rect 7373 28656 12499 28658
rect 7373 28600 7378 28656
rect 7434 28600 12438 28656
rect 12494 28600 12499 28656
rect 7373 28598 12499 28600
rect 7373 28595 7439 28598
rect 12433 28595 12499 28598
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 5257 28114 5323 28117
rect 7649 28114 7715 28117
rect 10409 28114 10475 28117
rect 5257 28112 10475 28114
rect 5257 28056 5262 28112
rect 5318 28056 7654 28112
rect 7710 28056 10414 28112
rect 10470 28056 10475 28112
rect 5257 28054 10475 28056
rect 5257 28051 5323 28054
rect 7649 28051 7715 28054
rect 10409 28051 10475 28054
rect 1669 27842 1735 27845
rect 5533 27842 5599 27845
rect 1669 27840 5599 27842
rect 1669 27784 1674 27840
rect 1730 27784 5538 27840
rect 5594 27784 5599 27840
rect 1669 27782 5599 27784
rect 1669 27779 1735 27782
rect 5533 27779 5599 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 5349 27570 5415 27573
rect 8293 27570 8359 27573
rect 5349 27568 8359 27570
rect 5349 27512 5354 27568
rect 5410 27512 8298 27568
rect 8354 27512 8359 27568
rect 5349 27510 8359 27512
rect 5349 27507 5415 27510
rect 8293 27507 8359 27510
rect 6729 27434 6795 27437
rect 7281 27434 7347 27437
rect 9857 27434 9923 27437
rect 6729 27432 9923 27434
rect 6729 27376 6734 27432
rect 6790 27376 7286 27432
rect 7342 27376 9862 27432
rect 9918 27376 9923 27432
rect 6729 27374 9923 27376
rect 6729 27371 6795 27374
rect 7281 27371 7347 27374
rect 9857 27371 9923 27374
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 0 27026 480 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 480 26966
rect 1577 26963 1643 26966
rect 4521 27026 4587 27029
rect 10041 27026 10107 27029
rect 4521 27024 10107 27026
rect 4521 26968 4526 27024
rect 4582 26968 10046 27024
rect 10102 26968 10107 27024
rect 4521 26966 10107 26968
rect 4521 26963 4587 26966
rect 10041 26963 10107 26966
rect 10133 26892 10199 26893
rect 10133 26890 10180 26892
rect 10088 26888 10180 26890
rect 10088 26832 10138 26888
rect 10088 26830 10180 26832
rect 10133 26828 10180 26830
rect 10244 26828 10250 26892
rect 10133 26827 10199 26828
rect 8017 26754 8083 26757
rect 10133 26754 10199 26757
rect 8017 26752 10199 26754
rect 8017 26696 8022 26752
rect 8078 26696 10138 26752
rect 10194 26696 10199 26752
rect 8017 26694 10199 26696
rect 8017 26691 8083 26694
rect 10133 26691 10199 26694
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 7557 26620 7623 26621
rect 7557 26616 7604 26620
rect 7668 26618 7674 26620
rect 7557 26560 7562 26616
rect 7557 26556 7604 26560
rect 7668 26558 7714 26618
rect 7668 26556 7674 26558
rect 7557 26555 7623 26556
rect 2221 26346 2287 26349
rect 4337 26346 4403 26349
rect 2221 26344 4403 26346
rect 2221 26288 2226 26344
rect 2282 26288 4342 26344
rect 4398 26288 4403 26344
rect 2221 26286 4403 26288
rect 2221 26283 2287 26286
rect 4337 26283 4403 26286
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 7465 25938 7531 25941
rect 9121 25938 9187 25941
rect 7465 25936 9187 25938
rect 7465 25880 7470 25936
rect 7526 25880 9126 25936
rect 9182 25880 9187 25936
rect 7465 25878 9187 25880
rect 7465 25875 7531 25878
rect 9121 25875 9187 25878
rect 2957 25802 3023 25805
rect 6821 25802 6887 25805
rect 2957 25800 6887 25802
rect 2957 25744 2962 25800
rect 3018 25744 6826 25800
rect 6882 25744 6887 25800
rect 2957 25742 6887 25744
rect 2957 25739 3023 25742
rect 6821 25739 6887 25742
rect 2589 25666 2655 25669
rect 4337 25666 4403 25669
rect 2589 25664 4403 25666
rect 2589 25608 2594 25664
rect 2650 25608 4342 25664
rect 4398 25608 4403 25664
rect 2589 25606 4403 25608
rect 2589 25603 2655 25606
rect 4337 25603 4403 25606
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 8017 25530 8083 25533
rect 8293 25530 8359 25533
rect 9397 25530 9463 25533
rect 8017 25528 9463 25530
rect 8017 25472 8022 25528
rect 8078 25472 8298 25528
rect 8354 25472 9402 25528
rect 9458 25472 9463 25528
rect 8017 25470 9463 25472
rect 8017 25467 8083 25470
rect 8293 25467 8359 25470
rect 9397 25467 9463 25470
rect 10961 25394 11027 25397
rect 12525 25394 12591 25397
rect 10961 25392 12591 25394
rect 10961 25336 10966 25392
rect 11022 25336 12530 25392
rect 12586 25336 12591 25392
rect 10961 25334 12591 25336
rect 10961 25331 11027 25334
rect 12525 25331 12591 25334
rect 4613 25258 4679 25261
rect 13261 25258 13327 25261
rect 4613 25256 13327 25258
rect 4613 25200 4618 25256
rect 4674 25200 13266 25256
rect 13322 25200 13327 25256
rect 4613 25198 13327 25200
rect 4613 25195 4679 25198
rect 13261 25195 13327 25198
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 8109 24850 8175 24853
rect 8569 24850 8635 24853
rect 8109 24848 8635 24850
rect 8109 24792 8114 24848
rect 8170 24792 8574 24848
rect 8630 24792 8635 24848
rect 8109 24790 8635 24792
rect 8109 24787 8175 24790
rect 8569 24787 8635 24790
rect 3417 24714 3483 24717
rect 10777 24714 10843 24717
rect 11789 24714 11855 24717
rect 12341 24714 12407 24717
rect 3417 24712 12407 24714
rect 3417 24656 3422 24712
rect 3478 24656 10782 24712
rect 10838 24656 11794 24712
rect 11850 24656 12346 24712
rect 12402 24656 12407 24712
rect 3417 24654 12407 24656
rect 3417 24651 3483 24654
rect 10777 24651 10843 24654
rect 11789 24651 11855 24654
rect 12341 24651 12407 24654
rect 0 24578 480 24608
rect 1669 24578 1735 24581
rect 0 24576 1735 24578
rect 0 24520 1674 24576
rect 1730 24520 1735 24576
rect 0 24518 1735 24520
rect 0 24488 480 24518
rect 1669 24515 1735 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 5901 24306 5967 24309
rect 12709 24306 12775 24309
rect 5901 24304 12775 24306
rect 5901 24248 5906 24304
rect 5962 24248 12714 24304
rect 12770 24248 12775 24304
rect 5901 24246 12775 24248
rect 5901 24243 5967 24246
rect 12709 24243 12775 24246
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 9438 23836 9444 23900
rect 9508 23898 9514 23900
rect 9581 23898 9647 23901
rect 9508 23896 9647 23898
rect 9508 23840 9586 23896
rect 9642 23840 9647 23896
rect 9508 23838 9647 23840
rect 9508 23836 9514 23838
rect 9581 23835 9647 23838
rect 3141 23762 3207 23765
rect 7557 23762 7623 23765
rect 3141 23760 7623 23762
rect 3141 23704 3146 23760
rect 3202 23704 7562 23760
rect 7618 23704 7623 23760
rect 3141 23702 7623 23704
rect 3141 23699 3207 23702
rect 7557 23699 7623 23702
rect 8753 23762 8819 23765
rect 9581 23762 9647 23765
rect 10593 23762 10659 23765
rect 8753 23760 10659 23762
rect 8753 23704 8758 23760
rect 8814 23704 9586 23760
rect 9642 23704 10598 23760
rect 10654 23704 10659 23760
rect 8753 23702 10659 23704
rect 8753 23699 8819 23702
rect 9581 23699 9647 23702
rect 10593 23699 10659 23702
rect 4153 23626 4219 23629
rect 4889 23626 4955 23629
rect 8385 23626 8451 23629
rect 4153 23624 8451 23626
rect 4153 23568 4158 23624
rect 4214 23568 4894 23624
rect 4950 23568 8390 23624
rect 8446 23568 8451 23624
rect 4153 23566 8451 23568
rect 4153 23563 4219 23566
rect 4889 23563 4955 23566
rect 8385 23563 8451 23566
rect 6821 23490 6887 23493
rect 9857 23490 9923 23493
rect 6821 23488 9923 23490
rect 6821 23432 6826 23488
rect 6882 23432 9862 23488
rect 9918 23432 9923 23488
rect 6821 23430 9923 23432
rect 6821 23427 6887 23430
rect 9857 23427 9923 23430
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 2957 23082 3023 23085
rect 7925 23082 7991 23085
rect 8385 23082 8451 23085
rect 2957 23080 8451 23082
rect 2957 23024 2962 23080
rect 3018 23024 7930 23080
rect 7986 23024 8390 23080
rect 8446 23024 8451 23080
rect 2957 23022 8451 23024
rect 2957 23019 3023 23022
rect 7925 23019 7991 23022
rect 8385 23019 8451 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 9489 22812 9555 22813
rect 9438 22748 9444 22812
rect 9508 22810 9555 22812
rect 9508 22808 9600 22810
rect 9550 22752 9600 22808
rect 9508 22750 9600 22752
rect 9508 22748 9555 22750
rect 9489 22747 9555 22748
rect 4613 22538 4679 22541
rect 7833 22538 7899 22541
rect 4613 22536 7899 22538
rect 4613 22480 4618 22536
rect 4674 22480 7838 22536
rect 7894 22480 7899 22536
rect 4613 22478 7899 22480
rect 4613 22475 4679 22478
rect 7833 22475 7899 22478
rect 8109 22538 8175 22541
rect 10133 22538 10199 22541
rect 8109 22536 10199 22538
rect 8109 22480 8114 22536
rect 8170 22480 10138 22536
rect 10194 22480 10199 22536
rect 8109 22478 10199 22480
rect 8109 22475 8175 22478
rect 10133 22475 10199 22478
rect 6277 22336 6597 22337
rect 0 22266 480 22296
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 1669 22266 1735 22269
rect 0 22264 1735 22266
rect 0 22208 1674 22264
rect 1730 22208 1735 22264
rect 0 22206 1735 22208
rect 0 22176 480 22206
rect 1669 22203 1735 22206
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 1393 21042 1459 21045
rect 5717 21042 5783 21045
rect 1393 21040 5783 21042
rect 1393 20984 1398 21040
rect 1454 20984 5722 21040
rect 5778 20984 5783 21040
rect 1393 20982 5783 20984
rect 1393 20979 1459 20982
rect 5717 20979 5783 20982
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 2221 20498 2287 20501
rect 9765 20498 9831 20501
rect 2221 20496 9831 20498
rect 2221 20440 2226 20496
rect 2282 20440 9770 20496
rect 9826 20440 9831 20496
rect 2221 20438 9831 20440
rect 2221 20435 2287 20438
rect 9765 20435 9831 20438
rect 3877 20362 3943 20365
rect 6177 20362 6243 20365
rect 11513 20362 11579 20365
rect 3877 20360 11579 20362
rect 3877 20304 3882 20360
rect 3938 20304 6182 20360
rect 6238 20304 11518 20360
rect 11574 20304 11579 20360
rect 3877 20302 11579 20304
rect 3877 20299 3943 20302
rect 6177 20299 6243 20302
rect 11513 20299 11579 20302
rect 7557 20228 7623 20229
rect 7557 20226 7604 20228
rect 7512 20224 7604 20226
rect 7512 20168 7562 20224
rect 7512 20166 7604 20168
rect 7557 20164 7604 20166
rect 7668 20164 7674 20228
rect 7557 20163 7623 20164
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 9397 20090 9463 20093
rect 9949 20090 10015 20093
rect 11053 20090 11119 20093
rect 9397 20088 11119 20090
rect 9397 20032 9402 20088
rect 9458 20032 9954 20088
rect 10010 20032 11058 20088
rect 11114 20032 11119 20088
rect 9397 20030 11119 20032
rect 9397 20027 9463 20030
rect 9949 20027 10015 20030
rect 11053 20027 11119 20030
rect 0 19954 480 19984
rect 1669 19954 1735 19957
rect 0 19952 1735 19954
rect 0 19896 1674 19952
rect 1730 19896 1735 19952
rect 0 19894 1735 19896
rect 0 19864 480 19894
rect 1669 19891 1735 19894
rect 7925 19954 7991 19957
rect 11421 19954 11487 19957
rect 7925 19952 11487 19954
rect 7925 19896 7930 19952
rect 7986 19896 11426 19952
rect 11482 19896 11487 19952
rect 7925 19894 11487 19896
rect 7925 19891 7991 19894
rect 11421 19891 11487 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 3233 19410 3299 19413
rect 3190 19408 3299 19410
rect 3190 19352 3238 19408
rect 3294 19352 3299 19408
rect 3190 19347 3299 19352
rect 3969 19410 4035 19413
rect 7097 19410 7163 19413
rect 3969 19408 7163 19410
rect 3969 19352 3974 19408
rect 4030 19352 7102 19408
rect 7158 19352 7163 19408
rect 3969 19350 7163 19352
rect 3969 19347 4035 19350
rect 7097 19347 7163 19350
rect 3190 19276 3250 19347
rect 3182 19212 3188 19276
rect 3252 19212 3258 19276
rect 4429 19274 4495 19277
rect 9213 19274 9279 19277
rect 4429 19272 9279 19274
rect 4429 19216 4434 19272
rect 4490 19216 9218 19272
rect 9274 19216 9279 19272
rect 4429 19214 9279 19216
rect 4429 19211 4495 19214
rect 9213 19211 9279 19214
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 4521 17778 4587 17781
rect 10685 17778 10751 17781
rect 4521 17776 10751 17778
rect 4521 17720 4526 17776
rect 4582 17720 10690 17776
rect 10746 17720 10751 17776
rect 4521 17718 10751 17720
rect 4521 17715 4587 17718
rect 10685 17715 10751 17718
rect 0 17642 480 17672
rect 1577 17642 1643 17645
rect 0 17640 1643 17642
rect 0 17584 1582 17640
rect 1638 17584 1643 17640
rect 0 17582 1643 17584
rect 0 17552 480 17582
rect 1577 17579 1643 17582
rect 8661 17642 8727 17645
rect 10593 17642 10659 17645
rect 8661 17640 10659 17642
rect 8661 17584 8666 17640
rect 8722 17584 10598 17640
rect 10654 17584 10659 17640
rect 8661 17582 10659 17584
rect 8661 17579 8727 17582
rect 10593 17579 10659 17582
rect 10409 17506 10475 17509
rect 12709 17506 12775 17509
rect 10409 17504 12775 17506
rect 10409 17448 10414 17504
rect 10470 17448 12714 17504
rect 12770 17448 12775 17504
rect 10409 17446 12775 17448
rect 10409 17443 10475 17446
rect 12709 17443 12775 17446
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 4613 17234 4679 17237
rect 11513 17234 11579 17237
rect 4613 17232 11579 17234
rect 4613 17176 4618 17232
rect 4674 17176 11518 17232
rect 11574 17176 11579 17232
rect 4613 17174 11579 17176
rect 4613 17171 4679 17174
rect 11513 17171 11579 17174
rect 5073 17098 5139 17101
rect 8293 17098 8359 17101
rect 5073 17096 8359 17098
rect 5073 17040 5078 17096
rect 5134 17040 8298 17096
rect 8354 17040 8359 17096
rect 5073 17038 8359 17040
rect 5073 17035 5139 17038
rect 8293 17035 8359 17038
rect 2129 16962 2195 16965
rect 4429 16962 4495 16965
rect 2129 16960 4495 16962
rect 2129 16904 2134 16960
rect 2190 16904 4434 16960
rect 4490 16904 4495 16960
rect 2129 16902 4495 16904
rect 2129 16899 2195 16902
rect 4429 16899 4495 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 5717 16690 5783 16693
rect 8017 16690 8083 16693
rect 9673 16690 9739 16693
rect 5717 16688 9739 16690
rect 5717 16632 5722 16688
rect 5778 16632 8022 16688
rect 8078 16632 9678 16688
rect 9734 16632 9739 16688
rect 5717 16630 9739 16632
rect 5717 16627 5783 16630
rect 8017 16627 8083 16630
rect 9673 16627 9739 16630
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 1393 16146 1459 16149
rect 6913 16146 6979 16149
rect 1393 16144 6979 16146
rect 1393 16088 1398 16144
rect 1454 16088 6918 16144
rect 6974 16088 6979 16144
rect 1393 16086 6979 16088
rect 1393 16083 1459 16086
rect 6913 16083 6979 16086
rect 4061 16010 4127 16013
rect 5073 16010 5139 16013
rect 4061 16008 5139 16010
rect 4061 15952 4066 16008
rect 4122 15952 5078 16008
rect 5134 15952 5139 16008
rect 4061 15950 5139 15952
rect 4061 15947 4127 15950
rect 5073 15947 5139 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3601 15602 3667 15605
rect 11145 15602 11211 15605
rect 3601 15600 11211 15602
rect 3601 15544 3606 15600
rect 3662 15544 11150 15600
rect 11206 15544 11211 15600
rect 3601 15542 11211 15544
rect 3601 15539 3667 15542
rect 11145 15539 11211 15542
rect 3610 15264 3930 15265
rect 0 15194 480 15224
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 480 15134
rect 1669 15131 1735 15134
rect 5349 15194 5415 15197
rect 5717 15194 5783 15197
rect 6637 15194 6703 15197
rect 5349 15192 6703 15194
rect 5349 15136 5354 15192
rect 5410 15136 5722 15192
rect 5778 15136 6642 15192
rect 6698 15136 6703 15192
rect 5349 15134 6703 15136
rect 5349 15131 5415 15134
rect 5717 15131 5783 15134
rect 6637 15131 6703 15134
rect 5809 15060 5875 15061
rect 5758 15058 5764 15060
rect 5718 14998 5764 15058
rect 5828 15056 5875 15060
rect 5870 15000 5875 15056
rect 5758 14996 5764 14998
rect 5828 14996 5875 15000
rect 5809 14995 5875 14996
rect 8569 15058 8635 15061
rect 12341 15058 12407 15061
rect 8569 15056 12407 15058
rect 8569 15000 8574 15056
rect 8630 15000 12346 15056
rect 12402 15000 12407 15056
rect 8569 14998 12407 15000
rect 8569 14995 8635 14998
rect 12341 14995 12407 14998
rect 3417 14922 3483 14925
rect 3601 14922 3667 14925
rect 12065 14922 12131 14925
rect 3417 14920 12131 14922
rect 3417 14864 3422 14920
rect 3478 14864 3606 14920
rect 3662 14864 12070 14920
rect 12126 14864 12131 14920
rect 3417 14862 12131 14864
rect 3417 14859 3483 14862
rect 3601 14859 3667 14862
rect 12065 14859 12131 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 12341 14650 12407 14653
rect 13813 14650 13879 14653
rect 12341 14648 13879 14650
rect 12341 14592 12346 14648
rect 12402 14592 13818 14648
rect 13874 14592 13879 14648
rect 12341 14590 13879 14592
rect 12341 14587 12407 14590
rect 13813 14587 13879 14590
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 2221 13970 2287 13973
rect 7005 13970 7071 13973
rect 2221 13968 7071 13970
rect 2221 13912 2226 13968
rect 2282 13912 7010 13968
rect 7066 13912 7071 13968
rect 2221 13910 7071 13912
rect 2221 13907 2287 13910
rect 7005 13907 7071 13910
rect 3785 13834 3851 13837
rect 9949 13834 10015 13837
rect 3785 13832 10015 13834
rect 3785 13776 3790 13832
rect 3846 13776 9954 13832
rect 10010 13776 10015 13832
rect 3785 13774 10015 13776
rect 3785 13771 3851 13774
rect 9949 13771 10015 13774
rect 5717 13700 5783 13701
rect 5717 13698 5764 13700
rect 5672 13696 5764 13698
rect 5672 13640 5722 13696
rect 5672 13638 5764 13640
rect 5717 13636 5764 13638
rect 5828 13636 5834 13700
rect 8017 13698 8083 13701
rect 10174 13698 10180 13700
rect 8017 13696 10180 13698
rect 8017 13640 8022 13696
rect 8078 13640 10180 13696
rect 8017 13638 10180 13640
rect 5717 13635 5783 13636
rect 8017 13635 8083 13638
rect 10174 13636 10180 13638
rect 10244 13636 10250 13700
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 0 12882 480 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 480 12822
rect 1577 12819 1643 12822
rect 3049 12882 3115 12885
rect 5349 12882 5415 12885
rect 3049 12880 5415 12882
rect 3049 12824 3054 12880
rect 3110 12824 5354 12880
rect 5410 12824 5415 12880
rect 3049 12822 5415 12824
rect 3049 12819 3115 12822
rect 5349 12819 5415 12822
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 2681 12202 2747 12205
rect 8385 12202 8451 12205
rect 2681 12200 8451 12202
rect 2681 12144 2686 12200
rect 2742 12144 8390 12200
rect 8446 12144 8451 12200
rect 2681 12142 8451 12144
rect 2681 12139 2747 12142
rect 8385 12139 8451 12142
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 1393 11794 1459 11797
rect 4521 11794 4587 11797
rect 1393 11792 4587 11794
rect 1393 11736 1398 11792
rect 1454 11736 4526 11792
rect 4582 11736 4587 11792
rect 1393 11734 4587 11736
rect 1393 11731 1459 11734
rect 4521 11731 4587 11734
rect 7373 11522 7439 11525
rect 7557 11522 7623 11525
rect 7373 11520 7623 11522
rect 7373 11464 7378 11520
rect 7434 11464 7562 11520
rect 7618 11464 7623 11520
rect 7373 11462 7623 11464
rect 7373 11459 7439 11462
rect 7557 11459 7623 11462
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 5625 11114 5691 11117
rect 10317 11114 10383 11117
rect 5625 11112 10383 11114
rect 5625 11056 5630 11112
rect 5686 11056 10322 11112
rect 10378 11056 10383 11112
rect 5625 11054 10383 11056
rect 5625 11051 5691 11054
rect 10317 11051 10383 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 4337 10706 4403 10709
rect 10041 10706 10107 10709
rect 4337 10704 10107 10706
rect 4337 10648 4342 10704
rect 4398 10648 10046 10704
rect 10102 10648 10107 10704
rect 4337 10646 10107 10648
rect 4337 10643 4403 10646
rect 10041 10643 10107 10646
rect 10409 10704 10475 10709
rect 10409 10648 10414 10704
rect 10470 10648 10475 10704
rect 10409 10643 10475 10648
rect 0 10570 480 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 480 10510
rect 1577 10507 1643 10510
rect 2497 10570 2563 10573
rect 10412 10570 10472 10643
rect 12341 10570 12407 10573
rect 2497 10568 12407 10570
rect 2497 10512 2502 10568
rect 2558 10512 12346 10568
rect 12402 10512 12407 10568
rect 2497 10510 12407 10512
rect 2497 10507 2563 10510
rect 12341 10507 12407 10510
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 5257 10162 5323 10165
rect 5625 10162 5691 10165
rect 5257 10160 5691 10162
rect 5257 10104 5262 10160
rect 5318 10104 5630 10160
rect 5686 10104 5691 10160
rect 5257 10102 5691 10104
rect 5257 10099 5323 10102
rect 5625 10099 5691 10102
rect 5993 10162 6059 10165
rect 11329 10162 11395 10165
rect 5993 10160 11395 10162
rect 5993 10104 5998 10160
rect 6054 10104 11334 10160
rect 11390 10104 11395 10160
rect 5993 10102 11395 10104
rect 5993 10099 6059 10102
rect 11329 10099 11395 10102
rect 3141 10026 3207 10029
rect 5625 10026 5691 10029
rect 9581 10026 9647 10029
rect 3141 10024 9647 10026
rect 3141 9968 3146 10024
rect 3202 9968 5630 10024
rect 5686 9968 9586 10024
rect 9642 9968 9647 10024
rect 3141 9966 9647 9968
rect 3141 9963 3207 9966
rect 5625 9963 5691 9966
rect 9581 9963 9647 9966
rect 13169 10026 13235 10029
rect 15520 10026 16000 10056
rect 13169 10024 16000 10026
rect 13169 9968 13174 10024
rect 13230 9968 16000 10024
rect 13169 9966 16000 9968
rect 13169 9963 13235 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 2589 9754 2655 9757
rect 2589 9752 2882 9754
rect 2589 9696 2594 9752
rect 2650 9696 2882 9752
rect 2589 9694 2882 9696
rect 2589 9691 2655 9694
rect 2681 9618 2747 9621
rect 2822 9618 2882 9694
rect 3182 9692 3188 9756
rect 3252 9692 3258 9756
rect 3190 9620 3250 9692
rect 2681 9616 2882 9618
rect 2681 9560 2686 9616
rect 2742 9560 2882 9616
rect 2681 9558 2882 9560
rect 2681 9555 2747 9558
rect 3182 9556 3188 9620
rect 3252 9556 3258 9620
rect 7281 9618 7347 9621
rect 11789 9618 11855 9621
rect 7281 9616 11898 9618
rect 7281 9560 7286 9616
rect 7342 9560 11794 9616
rect 11850 9560 11898 9616
rect 7281 9558 11898 9560
rect 7281 9555 7347 9558
rect 11789 9555 11898 9558
rect 2313 9482 2379 9485
rect 3785 9482 3851 9485
rect 2313 9480 3851 9482
rect 2313 9424 2318 9480
rect 2374 9424 3790 9480
rect 3846 9424 3851 9480
rect 2313 9422 3851 9424
rect 2313 9419 2379 9422
rect 3785 9419 3851 9422
rect 7189 9482 7255 9485
rect 10133 9482 10199 9485
rect 7189 9480 10199 9482
rect 7189 9424 7194 9480
rect 7250 9424 10138 9480
rect 10194 9424 10199 9480
rect 7189 9422 10199 9424
rect 11838 9482 11898 9555
rect 12985 9482 13051 9485
rect 11838 9480 13051 9482
rect 11838 9424 12990 9480
rect 13046 9424 13051 9480
rect 11838 9422 13051 9424
rect 7189 9419 7255 9422
rect 10133 9419 10199 9422
rect 12985 9419 13051 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 4337 9212 4403 9213
rect 4286 9148 4292 9212
rect 4356 9210 4403 9212
rect 4356 9208 4448 9210
rect 4398 9152 4448 9208
rect 4356 9150 4448 9152
rect 4356 9148 4403 9150
rect 4337 9147 4403 9148
rect 5073 9074 5139 9077
rect 7005 9074 7071 9077
rect 5073 9072 7071 9074
rect 5073 9016 5078 9072
rect 5134 9016 7010 9072
rect 7066 9016 7071 9072
rect 5073 9014 7071 9016
rect 5073 9011 5139 9014
rect 7005 9011 7071 9014
rect 7465 8938 7531 8941
rect 9857 8938 9923 8941
rect 7465 8936 9923 8938
rect 7465 8880 7470 8936
rect 7526 8880 9862 8936
rect 9918 8880 9923 8936
rect 7465 8878 9923 8880
rect 7465 8875 7531 8878
rect 9857 8875 9923 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 4705 8666 4771 8669
rect 5349 8666 5415 8669
rect 8201 8666 8267 8669
rect 4705 8664 8267 8666
rect 4705 8608 4710 8664
rect 4766 8608 5354 8664
rect 5410 8608 8206 8664
rect 8262 8608 8267 8664
rect 4705 8606 8267 8608
rect 4705 8603 4771 8606
rect 5349 8603 5415 8606
rect 8201 8603 8267 8606
rect 2129 8530 2195 8533
rect 7833 8530 7899 8533
rect 2129 8528 7899 8530
rect 2129 8472 2134 8528
rect 2190 8472 7838 8528
rect 7894 8472 7899 8528
rect 2129 8470 7899 8472
rect 2129 8467 2195 8470
rect 7833 8467 7899 8470
rect 7373 8394 7439 8397
rect 12709 8394 12775 8397
rect 13077 8394 13143 8397
rect 7373 8392 13143 8394
rect 7373 8336 7378 8392
rect 7434 8336 12714 8392
rect 12770 8336 13082 8392
rect 13138 8336 13143 8392
rect 7373 8334 13143 8336
rect 7373 8331 7439 8334
rect 12709 8331 12775 8334
rect 13077 8331 13143 8334
rect 6277 8192 6597 8193
rect 0 8122 480 8152
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 480 8062
rect 1577 8059 1643 8062
rect 3049 7986 3115 7989
rect 7189 7986 7255 7989
rect 8569 7986 8635 7989
rect 3049 7984 8635 7986
rect 3049 7928 3054 7984
rect 3110 7928 7194 7984
rect 7250 7928 8574 7984
rect 8630 7928 8635 7984
rect 3049 7926 8635 7928
rect 3049 7923 3115 7926
rect 7189 7923 7255 7926
rect 8569 7923 8635 7926
rect 4061 7850 4127 7853
rect 10041 7850 10107 7853
rect 4061 7848 10107 7850
rect 4061 7792 4066 7848
rect 4122 7792 10046 7848
rect 10102 7792 10107 7848
rect 4061 7790 10107 7792
rect 4061 7787 4127 7790
rect 10041 7787 10107 7790
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 2313 7442 2379 7445
rect 9857 7442 9923 7445
rect 2313 7440 9923 7442
rect 2313 7384 2318 7440
rect 2374 7384 9862 7440
rect 9918 7384 9923 7440
rect 2313 7382 9923 7384
rect 2313 7379 2379 7382
rect 9857 7379 9923 7382
rect 4797 7306 4863 7309
rect 7925 7306 7991 7309
rect 4797 7304 7991 7306
rect 4797 7248 4802 7304
rect 4858 7248 7930 7304
rect 7986 7248 7991 7304
rect 4797 7246 7991 7248
rect 4797 7243 4863 7246
rect 7925 7243 7991 7246
rect 7189 7170 7255 7173
rect 11421 7170 11487 7173
rect 7189 7168 11487 7170
rect 7189 7112 7194 7168
rect 7250 7112 11426 7168
rect 11482 7112 11487 7168
rect 7189 7110 11487 7112
rect 7189 7107 7255 7110
rect 11421 7107 11487 7110
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 7925 7034 7991 7037
rect 10225 7034 10291 7037
rect 7925 7032 10291 7034
rect 7925 6976 7930 7032
rect 7986 6976 10230 7032
rect 10286 6976 10291 7032
rect 7925 6974 10291 6976
rect 7925 6971 7991 6974
rect 10225 6971 10291 6974
rect 4613 6898 4679 6901
rect 7465 6898 7531 6901
rect 4613 6896 7531 6898
rect 4613 6840 4618 6896
rect 4674 6840 7470 6896
rect 7526 6840 7531 6896
rect 4613 6838 7531 6840
rect 4613 6835 4679 6838
rect 7465 6835 7531 6838
rect 7741 6898 7807 6901
rect 12801 6898 12867 6901
rect 7741 6896 12867 6898
rect 7741 6840 7746 6896
rect 7802 6840 12806 6896
rect 12862 6840 12867 6896
rect 7741 6838 12867 6840
rect 7741 6835 7807 6838
rect 12801 6835 12867 6838
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 8293 6218 8359 6221
rect 9673 6218 9739 6221
rect 8293 6216 9739 6218
rect 8293 6160 8298 6216
rect 8354 6160 9678 6216
rect 9734 6160 9739 6216
rect 8293 6158 9739 6160
rect 8293 6155 8359 6158
rect 9673 6155 9739 6158
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 0 5810 480 5840
rect 2773 5810 2839 5813
rect 0 5808 2839 5810
rect 0 5752 2778 5808
rect 2834 5752 2839 5808
rect 0 5750 2839 5752
rect 0 5720 480 5750
rect 2773 5747 2839 5750
rect 10041 5810 10107 5813
rect 12617 5810 12683 5813
rect 10041 5808 12683 5810
rect 10041 5752 10046 5808
rect 10102 5752 12622 5808
rect 12678 5752 12683 5808
rect 10041 5750 12683 5752
rect 10041 5747 10107 5750
rect 12617 5747 12683 5750
rect 2957 5674 3023 5677
rect 6913 5674 6979 5677
rect 2957 5672 6979 5674
rect 2957 5616 2962 5672
rect 3018 5616 6918 5672
rect 6974 5616 6979 5672
rect 2957 5614 6979 5616
rect 2957 5611 3023 5614
rect 6913 5611 6979 5614
rect 5349 5538 5415 5541
rect 6729 5538 6795 5541
rect 5349 5536 6795 5538
rect 5349 5480 5354 5536
rect 5410 5480 6734 5536
rect 6790 5480 6795 5536
rect 5349 5478 6795 5480
rect 5349 5475 5415 5478
rect 6729 5475 6795 5478
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 4521 5402 4587 5405
rect 7005 5402 7071 5405
rect 4521 5400 7071 5402
rect 4521 5344 4526 5400
rect 4582 5344 7010 5400
rect 7066 5344 7071 5400
rect 4521 5342 7071 5344
rect 4521 5339 4587 5342
rect 7005 5339 7071 5342
rect 4429 5266 4495 5269
rect 8017 5266 8083 5269
rect 4429 5264 8083 5266
rect 4429 5208 4434 5264
rect 4490 5208 8022 5264
rect 8078 5208 8083 5264
rect 4429 5206 8083 5208
rect 4429 5203 4495 5206
rect 8017 5203 8083 5206
rect 11145 5130 11211 5133
rect 12433 5130 12499 5133
rect 11145 5128 12499 5130
rect 11145 5072 11150 5128
rect 11206 5072 12438 5128
rect 12494 5072 12499 5128
rect 11145 5070 12499 5072
rect 11145 5067 11211 5070
rect 12433 5067 12499 5070
rect 2405 4994 2471 4997
rect 4153 4994 4219 4997
rect 2405 4992 4219 4994
rect 2405 4936 2410 4992
rect 2466 4936 4158 4992
rect 4214 4936 4219 4992
rect 2405 4934 4219 4936
rect 2405 4931 2471 4934
rect 4153 4931 4219 4934
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 8661 4858 8727 4861
rect 10961 4858 11027 4861
rect 8661 4856 11027 4858
rect 8661 4800 8666 4856
rect 8722 4800 10966 4856
rect 11022 4800 11027 4856
rect 8661 4798 11027 4800
rect 8661 4795 8727 4798
rect 10961 4795 11027 4798
rect 2681 4722 2747 4725
rect 4429 4722 4495 4725
rect 2681 4720 4495 4722
rect 2681 4664 2686 4720
rect 2742 4664 4434 4720
rect 4490 4664 4495 4720
rect 2681 4662 4495 4664
rect 2681 4659 2747 4662
rect 4429 4659 4495 4662
rect 2497 4586 2563 4589
rect 4521 4586 4587 4589
rect 2497 4584 4587 4586
rect 2497 4528 2502 4584
rect 2558 4528 4526 4584
rect 4582 4528 4587 4584
rect 2497 4526 4587 4528
rect 2497 4523 2563 4526
rect 4521 4523 4587 4526
rect 7097 4586 7163 4589
rect 15745 4586 15811 4589
rect 7097 4584 15811 4586
rect 7097 4528 7102 4584
rect 7158 4528 15750 4584
rect 15806 4528 15811 4584
rect 7097 4526 15811 4528
rect 7097 4523 7163 4526
rect 15745 4523 15811 4526
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 9949 4314 10015 4317
rect 13077 4314 13143 4317
rect 9949 4312 13143 4314
rect 9949 4256 9954 4312
rect 10010 4256 13082 4312
rect 13138 4256 13143 4312
rect 9949 4254 13143 4256
rect 9949 4251 10015 4254
rect 13077 4251 13143 4254
rect 8661 4178 8727 4181
rect 10501 4178 10567 4181
rect 8661 4176 10567 4178
rect 8661 4120 8666 4176
rect 8722 4120 10506 4176
rect 10562 4120 10567 4176
rect 8661 4118 10567 4120
rect 8661 4115 8727 4118
rect 10501 4115 10567 4118
rect 2865 4042 2931 4045
rect 5257 4042 5323 4045
rect 2865 4040 5323 4042
rect 2865 3984 2870 4040
rect 2926 3984 5262 4040
rect 5318 3984 5323 4040
rect 2865 3982 5323 3984
rect 2865 3979 2931 3982
rect 5257 3979 5323 3982
rect 8201 4042 8267 4045
rect 11881 4042 11947 4045
rect 8201 4040 11947 4042
rect 8201 3984 8206 4040
rect 8262 3984 11886 4040
rect 11942 3984 11947 4040
rect 8201 3982 11947 3984
rect 8201 3979 8267 3982
rect 11881 3979 11947 3982
rect 13537 4042 13603 4045
rect 14917 4042 14983 4045
rect 13537 4040 14983 4042
rect 13537 3984 13542 4040
rect 13598 3984 14922 4040
rect 14978 3984 14983 4040
rect 13537 3982 14983 3984
rect 13537 3979 13603 3982
rect 14917 3979 14983 3982
rect 4889 3906 4955 3909
rect 5993 3906 6059 3909
rect 4889 3904 6059 3906
rect 4889 3848 4894 3904
rect 4950 3848 5998 3904
rect 6054 3848 6059 3904
rect 4889 3846 6059 3848
rect 4889 3843 4955 3846
rect 5993 3843 6059 3846
rect 13261 3906 13327 3909
rect 14641 3906 14707 3909
rect 13261 3904 14707 3906
rect 13261 3848 13266 3904
rect 13322 3848 14646 3904
rect 14702 3848 14707 3904
rect 13261 3846 14707 3848
rect 13261 3843 13327 3846
rect 14641 3843 14707 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 6821 3770 6887 3773
rect 10041 3770 10107 3773
rect 6821 3768 10107 3770
rect 6821 3712 6826 3768
rect 6882 3712 10046 3768
rect 10102 3712 10107 3768
rect 6821 3710 10107 3712
rect 6821 3707 6887 3710
rect 10041 3707 10107 3710
rect 933 3634 999 3637
rect 4286 3634 4292 3636
rect 933 3632 4292 3634
rect 933 3576 938 3632
rect 994 3576 4292 3632
rect 933 3574 4292 3576
rect 933 3571 999 3574
rect 4286 3572 4292 3574
rect 4356 3634 4362 3636
rect 9673 3634 9739 3637
rect 10685 3634 10751 3637
rect 4356 3632 10751 3634
rect 4356 3576 9678 3632
rect 9734 3576 10690 3632
rect 10746 3576 10751 3632
rect 4356 3574 10751 3576
rect 4356 3572 4362 3574
rect 9673 3571 9739 3574
rect 10685 3571 10751 3574
rect 11513 3634 11579 3637
rect 15377 3634 15443 3637
rect 11513 3632 15443 3634
rect 11513 3576 11518 3632
rect 11574 3576 15382 3632
rect 15438 3576 15443 3632
rect 11513 3574 15443 3576
rect 11513 3571 11579 3574
rect 15377 3571 15443 3574
rect 0 3498 480 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 2957 3498 3023 3501
rect 3182 3498 3188 3500
rect 2957 3496 3188 3498
rect 2957 3440 2962 3496
rect 3018 3440 3188 3496
rect 2957 3438 3188 3440
rect 2957 3435 3023 3438
rect 3182 3436 3188 3438
rect 3252 3436 3258 3500
rect 12801 3498 12867 3501
rect 3374 3496 12867 3498
rect 3374 3440 12806 3496
rect 12862 3440 12867 3496
rect 3374 3438 12867 3440
rect 1669 3362 1735 3365
rect 3374 3362 3434 3438
rect 12801 3435 12867 3438
rect 1669 3360 3434 3362
rect 1669 3304 1674 3360
rect 1730 3304 3434 3360
rect 1669 3302 3434 3304
rect 1669 3299 1735 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 4797 3226 4863 3229
rect 10133 3226 10199 3229
rect 12617 3226 12683 3229
rect 4797 3224 8770 3226
rect 4797 3168 4802 3224
rect 4858 3168 8770 3224
rect 4797 3166 8770 3168
rect 4797 3163 4863 3166
rect 4245 3090 4311 3093
rect 8569 3090 8635 3093
rect 4245 3088 8635 3090
rect 4245 3032 4250 3088
rect 4306 3032 8574 3088
rect 8630 3032 8635 3088
rect 4245 3030 8635 3032
rect 8710 3090 8770 3166
rect 10133 3224 12683 3226
rect 10133 3168 10138 3224
rect 10194 3168 12622 3224
rect 12678 3168 12683 3224
rect 10133 3166 12683 3168
rect 10133 3163 10199 3166
rect 12617 3163 12683 3166
rect 12433 3090 12499 3093
rect 8710 3088 12499 3090
rect 8710 3032 12438 3088
rect 12494 3032 12499 3088
rect 8710 3030 12499 3032
rect 4245 3027 4311 3030
rect 8569 3027 8635 3030
rect 12433 3027 12499 3030
rect 10961 2954 11027 2957
rect 12617 2954 12683 2957
rect 10961 2952 12683 2954
rect 10961 2896 10966 2952
rect 11022 2896 12622 2952
rect 12678 2896 12683 2952
rect 10961 2894 12683 2896
rect 10961 2891 11027 2894
rect 12617 2891 12683 2894
rect 3417 2818 3483 2821
rect 12065 2818 12131 2821
rect 13353 2818 13419 2821
rect 3417 2816 4170 2818
rect 3417 2760 3422 2816
rect 3478 2760 4170 2816
rect 3417 2758 4170 2760
rect 3417 2755 3483 2758
rect 4110 2682 4170 2758
rect 12065 2816 13419 2818
rect 12065 2760 12070 2816
rect 12126 2760 13358 2816
rect 13414 2760 13419 2816
rect 12065 2758 13419 2760
rect 12065 2755 12131 2758
rect 13353 2755 13419 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 5533 2682 5599 2685
rect 4110 2680 5599 2682
rect 4110 2624 5538 2680
rect 5594 2624 5599 2680
rect 4110 2622 5599 2624
rect 5533 2619 5599 2622
rect 7465 2682 7531 2685
rect 9949 2682 10015 2685
rect 7465 2680 10015 2682
rect 7465 2624 7470 2680
rect 7526 2624 9954 2680
rect 10010 2624 10015 2680
rect 7465 2622 10015 2624
rect 7465 2619 7531 2622
rect 9949 2619 10015 2622
rect 6085 2546 6151 2549
rect 12617 2546 12683 2549
rect 6085 2544 12683 2546
rect 6085 2488 6090 2544
rect 6146 2488 12622 2544
rect 12678 2488 12683 2544
rect 6085 2486 12683 2488
rect 6085 2483 6151 2486
rect 12617 2483 12683 2486
rect 10869 2410 10935 2413
rect 12709 2410 12775 2413
rect 10869 2408 12775 2410
rect 10869 2352 10874 2408
rect 10930 2352 12714 2408
rect 12770 2352 12775 2408
rect 10869 2350 12775 2352
rect 10869 2347 10935 2350
rect 12709 2347 12775 2350
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 6913 1458 6979 1461
rect 10777 1458 10843 1461
rect 6913 1456 10843 1458
rect 6913 1400 6918 1456
rect 6974 1400 10782 1456
rect 10838 1400 10843 1456
rect 6913 1398 10843 1400
rect 6913 1395 6979 1398
rect 10777 1395 10843 1398
rect 11329 1458 11395 1461
rect 12801 1458 12867 1461
rect 11329 1456 12867 1458
rect 11329 1400 11334 1456
rect 11390 1400 12806 1456
rect 12862 1400 12867 1456
rect 11329 1398 12867 1400
rect 11329 1395 11395 1398
rect 12801 1395 12867 1398
rect 0 1186 480 1216
rect 1485 1186 1551 1189
rect 0 1184 1551 1186
rect 0 1128 1490 1184
rect 1546 1128 1551 1184
rect 0 1126 1551 1128
rect 0 1096 480 1126
rect 1485 1123 1551 1126
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 10180 26888 10244 26892
rect 10180 26832 10194 26888
rect 10194 26832 10244 26888
rect 10180 26828 10244 26832
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 7604 26616 7668 26620
rect 7604 26560 7618 26616
rect 7618 26560 7668 26616
rect 7604 26556 7668 26560
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 9444 23836 9508 23900
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 9444 22808 9508 22812
rect 9444 22752 9494 22808
rect 9494 22752 9508 22808
rect 9444 22748 9508 22752
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 7604 20224 7668 20228
rect 7604 20168 7618 20224
rect 7618 20168 7668 20224
rect 7604 20164 7668 20168
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 3188 19212 3252 19276
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 5764 15056 5828 15060
rect 5764 15000 5814 15056
rect 5814 15000 5828 15056
rect 5764 14996 5828 15000
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 5764 13696 5828 13700
rect 5764 13640 5778 13696
rect 5778 13640 5828 13696
rect 5764 13636 5828 13640
rect 10180 13636 10244 13700
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 3188 9692 3252 9756
rect 3188 9556 3252 9620
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 4292 9208 4356 9212
rect 4292 9152 4342 9208
rect 4342 9152 4356 9208
rect 4292 9148 4356 9152
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 4292 3572 4356 3636
rect 3188 3436 3252 3500
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3187 19276 3253 19277
rect 3187 19212 3188 19276
rect 3252 19212 3253 19276
rect 3187 19211 3253 19212
rect 3190 9757 3250 19211
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 7603 26620 7669 26621
rect 7603 26556 7604 26620
rect 7668 26556 7669 26620
rect 7603 26555 7669 26556
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 7606 20229 7666 26555
rect 8944 26144 9264 27168
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 10179 26892 10245 26893
rect 10179 26828 10180 26892
rect 10244 26828 10245 26892
rect 10179 26827 10245 26828
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 9443 23900 9509 23901
rect 9443 23836 9444 23900
rect 9508 23836 9509 23900
rect 9443 23835 9509 23836
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 9446 22813 9506 23835
rect 9443 22812 9509 22813
rect 9443 22748 9444 22812
rect 9508 22748 9509 22812
rect 9443 22747 9509 22748
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 7603 20228 7669 20229
rect 7603 20164 7604 20228
rect 7668 20164 7669 20228
rect 7603 20163 7669 20164
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 5763 15060 5829 15061
rect 5763 14996 5764 15060
rect 5828 14996 5829 15060
rect 5763 14995 5829 14996
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 5766 13701 5826 14995
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 5763 13700 5829 13701
rect 5763 13636 5764 13700
rect 5828 13636 5829 13700
rect 5763 13635 5829 13636
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3187 9756 3253 9757
rect 3187 9692 3188 9756
rect 3252 9692 3253 9756
rect 3187 9691 3253 9692
rect 3187 9620 3253 9621
rect 3187 9556 3188 9620
rect 3252 9556 3253 9620
rect 3187 9555 3253 9556
rect 3190 3501 3250 9555
rect 3610 8736 3931 9760
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 4291 9212 4357 9213
rect 4291 9148 4292 9212
rect 4356 9148 4357 9212
rect 4291 9147 4357 9148
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3187 3500 3253 3501
rect 3187 3436 3188 3500
rect 3252 3436 3253 3500
rect 3187 3435 3253 3436
rect 3610 3296 3931 4320
rect 4294 3637 4354 9147
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 4291 3636 4357 3637
rect 4291 3572 4292 3636
rect 4356 3572 4357 3636
rect 4291 3571 4357 3572
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 10182 13701 10242 26827
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 10179 13700 10245 13701
rect 10179 13636 10180 13700
rect 10244 13636 10245 13700
rect 10179 13635 10245 13636
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_fill_2  FILLER_1_9 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_1.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l2_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_52
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _53_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_92
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_115 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_133 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_139 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_145
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_40
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_98
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_9
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 130 592
use scs8hd_conb_1  _22_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_20
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_24
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_134
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_21
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_91
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_7_28
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_35
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_39
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_67
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_81
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 1786 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_131
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use scs8hd_buf_4  mux_right_ipin_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_9
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_13
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_20
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_24
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_89
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 1786 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_4  mux_left_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_9
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_21
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_137
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_131
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_14
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_38
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_110
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_114
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_43
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_138
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_21
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_76
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_103
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_13
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_26
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_101
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_4  mux_right_ipin_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_9
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_32
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l4_in_0_
timestamp 1586364061
transform 1 0 6900 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_72
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_76
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_12
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_18
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_25
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l2_in_2_
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_8
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_67
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_85
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_89
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_103
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_9
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_48
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_24_60
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_4  mux_right_ipin_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_9
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_13
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_17
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_55
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_6.mux_l3_in_1_
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_20
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_84
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_87
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_8
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_49
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_70
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_49
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_104
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_120
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_35
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_42
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_54
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_7.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_114
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_126
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2300 0 1 19040
box -38 -48 1786 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_42
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_85
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_29
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_32_101
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_135
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 590 592
use scs8hd_buf_4  mux_right_ipin_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_16
timestamp 1586364061
transform 1 0 2576 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_13
timestamp 1586364061
transform 1 0 2300 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_9
timestamp 1586364061
transform 1 0 1932 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_33_13
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_9
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_28
timestamp 1586364061
transform 1 0 3680 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_24
timestamp 1586364061
transform 1 0 3312 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3496 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_55
timestamp 1586364061
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_51
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_65
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_78
timestamp 1586364061
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_90
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_124
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_136
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_144
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_9
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_16
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3496 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_45
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_49
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8096 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_68
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_72
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_85
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_89
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_102
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_108
timestamp 1586364061
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_11
timestamp 1586364061
transform 1 0 2116 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_41
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_8  FILLER_36_58
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_79
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_97
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_36_101
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_24
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_36
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_44
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_48
timestamp 1586364061
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_52
timestamp 1586364061
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_56
timestamp 1586364061
transform 1 0 6256 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_60
timestamp 1586364061
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_67
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_84
timestamp 1586364061
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_105
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_10
timestamp 1586364061
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_6  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_38
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5336 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5060 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_41
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_45
timestamp 1586364061
transform 1 0 5244 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_55
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_63
timestamp 1586364061
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_97
timestamp 1586364061
transform 1 0 10028 0 -1 23392
box -38 -48 406 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_101
timestamp 1586364061
transform 1 0 10396 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_111
timestamp 1586364061
transform 1 0 11316 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_115
timestamp 1586364061
transform 1 0 11684 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_122
timestamp 1586364061
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_130
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_142
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1932 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_26
timestamp 1586364061
transform 1 0 3496 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_22
timestamp 1586364061
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_29
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_25
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3312 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 222 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4508 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_35
timestamp 1586364061
transform 1 0 4324 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_39
timestamp 1586364061
transform 1 0 4692 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6072 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_48
timestamp 1586364061
transform 1 0 5520 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_52
timestamp 1586364061
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_56
timestamp 1586364061
transform 1 0 6256 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_43
timestamp 1586364061
transform 1 0 5060 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_55
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_63
timestamp 1586364061
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_69
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_65
timestamp 1586364061
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_60
timestamp 1586364061
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 24480
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11132 0 -1 24480
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_107
timestamp 1586364061
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_144
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l3_in_1_
timestamp 1586364061
transform 1 0 2668 0 1 24480
box -38 -48 866 592
use scs8hd_buf_4  mux_right_ipin_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 590 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_9
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_13
timestamp 1586364061
transform 1 0 2300 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_16
timestamp 1586364061
transform 1 0 2576 0 1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4232 0 1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_26
timestamp 1586364061
transform 1 0 3496 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_30
timestamp 1586364061
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6992 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_66
timestamp 1586364061
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_70
timestamp 1586364061
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_83
timestamp 1586364061
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_87
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_100
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_104
timestamp 1586364061
transform 1 0 10672 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_107
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_111
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_115
timestamp 1586364061
transform 1 0 11684 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_144
timestamp 1586364061
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 2208 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_7
timestamp 1586364061
transform 1 0 1748 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_10
timestamp 1586364061
transform 1 0 2024 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_10.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5796 0 -1 25568
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_41
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_45
timestamp 1586364061
transform 1 0 5244 0 -1 25568
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_70
timestamp 1586364061
transform 1 0 7544 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_76
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_88
timestamp 1586364061
transform 1 0 9200 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_97
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_42_101
timestamp 1586364061
transform 1 0 10396 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 12696 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_124
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_128
timestamp 1586364061
transform 1 0 12880 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_140
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2668 0 1 25568
box -38 -48 1786 592
use scs8hd_buf_4  mux_right_ipin_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 590 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2116 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_9
timestamp 1586364061
transform 1 0 1932 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_13
timestamp 1586364061
transform 1 0 2300 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4600 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_36
timestamp 1586364061
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5336 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_40
timestamp 1586364061
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_44
timestamp 1586364061
transform 1 0 5152 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_48
timestamp 1586364061
transform 1 0 5520 0 1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_43_54
timestamp 1586364061
transform 1 0 6072 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_57
timestamp 1586364061
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7268 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8280 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_66
timestamp 1586364061
transform 1 0 7176 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_76
timestamp 1586364061
transform 1 0 8096 0 1 25568
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9844 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9660 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8924 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_80
timestamp 1586364061
transform 1 0 8464 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_84
timestamp 1586364061
transform 1 0 8832 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_87
timestamp 1586364061
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_91
timestamp 1586364061
transform 1 0 9476 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_104
timestamp 1586364061
transform 1 0 10672 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_120
timestamp 1586364061
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2668 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_19
timestamp 1586364061
transform 1 0 2852 0 -1 26656
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4232 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5244 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6440 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_43
timestamp 1586364061
transform 1 0 5060 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_47
timestamp 1586364061
transform 1 0 5428 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_44_55
timestamp 1586364061
transform 1 0 6164 0 -1 26656
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6992 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6808 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8004 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_60
timestamp 1586364061
transform 1 0 6624 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_73
timestamp 1586364061
transform 1 0 7820 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_77
timestamp 1586364061
transform 1 0 8188 0 -1 26656
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_44_89
timestamp 1586364061
transform 1 0 9292 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_102
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_114
timestamp 1586364061
transform 1 0 11592 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_126
timestamp 1586364061
transform 1 0 12696 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_44_138
timestamp 1586364061
transform 1 0 13800 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4508 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3956 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_29
timestamp 1586364061
transform 1 0 3772 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_33
timestamp 1586364061
transform 1 0 4140 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5520 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_46
timestamp 1586364061
transform 1 0 5336 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_50
timestamp 1586364061
transform 1 0 5704 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_54
timestamp 1586364061
transform 1 0 6072 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_58
timestamp 1586364061
transform 1 0 6440 0 1 26656
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_71
timestamp 1586364061
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_75
timestamp 1586364061
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_79
timestamp 1586364061
transform 1 0 8372 0 1 26656
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9660 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10028 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_91
timestamp 1586364061
transform 1 0 9476 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_95
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_99
timestamp 1586364061
transform 1 0 10212 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_103
timestamp 1586364061
transform 1 0 10580 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_45_115
timestamp 1586364061
transform 1 0 11684 0 1 26656
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_45_121
timestamp 1586364061
transform 1 0 12236 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_47_7
timestamp 1586364061
transform 1 0 1748 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_11
timestamp 1586364061
transform 1 0 2116 0 1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_46_11
timestamp 1586364061
transform 1 0 2116 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2392 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2208 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_16
timestamp 1586364061
transform 1 0 2576 0 -1 27744
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2392 0 1 27744
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4324 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_28
timestamp 1586364061
transform 1 0 3680 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_33
timestamp 1586364061
transform 1 0 4140 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_37
timestamp 1586364061
transform 1 0 4508 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 -1 27744
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4968 0 -1 27744
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4876 0 1 27744
box -38 -48 866 592
use scs8hd_decap_3  FILLER_47_58
timestamp 1586364061
transform 1 0 6440 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_54
timestamp 1586364061
transform 1 0 6072 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_50
timestamp 1586364061
transform 1 0 5704 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_46_51
timestamp 1586364061
transform 1 0 5796 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6256 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5888 0 1 27744
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l4_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_68
timestamp 1586364061
transform 1 0 7360 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 7084 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_72
timestamp 1586364061
transform 1 0 7728 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_72
timestamp 1586364061
transform 1 0 7728 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8096 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7544 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7544 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_78
timestamp 1586364061
transform 1 0 8280 0 -1 27744
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_90
timestamp 1586364061
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_95
timestamp 1586364061
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_99
timestamp 1586364061
transform 1 0 10212 0 1 27744
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10580 0 1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10396 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10948 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_106
timestamp 1586364061
transform 1 0 10856 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_109
timestamp 1586364061
transform 1 0 11132 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_112
timestamp 1586364061
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_47_116
timestamp 1586364061
transform 1 0 11776 0 1 27744
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_121
timestamp 1586364061
transform 1 0 12236 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_133
timestamp 1586364061
transform 1 0 13340 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 590 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_9
timestamp 1586364061
transform 1 0 1932 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_21
timestamp 1586364061
transform 1 0 3036 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_29
timestamp 1586364061
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_36
timestamp 1586364061
transform 1 0 4416 0 -1 28832
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4784 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5796 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6440 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_49
timestamp 1586364061
transform 1 0 5612 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_53
timestamp 1586364061
transform 1 0 5980 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_57
timestamp 1586364061
transform 1 0 6348 0 -1 28832
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7084 0 -1 28832
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6808 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_60
timestamp 1586364061
transform 1 0 6624 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_64
timestamp 1586364061
transform 1 0 6992 0 -1 28832
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10212 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_84
timestamp 1586364061
transform 1 0 8832 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_6  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10948 0 -1 28832
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_101
timestamp 1586364061
transform 1 0 10396 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_126
timestamp 1586364061
transform 1 0 12696 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_138
timestamp 1586364061
transform 1 0 13800 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 28832
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_31
timestamp 1586364061
transform 1 0 3956 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_53
timestamp 1586364061
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_71
timestamp 1586364061
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_75
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8556 0 1 28832
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10488 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10856 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_100
timestamp 1586364061
transform 1 0 10304 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_104
timestamp 1586364061
transform 1 0 10672 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_108
timestamp 1586364061
transform 1 0 11040 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_118
timestamp 1586364061
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_127
timestamp 1586364061
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_49_139
timestamp 1586364061
transform 1 0 13892 0 1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_49_145
timestamp 1586364061
transform 1 0 14444 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_23
timestamp 1586364061
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7636 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7084 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_63
timestamp 1586364061
transform 1 0 6900 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_67
timestamp 1586364061
transform 1 0 7268 0 -1 29920
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10212 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8648 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_84
timestamp 1586364061
transform 1 0 8832 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_97
timestamp 1586364061
transform 1 0 10028 0 -1 29920
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11776 0 -1 29920
box -38 -48 866 592
use scs8hd_decap_8  FILLER_50_108
timestamp 1586364061
transform 1 0 11040 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_12  FILLER_50_125
timestamp 1586364061
transform 1 0 12604 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_137
timestamp 1586364061
transform 1 0 13708 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_7
timestamp 1586364061
transform 1 0 1748 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_51_19
timestamp 1586364061
transform 1 0 2852 0 1 29920
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3404 0 1 29920
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3220 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_44
timestamp 1586364061
transform 1 0 5152 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  FILLER_51_52
timestamp 1586364061
transform 1 0 5888 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_57
timestamp 1586364061
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_12.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_71
timestamp 1586364061
transform 1 0 7636 0 1 29920
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9752 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9568 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_83
timestamp 1586364061
transform 1 0 8740 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_87
timestamp 1586364061
transform 1 0 9108 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_90
timestamp 1586364061
transform 1 0 9384 0 1 29920
box -38 -48 222 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 11316 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11040 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_103
timestamp 1586364061
transform 1 0 10580 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_107
timestamp 1586364061
transform 1 0 10948 0 1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_114
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_118
timestamp 1586364061
transform 1 0 11960 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_9
timestamp 1586364061
transform 1 0 1932 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_8  FILLER_52_21
timestamp 1586364061
transform 1 0 3036 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_52_29
timestamp 1586364061
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6808 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_64
timestamp 1586364061
transform 1 0 6992 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_76
timestamp 1586364061
transform 1 0 8096 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_66
timestamp 1586364061
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_70
timestamp 1586364061
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_84
timestamp 1586364061
transform 1 0 8832 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8648 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_97
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_97
timestamp 1586364061
transform 1 0 10028 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_90
timestamp 1586364061
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_101
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_107
timestamp 1586364061
transform 1 0 10948 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_101
timestamp 1586364061
transform 1 0 10396 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l2_in_2_
timestamp 1586364061
transform 1 0 10764 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_118
timestamp 1586364061
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_114
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11040 0 -1 31008
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 13432 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_127
timestamp 1586364061
transform 1 0 12788 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_132
timestamp 1586364061
transform 1 0 13248 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_53_136
timestamp 1586364061
transform 1 0 13616 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_decap_6  FILLER_52_139
timestamp 1586364061
transform 1 0 13892 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_144
timestamp 1586364061
transform 1 0 14352 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2300 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 1932 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_7
timestamp 1586364061
transform 1 0 1748 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_11
timestamp 1586364061
transform 1 0 2116 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4232 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3036 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_23
timestamp 1586364061
transform 1 0 3220 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_36
timestamp 1586364061
transform 1 0 4416 0 -1 32096
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5980 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_46
timestamp 1586364061
transform 1 0 5336 0 -1 32096
box -38 -48 590 592
use scs8hd_fill_1  FILLER_54_52
timestamp 1586364061
transform 1 0 5888 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_55
timestamp 1586364061
transform 1 0 6164 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_59
timestamp 1586364061
transform 1 0 6532 0 -1 32096
box -38 -48 314 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 8372 0 -1 32096
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 8188 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_71
timestamp 1586364061
transform 1 0 7636 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_75
timestamp 1586364061
transform 1 0 8004 0 -1 32096
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_82
timestamp 1586364061
transform 1 0 8648 0 -1 32096
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_ipin_13.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11040 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_119
timestamp 1586364061
transform 1 0 12052 0 -1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 12420 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 12788 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_125
timestamp 1586364061
transform 1 0 12604 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_buf_4  mux_right_ipin_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 590 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2300 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2668 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_9
timestamp 1586364061
transform 1 0 1932 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_19
timestamp 1586364061
transform 1 0 2852 0 1 32096
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3036 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4048 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4416 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_30
timestamp 1586364061
transform 1 0 3864 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_34
timestamp 1586364061
transform 1 0 4232 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_38
timestamp 1586364061
transform 1 0 4600 0 1 32096
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6900 0 1 32096
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_1  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9384 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8832 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_82
timestamp 1586364061
transform 1 0 8648 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_99
timestamp 1586364061
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 10948 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 10396 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10764 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_103
timestamp 1586364061
transform 1 0 10580 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_111
timestamp 1586364061
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_55_115
timestamp 1586364061
transform 1 0 11684 0 1 32096
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_fill_1  FILLER_55_121
timestamp 1586364061
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2300 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1656 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2024 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_8
timestamp 1586364061
transform 1 0 1840 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_12
timestamp 1586364061
transform 1 0 2208 0 -1 33184
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3312 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_22
timestamp 1586364061
transform 1 0 3128 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_26
timestamp 1586364061
transform 1 0 3496 0 -1 33184
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5980 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5060 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5796 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5428 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_41
timestamp 1586364061
transform 1 0 4876 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_45
timestamp 1586364061
transform 1 0 5244 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_49
timestamp 1586364061
transform 1 0 5612 0 -1 33184
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l2_in_2_
timestamp 1586364061
transform 1 0 7544 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6992 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_62
timestamp 1586364061
transform 1 0 6808 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_66
timestamp 1586364061
transform 1 0 7176 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_79
timestamp 1586364061
transform 1 0 8372 0 -1 33184
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10120 0 -1 33184
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9844 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8556 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_83
timestamp 1586364061
transform 1 0 8740 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_56_89
timestamp 1586364061
transform 1 0 9292 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_97
timestamp 1586364061
transform 1 0 10028 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_145
timestamp 1586364061
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1564 0 1 33184
box -38 -48 1786 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 1 33184
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3864 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3496 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_24
timestamp 1586364061
transform 1 0 3312 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_28
timestamp 1586364061
transform 1 0 3680 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6992 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_73
timestamp 1586364061
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_77
timestamp 1586364061
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8556 0 1 33184
box -38 -48 1786 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 11040 0 1 33184
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_100
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_104
timestamp 1586364061
transform 1 0 10672 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_112
timestamp 1586364061
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_57_116
timestamp 1586364061
transform 1 0 11776 0 1 33184
box -38 -48 590 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 13432 0 1 33184
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 12696 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 314 592
use scs8hd_decap_6  FILLER_57_128
timestamp 1586364061
transform 1 0 12880 0 1 33184
box -38 -48 590 592
use scs8hd_fill_2  FILLER_57_138
timestamp 1586364061
transform 1 0 13800 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 13984 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_142
timestamp 1586364061
transform 1 0 14168 0 1 33184
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1656 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2668 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_19
timestamp 1586364061
transform 1 0 2852 0 -1 34272
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4324 0 -1 34272
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3036 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_23
timestamp 1586364061
transform 1 0 3220 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_3  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_58_54
timestamp 1586364061
transform 1 0 6072 0 -1 34272
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6808 0 -1 34272
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_81
timestamp 1586364061
transform 1 0 8556 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_85
timestamp 1586364061
transform 1 0 8924 0 -1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_58_91
timestamp 1586364061
transform 1 0 9476 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_112
timestamp 1586364061
transform 1 0 11408 0 -1 34272
box -38 -48 1142 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 12696 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_124
timestamp 1586364061
transform 1 0 12512 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_58_130
timestamp 1586364061
transform 1 0 13064 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_58_142
timestamp 1586364061
transform 1 0 14168 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_7
timestamp 1586364061
transform 1 0 1748 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_7
timestamp 1586364061
transform 1 0 1748 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1840 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_10
timestamp 1586364061
transform 1 0 2024 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2208 0 1 34272
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2116 0 -1 35360
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 1 34272
box -38 -48 866 592
use scs8hd_decap_6  FILLER_60_24
timestamp 1586364061
transform 1 0 3312 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_60_20
timestamp 1586364061
transform 1 0 2944 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_23
timestamp 1586364061
transform 1 0 3220 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_36
timestamp 1586364061
transform 1 0 4416 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_30
timestamp 1586364061
transform 1 0 3864 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3956 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_59_44
timestamp 1586364061
transform 1 0 5152 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_40
timestamp 1586364061
transform 1 0 4784 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5336 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 5520 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4968 0 -1 35360
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_60_65
timestamp 1586364061
transform 1 0 7084 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_61
timestamp 1586364061
transform 1 0 6716 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6900 0 -1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 866 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 7452 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_6  FILLER_60_73
timestamp 1586364061
transform 1 0 7820 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_75
timestamp 1586364061
transform 1 0 8004 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_71
timestamp 1586364061
transform 1 0 7636 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8372 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_ipin_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_81
timestamp 1586364061
transform 1 0 8556 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_59_88
timestamp 1586364061
transform 1 0 9200 0 1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_60_97
timestamp 1586364061
transform 1 0 10028 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_3  FILLER_60_89
timestamp 1586364061
transform 1 0 9292 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_59_92
timestamp 1586364061
transform 1 0 9568 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 9936 0 1 34272
box -38 -48 406 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_104
timestamp 1586364061
transform 1 0 10672 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_100
timestamp 1586364061
transform 1 0 10304 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 10488 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 10856 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 406 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 11040 0 1 34272
box -38 -48 406 592
use scs8hd_decap_4  FILLER_60_113
timestamp 1586364061
transform 1 0 11500 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_109
timestamp 1586364061
transform 1 0 11132 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_112
timestamp 1586364061
transform 1 0 11408 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 11316 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_116
timestamp 1586364061
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_8  FILLER_60_121
timestamp 1586364061
transform 1 0 12236 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_8  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_120
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_135
timestamp 1586364061
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_133
timestamp 1586364061
transform 1 0 13340 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 13156 0 -1 35360
box -38 -48 406 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 13432 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_138
timestamp 1586364061
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_142
timestamp 1586364061
transform 1 0 14168 0 1 34272
box -38 -48 406 592
use scs8hd_decap_3  FILLER_60_143
timestamp 1586364061
transform 1 0 14260 0 -1 35360
box -38 -48 314 592
use scs8hd_buf_4  mux_right_ipin_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 590 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2116 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_9
timestamp 1586364061
transform 1 0 1932 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_13
timestamp 1586364061
transform 1 0 2300 0 1 35360
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_ipin_15.mux_l2_in_3_
timestamp 1586364061
transform 1 0 3956 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3772 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3404 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_40
timestamp 1586364061
transform 1 0 4784 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_52
timestamp 1586364061
transform 1 0 5888 0 1 35360
box -38 -48 774 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 7820 0 1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 8372 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_60
timestamp 1586364061
transform 1 0 6624 0 1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  FILLER_61_70
timestamp 1586364061
transform 1 0 7544 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_77
timestamp 1586364061
transform 1 0 8188 0 1 35360
box -38 -48 222 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 8924 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 9476 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 9844 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_81
timestamp 1586364061
transform 1 0 8556 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_89
timestamp 1586364061
transform 1 0 9292 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_93
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 11132 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 10764 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 11868 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_101
timestamp 1586364061
transform 1 0 10396 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_107
timestamp 1586364061
transform 1 0 10948 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_113
timestamp 1586364061
transform 1 0 11500 0 1 35360
box -38 -48 406 592
use scs8hd_decap_3  FILLER_61_119
timestamp 1586364061
transform 1 0 12052 0 1 35360
box -38 -48 314 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 12972 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_127
timestamp 1586364061
transform 1 0 12788 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_131
timestamp 1586364061
transform 1 0 13156 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4232 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_36
timestamp 1586364061
transform 1 0 4416 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_48
timestamp 1586364061
transform 1 0 5520 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_60
timestamp 1586364061
transform 1 0 6624 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_72
timestamp 1586364061
transform 1 0 7728 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_84
timestamp 1586364061
transform 1 0 8832 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 406 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_8  FILLER_62_109
timestamp 1586364061
transform 1 0 11132 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_12  FILLER_62_121
timestamp 1586364061
transform 1 0 12236 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_133
timestamp 1586364061
transform 1 0 13340 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 774 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 11132 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 11684 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_106
timestamp 1586364061
transform 1 0 10856 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_113
timestamp 1586364061
transform 1 0 11500 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_117
timestamp 1586364061
transform 1 0 11868 0 1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_63_121
timestamp 1586364061
transform 1 0 12236 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 15750 39520 15806 40000 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 38632 480 38752 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 570 0 626 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 202 39520 258 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 4066 39520 4122 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 4434 39520 4490 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 4802 39520 4858 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 5262 39520 5318 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 5630 39520 5686 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 5998 39520 6054 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 6366 39520 6422 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 6826 39520 6882 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 7194 39520 7250 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 7562 39520 7618 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 570 39520 626 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 938 39520 994 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 1306 39520 1362 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 1674 39520 1730 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 2502 39520 2558 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 2870 39520 2926 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 3238 39520 3294 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 3698 39520 3754 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 7930 39520 7986 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 11886 39520 11942 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 12254 39520 12310 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 12622 39520 12678 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 13082 39520 13138 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 13450 39520 13506 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 13818 39520 13874 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 14646 39520 14702 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 15014 39520 15070 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 8390 39520 8446 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 8758 39520 8814 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 9126 39520 9182 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 9494 39520 9550 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 9954 39520 10010 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 10322 39520 10378 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 10690 39520 10746 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 11058 39520 11114 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 11518 39520 11574 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 1096 480 1216 6 left_grid_pin_0_
port 82 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 left_grid_pin_10_
port 83 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_11_
port 84 nsew default tristate
rlabel metal3 s 0 29248 480 29368 6 left_grid_pin_12_
port 85 nsew default tristate
rlabel metal3 s 0 31560 480 31680 6 left_grid_pin_13_
port 86 nsew default tristate
rlabel metal3 s 0 34008 480 34128 6 left_grid_pin_14_
port 87 nsew default tristate
rlabel metal3 s 0 36320 480 36440 6 left_grid_pin_15_
port 88 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_1_
port 89 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 left_grid_pin_2_
port 90 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_3_
port 91 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 left_grid_pin_4_
port 92 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_5_
port 93 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_6_
port 94 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_7_
port 95 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 left_grid_pin_8_
port 96 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 left_grid_pin_9_
port 97 nsew default tristate
rlabel metal3 s 15520 29928 16000 30048 6 prog_clk
port 98 nsew default input
rlabel metal3 s 15520 9936 16000 10056 6 right_grid_pin_52_
port 99 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 100 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
