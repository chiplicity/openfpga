magic
tech sky130A
magscale 1 2
timestamp 1606928588
<< locali >>
rect 7941 13855 7975 14025
rect 13277 11611 13311 11849
rect 13553 9979 13587 10081
rect 10517 8959 10551 9061
rect 10183 8517 10275 8551
rect 6561 8347 6595 8449
rect 10241 8415 10275 8517
rect 3893 7803 3927 8041
rect 13093 7191 13127 7293
rect 8769 6103 8803 6409
rect 8493 5627 8527 5729
rect 7665 5151 7699 5321
rect 10149 4607 10183 4777
rect 3525 2907 3559 3145
rect 3617 2839 3651 3077
rect 6561 2907 6595 3145
rect 7481 2907 7515 3009
<< viali >>
rect 2513 14569 2547 14603
rect 5457 14569 5491 14603
rect 1593 14433 1627 14467
rect 2329 14433 2363 14467
rect 5273 14433 5307 14467
rect 1777 14365 1811 14399
rect 5181 14229 5215 14263
rect 3249 14025 3283 14059
rect 4077 14025 4111 14059
rect 7941 14025 7975 14059
rect 17601 14025 17635 14059
rect 18245 14025 18279 14059
rect 2605 13889 2639 13923
rect 6377 13889 6411 13923
rect 7573 13889 7607 13923
rect 17049 13957 17083 13991
rect 8309 13889 8343 13923
rect 14381 13889 14415 13923
rect 1593 13821 1627 13855
rect 1869 13821 1903 13855
rect 2329 13821 2363 13855
rect 3065 13821 3099 13855
rect 3893 13821 3927 13855
rect 6193 13821 6227 13855
rect 7941 13821 7975 13855
rect 8033 13821 8067 13855
rect 14115 13821 14149 13855
rect 16865 13821 16899 13855
rect 17417 13821 17451 13855
rect 18061 13821 18095 13855
rect 6101 13753 6135 13787
rect 5733 13685 5767 13719
rect 7021 13685 7055 13719
rect 7389 13685 7423 13719
rect 7481 13685 7515 13719
rect 2513 13481 2547 13515
rect 5273 13481 5307 13515
rect 6929 13481 6963 13515
rect 7389 13481 7423 13515
rect 1869 13413 1903 13447
rect 1593 13345 1627 13379
rect 2329 13345 2363 13379
rect 6285 13345 6319 13379
rect 7297 13345 7331 13379
rect 8769 13345 8803 13379
rect 10885 13345 10919 13379
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 6377 13277 6411 13311
rect 6469 13277 6503 13311
rect 7573 13277 7607 13311
rect 8861 13277 8895 13311
rect 8953 13277 8987 13311
rect 10977 13277 11011 13311
rect 11069 13277 11103 13311
rect 5917 13209 5951 13243
rect 8401 13209 8435 13243
rect 4905 13141 4939 13175
rect 10517 13141 10551 13175
rect 1869 12937 1903 12971
rect 5733 12937 5767 12971
rect 6837 12937 6871 12971
rect 3249 12869 3283 12903
rect 2789 12801 2823 12835
rect 3801 12801 3835 12835
rect 4905 12801 4939 12835
rect 6377 12801 6411 12835
rect 7481 12801 7515 12835
rect 8585 12801 8619 12835
rect 10333 12801 10367 12835
rect 10517 12801 10551 12835
rect 11529 12801 11563 12835
rect 12817 12801 12851 12835
rect 1685 12733 1719 12767
rect 4813 12733 4847 12767
rect 12449 12733 12483 12767
rect 6101 12665 6135 12699
rect 7205 12665 7239 12699
rect 11345 12665 11379 12699
rect 2237 12597 2271 12631
rect 2605 12597 2639 12631
rect 2697 12597 2731 12631
rect 3617 12597 3651 12631
rect 3709 12597 3743 12631
rect 4353 12597 4387 12631
rect 4721 12597 4755 12631
rect 6193 12597 6227 12631
rect 7297 12597 7331 12631
rect 7941 12597 7975 12631
rect 8309 12597 8343 12631
rect 8401 12597 8435 12631
rect 9873 12597 9907 12631
rect 10241 12597 10275 12631
rect 10885 12597 10919 12631
rect 11253 12597 11287 12631
rect 1777 12393 1811 12427
rect 4077 12393 4111 12427
rect 4537 12393 4571 12427
rect 5089 12393 5123 12427
rect 5457 12393 5491 12427
rect 6101 12393 6135 12427
rect 6469 12393 6503 12427
rect 7481 12393 7515 12427
rect 10793 12393 10827 12427
rect 11345 12393 11379 12427
rect 16129 12393 16163 12427
rect 17601 12393 17635 12427
rect 3157 12325 3191 12359
rect 8401 12325 8435 12359
rect 8493 12325 8527 12359
rect 17509 12325 17543 12359
rect 2145 12257 2179 12291
rect 3249 12257 3283 12291
rect 4445 12257 4479 12291
rect 6561 12257 6595 12291
rect 10701 12257 10735 12291
rect 11713 12257 11747 12291
rect 2237 12189 2271 12223
rect 2421 12189 2455 12223
rect 3341 12189 3375 12223
rect 4629 12189 4663 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 6653 12189 6687 12223
rect 8677 12189 8711 12223
rect 10977 12189 11011 12223
rect 11805 12189 11839 12223
rect 11897 12189 11931 12223
rect 16221 12189 16255 12223
rect 16313 12189 16347 12223
rect 17693 12189 17727 12223
rect 18153 12189 18187 12223
rect 2789 12053 2823 12087
rect 8033 12053 8067 12087
rect 10333 12053 10367 12087
rect 15761 12053 15795 12087
rect 17141 12053 17175 12087
rect 6469 11849 6503 11883
rect 11529 11849 11563 11883
rect 13277 11849 13311 11883
rect 13369 11849 13403 11883
rect 4353 11713 4387 11747
rect 8493 11713 8527 11747
rect 2053 11645 2087 11679
rect 2320 11645 2354 11679
rect 4169 11645 4203 11679
rect 5089 11645 5123 11679
rect 6837 11645 6871 11679
rect 7093 11645 7127 11679
rect 10149 11645 10183 11679
rect 13921 11713 13955 11747
rect 16497 11713 16531 11747
rect 16681 11713 16715 11747
rect 13737 11645 13771 11679
rect 14381 11645 14415 11679
rect 17417 11645 17451 11679
rect 18061 11645 18095 11679
rect 5356 11577 5390 11611
rect 8760 11577 8794 11611
rect 10394 11577 10428 11611
rect 13277 11577 13311 11611
rect 14648 11577 14682 11611
rect 16405 11577 16439 11611
rect 3433 11509 3467 11543
rect 3801 11509 3835 11543
rect 4261 11509 4295 11543
rect 8217 11509 8251 11543
rect 9873 11509 9907 11543
rect 11805 11509 11839 11543
rect 13829 11509 13863 11543
rect 15761 11509 15795 11543
rect 16037 11509 16071 11543
rect 17601 11509 17635 11543
rect 18245 11509 18279 11543
rect 2053 11305 2087 11339
rect 2421 11305 2455 11339
rect 5457 11305 5491 11339
rect 5733 11305 5767 11339
rect 6193 11305 6227 11339
rect 8033 11305 8067 11339
rect 8953 11305 8987 11339
rect 9689 11305 9723 11339
rect 10057 11305 10091 11339
rect 10885 11305 10919 11339
rect 11253 11305 11287 11339
rect 11345 11305 11379 11339
rect 17693 11305 17727 11339
rect 1961 11237 1995 11271
rect 17785 11237 17819 11271
rect 2513 11169 2547 11203
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 6101 11169 6135 11203
rect 7941 11169 7975 11203
rect 12265 11169 12299 11203
rect 13093 11169 13127 11203
rect 13360 11169 13394 11203
rect 15925 11169 15959 11203
rect 2605 11101 2639 11135
rect 3065 11101 3099 11135
rect 6285 11101 6319 11135
rect 8217 11101 8251 11135
rect 9045 11101 9079 11135
rect 9229 11101 9263 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11529 11101 11563 11135
rect 12357 11101 12391 11135
rect 12541 11101 12575 11135
rect 15669 11101 15703 11135
rect 17877 11101 17911 11135
rect 7573 11033 7607 11067
rect 8585 11033 8619 11067
rect 11897 10965 11931 10999
rect 14473 10965 14507 10999
rect 17049 10965 17083 10999
rect 17325 10965 17359 10999
rect 2053 10761 2087 10795
rect 3065 10761 3099 10795
rect 4261 10761 4295 10795
rect 5273 10761 5307 10795
rect 7113 10761 7147 10795
rect 8769 10761 8803 10795
rect 9229 10761 9263 10795
rect 11621 10761 11655 10795
rect 14105 10761 14139 10795
rect 14381 10761 14415 10795
rect 1685 10693 1719 10727
rect 2697 10625 2731 10659
rect 3525 10625 3559 10659
rect 3617 10625 3651 10659
rect 4813 10625 4847 10659
rect 5917 10625 5951 10659
rect 9781 10625 9815 10659
rect 10241 10625 10275 10659
rect 15025 10625 15059 10659
rect 16037 10625 16071 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 1501 10557 1535 10591
rect 2421 10557 2455 10591
rect 4629 10557 4663 10591
rect 5733 10557 5767 10591
rect 7297 10557 7331 10591
rect 7389 10557 7423 10591
rect 7656 10557 7690 10591
rect 10508 10557 10542 10591
rect 12449 10557 12483 10591
rect 14289 10557 14323 10591
rect 14841 10557 14875 10591
rect 15853 10557 15887 10591
rect 16957 10557 16991 10591
rect 18061 10557 18095 10591
rect 2513 10489 2547 10523
rect 9597 10489 9631 10523
rect 12716 10489 12750 10523
rect 14749 10489 14783 10523
rect 15761 10489 15795 10523
rect 3433 10421 3467 10455
rect 4721 10421 4755 10455
rect 5641 10421 5675 10455
rect 9689 10421 9723 10455
rect 13829 10421 13863 10455
rect 15393 10421 15427 10455
rect 16589 10421 16623 10455
rect 18245 10421 18279 10455
rect 3617 10217 3651 10251
rect 7113 10217 7147 10251
rect 9873 10217 9907 10251
rect 10885 10217 10919 10251
rect 13277 10217 13311 10251
rect 14197 10217 14231 10251
rect 14657 10217 14691 10251
rect 17325 10217 17359 10251
rect 18153 10217 18187 10251
rect 1676 10149 1710 10183
rect 6000 10149 6034 10183
rect 8197 10149 8231 10183
rect 10241 10149 10275 10183
rect 17417 10149 17451 10183
rect 3065 10081 3099 10115
rect 3801 10081 3835 10115
rect 4445 10081 4479 10115
rect 5733 10081 5767 10115
rect 7941 10081 7975 10115
rect 11069 10081 11103 10115
rect 11529 10081 11563 10115
rect 11888 10081 11922 10115
rect 13461 10081 13495 10115
rect 13553 10081 13587 10115
rect 14565 10081 14599 10115
rect 15301 10081 15335 10115
rect 15568 10081 15602 10115
rect 17969 10081 18003 10115
rect 1409 10013 1443 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 5089 10013 5123 10047
rect 7481 10013 7515 10047
rect 10333 10013 10367 10047
rect 10517 10013 10551 10047
rect 11621 10013 11655 10047
rect 13737 10013 13771 10047
rect 14749 10013 14783 10047
rect 17509 10013 17543 10047
rect 2789 9945 2823 9979
rect 4077 9945 4111 9979
rect 9321 9945 9355 9979
rect 13553 9945 13587 9979
rect 3249 9877 3283 9911
rect 11345 9877 11379 9911
rect 13001 9877 13035 9911
rect 16681 9877 16715 9911
rect 16957 9877 16991 9911
rect 3617 9673 3651 9707
rect 16957 9673 16991 9707
rect 6285 9605 6319 9639
rect 8677 9605 8711 9639
rect 11069 9605 11103 9639
rect 11345 9605 11379 9639
rect 4077 9537 4111 9571
rect 4261 9537 4295 9571
rect 6837 9537 6871 9571
rect 9321 9537 9355 9571
rect 9689 9537 9723 9571
rect 11989 9537 12023 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 15025 9537 15059 9571
rect 15577 9537 15611 9571
rect 1777 9469 1811 9503
rect 4629 9469 4663 9503
rect 4896 9469 4930 9503
rect 6469 9469 6503 9503
rect 9956 9469 9990 9503
rect 14841 9469 14875 9503
rect 15844 9469 15878 9503
rect 17417 9469 17451 9503
rect 18061 9469 18095 9503
rect 2044 9401 2078 9435
rect 3985 9401 4019 9435
rect 7104 9401 7138 9435
rect 9137 9401 9171 9435
rect 12817 9401 12851 9435
rect 13829 9401 13863 9435
rect 14933 9401 14967 9435
rect 3157 9333 3191 9367
rect 6009 9333 6043 9367
rect 8217 9333 8251 9367
rect 9045 9333 9079 9367
rect 11713 9333 11747 9367
rect 11805 9333 11839 9367
rect 12449 9333 12483 9367
rect 13461 9333 13495 9367
rect 14473 9333 14507 9367
rect 17601 9333 17635 9367
rect 18245 9333 18279 9367
rect 5457 9129 5491 9163
rect 7389 9129 7423 9163
rect 9321 9129 9355 9163
rect 9689 9129 9723 9163
rect 12081 9129 12115 9163
rect 12541 9129 12575 9163
rect 14933 9129 14967 9163
rect 1676 9061 1710 9095
rect 8208 9061 8242 9095
rect 10517 9061 10551 9095
rect 10968 9061 11002 9095
rect 16764 9061 16798 9095
rect 1409 8993 1443 9027
rect 3065 8993 3099 9027
rect 4077 8993 4111 9027
rect 4344 8993 4378 9027
rect 6009 8993 6043 9027
rect 6276 8993 6310 9027
rect 7941 8993 7975 9027
rect 10057 8993 10091 9027
rect 12909 8993 12943 9027
rect 13553 8993 13587 9027
rect 13820 8993 13854 9027
rect 15853 8993 15887 9027
rect 15945 8993 15979 9027
rect 16497 8993 16531 9027
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 13001 8925 13035 8959
rect 13185 8925 13219 8959
rect 16129 8925 16163 8959
rect 2789 8789 2823 8823
rect 3249 8789 3283 8823
rect 15485 8789 15519 8823
rect 17877 8789 17911 8823
rect 1409 8585 1443 8619
rect 3801 8585 3835 8619
rect 4721 8585 4755 8619
rect 7021 8585 7055 8619
rect 8309 8585 8343 8619
rect 12633 8585 12667 8619
rect 16497 8585 16531 8619
rect 5733 8517 5767 8551
rect 9321 8517 9355 8551
rect 10149 8517 10183 8551
rect 10333 8517 10367 8551
rect 11345 8517 11379 8551
rect 18245 8517 18279 8551
rect 1869 8449 1903 8483
rect 2053 8449 2087 8483
rect 2421 8449 2455 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 8953 8449 8987 8483
rect 9965 8449 9999 8483
rect 1777 8381 1811 8415
rect 4077 8381 4111 8415
rect 5089 8381 5123 8415
rect 6101 8381 6135 8415
rect 6193 8381 6227 8415
rect 10793 8449 10827 8483
rect 10977 8449 11011 8483
rect 11989 8449 12023 8483
rect 13093 8449 13127 8483
rect 13277 8449 13311 8483
rect 14473 8449 14507 8483
rect 14841 8449 14875 8483
rect 16957 8449 16991 8483
rect 17049 8449 17083 8483
rect 8769 8381 8803 8415
rect 9781 8381 9815 8415
rect 10241 8381 10275 8415
rect 10701 8381 10735 8415
rect 11805 8381 11839 8415
rect 13001 8381 13035 8415
rect 14289 8381 14323 8415
rect 15108 8381 15142 8415
rect 18061 8381 18095 8415
rect 2666 8313 2700 8347
rect 6561 8313 6595 8347
rect 7389 8313 7423 8347
rect 9689 8313 9723 8347
rect 4261 8245 4295 8279
rect 8677 8245 8711 8279
rect 11713 8245 11747 8279
rect 13829 8245 13863 8279
rect 14197 8245 14231 8279
rect 16221 8245 16255 8279
rect 16865 8245 16899 8279
rect 17509 8245 17543 8279
rect 1593 8041 1627 8075
rect 3433 8041 3467 8075
rect 3893 8041 3927 8075
rect 5273 8041 5307 8075
rect 6653 8041 6687 8075
rect 6745 8041 6779 8075
rect 10333 8041 10367 8075
rect 14381 8041 14415 8075
rect 14841 8041 14875 8075
rect 15853 8041 15887 8075
rect 16405 8041 16439 8075
rect 16773 8041 16807 8075
rect 17417 8041 17451 8075
rect 17785 8041 17819 8075
rect 2329 7973 2363 8007
rect 1409 7905 1443 7939
rect 3341 7905 3375 7939
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 3617 7837 3651 7871
rect 5641 7973 5675 8007
rect 9689 7973 9723 8007
rect 15761 7973 15795 8007
rect 4629 7905 4663 7939
rect 7297 7905 7331 7939
rect 7849 7905 7883 7939
rect 8116 7905 8150 7939
rect 10701 7905 10735 7939
rect 11345 7905 11379 7939
rect 11612 7905 11646 7939
rect 13257 7905 13291 7939
rect 14657 7905 14691 7939
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 6837 7837 6871 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 13001 7837 13035 7871
rect 16037 7837 16071 7871
rect 16865 7837 16899 7871
rect 16957 7837 16991 7871
rect 17877 7837 17911 7871
rect 17969 7837 18003 7871
rect 3893 7769 3927 7803
rect 6285 7769 6319 7803
rect 12725 7769 12759 7803
rect 1961 7701 1995 7735
rect 2973 7701 3007 7735
rect 4261 7701 4295 7735
rect 7481 7701 7515 7735
rect 9229 7701 9263 7735
rect 15393 7701 15427 7735
rect 1685 7497 1719 7531
rect 3709 7497 3743 7531
rect 6101 7497 6135 7531
rect 11069 7497 11103 7531
rect 12081 7497 12115 7531
rect 16221 7497 16255 7531
rect 16957 7497 16991 7531
rect 2237 7361 2271 7395
rect 3341 7361 3375 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 4721 7361 4755 7395
rect 7389 7361 7423 7395
rect 10701 7361 10735 7395
rect 11713 7361 11747 7395
rect 13829 7361 13863 7395
rect 17601 7361 17635 7395
rect 2053 7293 2087 7327
rect 3065 7293 3099 7327
rect 6653 7293 6687 7327
rect 7849 7293 7883 7327
rect 8953 7293 8987 7327
rect 11897 7293 11931 7327
rect 12725 7293 12759 7327
rect 13093 7293 13127 7327
rect 13645 7293 13679 7327
rect 14289 7293 14323 7327
rect 14841 7293 14875 7327
rect 16497 7293 16531 7327
rect 17325 7293 17359 7327
rect 18061 7293 18095 7327
rect 4077 7225 4111 7259
rect 4988 7225 5022 7259
rect 7205 7225 7239 7259
rect 11437 7225 11471 7259
rect 13737 7225 13771 7259
rect 15108 7225 15142 7259
rect 17417 7225 17451 7259
rect 2145 7157 2179 7191
rect 2697 7157 2731 7191
rect 3157 7157 3191 7191
rect 6469 7157 6503 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 8033 7157 8067 7191
rect 11529 7157 11563 7191
rect 12909 7157 12943 7191
rect 13093 7157 13127 7191
rect 13277 7157 13311 7191
rect 14473 7157 14507 7191
rect 18245 7157 18279 7191
rect 10241 6953 10275 6987
rect 14933 6953 14967 6987
rect 17785 6953 17819 6987
rect 8392 6885 8426 6919
rect 11152 6885 11186 6919
rect 16028 6885 16062 6919
rect 1941 6817 1975 6851
rect 3341 6817 3375 6851
rect 4804 6817 4838 6851
rect 6552 6817 6586 6851
rect 12909 6817 12943 6851
rect 13809 6817 13843 6851
rect 15761 6817 15795 6851
rect 1685 6749 1719 6783
rect 4077 6749 4111 6783
rect 4537 6749 4571 6783
rect 6285 6749 6319 6783
rect 8125 6749 8159 6783
rect 10333 6749 10367 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 13001 6749 13035 6783
rect 13185 6749 13219 6783
rect 13553 6749 13587 6783
rect 15301 6749 15335 6783
rect 17877 6749 17911 6783
rect 17969 6749 18003 6783
rect 3065 6681 3099 6715
rect 12265 6681 12299 6715
rect 17417 6681 17451 6715
rect 3525 6613 3559 6647
rect 5917 6613 5951 6647
rect 7665 6613 7699 6647
rect 9505 6613 9539 6647
rect 9873 6613 9907 6647
rect 12541 6613 12575 6647
rect 17141 6613 17175 6647
rect 4445 6409 4479 6443
rect 8769 6409 8803 6443
rect 11161 6409 11195 6443
rect 12817 6409 12851 6443
rect 15853 6409 15887 6443
rect 7941 6341 7975 6375
rect 2697 6273 2731 6307
rect 5641 6273 5675 6307
rect 6377 6273 6411 6307
rect 6469 6273 6503 6307
rect 7665 6273 7699 6307
rect 8493 6273 8527 6307
rect 1501 6205 1535 6239
rect 2421 6205 2455 6239
rect 3065 6205 3099 6239
rect 4997 6205 5031 6239
rect 7481 6205 7515 6239
rect 7573 6205 7607 6239
rect 8309 6205 8343 6239
rect 3332 6137 3366 6171
rect 5457 6137 5491 6171
rect 13829 6341 13863 6375
rect 8861 6273 8895 6307
rect 11713 6273 11747 6307
rect 13277 6273 13311 6307
rect 13461 6273 13495 6307
rect 14289 6273 14323 6307
rect 14473 6273 14507 6307
rect 15301 6273 15335 6307
rect 15485 6273 15519 6307
rect 16313 6273 16347 6307
rect 16497 6273 16531 6307
rect 17325 6273 17359 6307
rect 17509 6273 17543 6307
rect 9128 6205 9162 6239
rect 10517 6205 10551 6239
rect 18061 6205 18095 6239
rect 11621 6137 11655 6171
rect 15209 6137 15243 6171
rect 1685 6069 1719 6103
rect 2053 6069 2087 6103
rect 2513 6069 2547 6103
rect 4813 6069 4847 6103
rect 5089 6069 5123 6103
rect 5549 6069 5583 6103
rect 5917 6069 5951 6103
rect 6285 6069 6319 6103
rect 7113 6069 7147 6103
rect 8401 6069 8435 6103
rect 8769 6069 8803 6103
rect 10241 6069 10275 6103
rect 11529 6069 11563 6103
rect 13185 6069 13219 6103
rect 14197 6069 14231 6103
rect 14841 6069 14875 6103
rect 16221 6069 16255 6103
rect 16865 6069 16899 6103
rect 17233 6069 17267 6103
rect 18245 6069 18279 6103
rect 2237 5865 2271 5899
rect 5733 5865 5767 5899
rect 6101 5865 6135 5899
rect 8401 5865 8435 5899
rect 9137 5865 9171 5899
rect 11069 5865 11103 5899
rect 11897 5865 11931 5899
rect 12909 5865 12943 5899
rect 15669 5865 15703 5899
rect 15761 5865 15795 5899
rect 18153 5865 18187 5899
rect 4344 5797 4378 5831
rect 13544 5797 13578 5831
rect 1685 5729 1719 5763
rect 2605 5729 2639 5763
rect 3249 5729 3283 5763
rect 6561 5729 6595 5763
rect 7288 5729 7322 5763
rect 8493 5729 8527 5763
rect 8585 5729 8619 5763
rect 8953 5729 8987 5763
rect 9945 5729 9979 5763
rect 12725 5729 12759 5763
rect 13277 5729 13311 5763
rect 15117 5729 15151 5763
rect 16753 5729 16787 5763
rect 2697 5661 2731 5695
rect 2881 5661 2915 5695
rect 4077 5661 4111 5695
rect 6193 5661 6227 5695
rect 6377 5661 6411 5695
rect 7021 5661 7055 5695
rect 9689 5661 9723 5695
rect 11989 5661 12023 5695
rect 12173 5661 12207 5695
rect 15945 5661 15979 5695
rect 16497 5661 16531 5695
rect 8493 5593 8527 5627
rect 1869 5525 1903 5559
rect 3433 5525 3467 5559
rect 5457 5525 5491 5559
rect 6745 5525 6779 5559
rect 8769 5525 8803 5559
rect 11529 5525 11563 5559
rect 14657 5525 14691 5559
rect 14933 5525 14967 5559
rect 15301 5525 15335 5559
rect 17877 5525 17911 5559
rect 6837 5321 6871 5355
rect 7665 5321 7699 5355
rect 10149 5321 10183 5355
rect 14473 5321 14507 5355
rect 14749 5321 14783 5355
rect 2329 5185 2363 5219
rect 4905 5185 4939 5219
rect 7389 5185 7423 5219
rect 8953 5253 8987 5287
rect 8309 5185 8343 5219
rect 8401 5185 8435 5219
rect 9505 5185 9539 5219
rect 10793 5185 10827 5219
rect 11805 5185 11839 5219
rect 15025 5185 15059 5219
rect 17509 5185 17543 5219
rect 1593 5117 1627 5151
rect 4169 5117 4203 5151
rect 5172 5117 5206 5151
rect 7665 5117 7699 5151
rect 9413 5117 9447 5151
rect 10517 5117 10551 5151
rect 11529 5117 11563 5151
rect 13093 5117 13127 5151
rect 14933 5117 14967 5151
rect 15292 5117 15326 5151
rect 18061 5117 18095 5151
rect 1869 5049 1903 5083
rect 2596 5049 2630 5083
rect 4445 5049 4479 5083
rect 9321 5049 9355 5083
rect 10609 5049 10643 5083
rect 13360 5049 13394 5083
rect 3709 4981 3743 5015
rect 6285 4981 6319 5015
rect 7205 4981 7239 5015
rect 7297 4981 7331 5015
rect 7849 4981 7883 5015
rect 8217 4981 8251 5015
rect 11161 4981 11195 5015
rect 11621 4981 11655 5015
rect 12449 4981 12483 5015
rect 16405 4981 16439 5015
rect 16957 4981 16991 5015
rect 17325 4981 17359 5015
rect 17417 4981 17451 5015
rect 18245 4981 18279 5015
rect 2973 4777 3007 4811
rect 4537 4777 4571 4811
rect 5089 4777 5123 4811
rect 6101 4777 6135 4811
rect 9045 4777 9079 4811
rect 9873 4777 9907 4811
rect 10149 4777 10183 4811
rect 10977 4777 11011 4811
rect 11529 4777 11563 4811
rect 14013 4777 14047 4811
rect 15669 4777 15703 4811
rect 16681 4777 16715 4811
rect 17509 4777 17543 4811
rect 2421 4709 2455 4743
rect 1409 4641 1443 4675
rect 2329 4641 2363 4675
rect 3341 4641 3375 4675
rect 4445 4641 4479 4675
rect 5457 4641 5491 4675
rect 6285 4641 6319 4675
rect 6633 4641 6667 4675
rect 8033 4641 8067 4675
rect 8953 4641 8987 4675
rect 9689 4641 9723 4675
rect 11897 4709 11931 4743
rect 17417 4709 17451 4743
rect 10425 4641 10459 4675
rect 10885 4641 10919 4675
rect 12889 4641 12923 4675
rect 14657 4641 14691 4675
rect 16497 4641 16531 4675
rect 18061 4641 18095 4675
rect 2513 4573 2547 4607
rect 3433 4573 3467 4607
rect 3617 4573 3651 4607
rect 4629 4573 4663 4607
rect 5549 4573 5583 4607
rect 5641 4573 5675 4607
rect 6377 4573 6411 4607
rect 9229 4573 9263 4607
rect 10149 4573 10183 4607
rect 11161 4573 11195 4607
rect 11989 4573 12023 4607
rect 12173 4573 12207 4607
rect 12633 4573 12667 4607
rect 15761 4573 15795 4607
rect 15853 4573 15887 4607
rect 17601 4573 17635 4607
rect 1961 4505 1995 4539
rect 7757 4505 7791 4539
rect 10517 4505 10551 4539
rect 14841 4505 14875 4539
rect 1593 4437 1627 4471
rect 4077 4437 4111 4471
rect 8217 4437 8251 4471
rect 8585 4437 8619 4471
rect 10241 4437 10275 4471
rect 15301 4437 15335 4471
rect 17049 4437 17083 4471
rect 18245 4437 18279 4471
rect 2789 4233 2823 4267
rect 13829 4233 13863 4267
rect 15945 4233 15979 4267
rect 1409 4097 1443 4131
rect 3985 4097 4019 4131
rect 6193 4097 6227 4131
rect 7389 4097 7423 4131
rect 10517 4097 10551 4131
rect 12449 4097 12483 4131
rect 14289 4097 14323 4131
rect 16497 4097 16531 4131
rect 17417 4097 17451 4131
rect 17601 4097 17635 4131
rect 3249 4029 3283 4063
rect 3525 4029 3559 4063
rect 6101 4029 6135 4063
rect 7297 4029 7331 4063
rect 7849 4029 7883 4063
rect 8401 4029 8435 4063
rect 14556 4029 14590 4063
rect 17325 4029 17359 4063
rect 18061 4029 18095 4063
rect 1654 3961 1688 3995
rect 4252 3961 4286 3995
rect 6009 3961 6043 3995
rect 8668 3961 8702 3995
rect 10762 3961 10796 3995
rect 12716 3961 12750 3995
rect 16313 3961 16347 3995
rect 5365 3893 5399 3927
rect 5641 3893 5675 3927
rect 6837 3893 6871 3927
rect 7205 3893 7239 3927
rect 8033 3893 8067 3927
rect 9781 3893 9815 3927
rect 10057 3893 10091 3927
rect 11897 3893 11931 3927
rect 15669 3893 15703 3927
rect 16405 3893 16439 3927
rect 16957 3893 16991 3927
rect 18245 3893 18279 3927
rect 2145 3689 2179 3723
rect 4997 3689 5031 3723
rect 7389 3689 7423 3723
rect 10149 3689 10183 3723
rect 10977 3689 11011 3723
rect 11989 3689 12023 3723
rect 12357 3689 12391 3723
rect 12449 3689 12483 3723
rect 13921 3689 13955 3723
rect 14381 3689 14415 3723
rect 1685 3621 1719 3655
rect 5089 3621 5123 3655
rect 7932 3621 7966 3655
rect 14289 3621 14323 3655
rect 17325 3621 17359 3655
rect 1409 3553 1443 3587
rect 2513 3553 2547 3587
rect 3157 3553 3191 3587
rect 4077 3553 4111 3587
rect 5989 3553 6023 3587
rect 7573 3553 7607 3587
rect 7665 3553 7699 3587
rect 10057 3553 10091 3587
rect 11345 3553 11379 3587
rect 13001 3553 13035 3587
rect 15301 3553 15335 3587
rect 16313 3553 16347 3587
rect 17049 3553 17083 3587
rect 17785 3553 17819 3587
rect 2605 3485 2639 3519
rect 2697 3485 2731 3519
rect 3433 3485 3467 3519
rect 5273 3485 5307 3519
rect 5733 3485 5767 3519
rect 10241 3485 10275 3519
rect 11437 3485 11471 3519
rect 11529 3485 11563 3519
rect 12541 3485 12575 3519
rect 13185 3485 13219 3519
rect 14565 3485 14599 3519
rect 15577 3485 15611 3519
rect 16589 3485 16623 3519
rect 18061 3485 18095 3519
rect 4261 3417 4295 3451
rect 4629 3349 4663 3383
rect 7113 3349 7147 3383
rect 9045 3349 9079 3383
rect 9689 3349 9723 3383
rect 1685 3145 1719 3179
rect 3525 3145 3559 3179
rect 2329 3009 2363 3043
rect 3249 3009 3283 3043
rect 6561 3145 6595 3179
rect 8585 3145 8619 3179
rect 9597 3145 9631 3179
rect 12449 3145 12483 3179
rect 13461 3145 13495 3179
rect 18245 3145 18279 3179
rect 3157 2873 3191 2907
rect 3525 2873 3559 2907
rect 3617 3077 3651 3111
rect 4261 3009 4295 3043
rect 5273 3009 5307 3043
rect 6285 3009 6319 3043
rect 4077 2941 4111 2975
rect 5181 2941 5215 2975
rect 7573 3077 7607 3111
rect 7481 3009 7515 3043
rect 8033 3009 8067 3043
rect 8217 3009 8251 3043
rect 9045 3009 9079 3043
rect 9137 3009 9171 3043
rect 10149 3009 10183 3043
rect 11069 3009 11103 3043
rect 11253 3009 11287 3043
rect 13001 3009 13035 3043
rect 14013 3009 14047 3043
rect 14657 3009 14691 3043
rect 17509 3009 17543 3043
rect 6837 2941 6871 2975
rect 7941 2941 7975 2975
rect 10977 2941 11011 2975
rect 11621 2941 11655 2975
rect 12817 2941 12851 2975
rect 13829 2941 13863 2975
rect 14473 2941 14507 2975
rect 15209 2941 15243 2975
rect 16497 2941 16531 2975
rect 17233 2941 17267 2975
rect 18061 2941 18095 2975
rect 4169 2873 4203 2907
rect 5089 2873 5123 2907
rect 6101 2873 6135 2907
rect 6561 2873 6595 2907
rect 7113 2873 7147 2907
rect 7481 2873 7515 2907
rect 8953 2873 8987 2907
rect 9965 2873 9999 2907
rect 11897 2873 11931 2907
rect 13921 2873 13955 2907
rect 15485 2873 15519 2907
rect 16773 2873 16807 2907
rect 2053 2805 2087 2839
rect 2145 2805 2179 2839
rect 2697 2805 2731 2839
rect 3065 2805 3099 2839
rect 3617 2805 3651 2839
rect 3709 2805 3743 2839
rect 4721 2805 4755 2839
rect 5733 2805 5767 2839
rect 6193 2805 6227 2839
rect 10057 2805 10091 2839
rect 10609 2805 10643 2839
rect 12909 2805 12943 2839
rect 1685 2601 1719 2635
rect 2697 2601 2731 2635
rect 3065 2601 3099 2635
rect 4261 2601 4295 2635
rect 4629 2601 4663 2635
rect 5273 2601 5307 2635
rect 5641 2601 5675 2635
rect 9137 2601 9171 2635
rect 10057 2601 10091 2635
rect 10425 2601 10459 2635
rect 16589 2601 16623 2635
rect 2145 2533 2179 2567
rect 2053 2465 2087 2499
rect 4721 2465 4755 2499
rect 5733 2465 5767 2499
rect 6285 2465 6319 2499
rect 7113 2465 7147 2499
rect 7941 2465 7975 2499
rect 9045 2465 9079 2499
rect 10517 2465 10551 2499
rect 11069 2465 11103 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 16773 2465 16807 2499
rect 17509 2465 17543 2499
rect 2329 2397 2363 2431
rect 3157 2397 3191 2431
rect 3249 2397 3283 2431
rect 4905 2397 4939 2431
rect 5825 2397 5859 2431
rect 7389 2397 7423 2431
rect 8217 2397 8251 2431
rect 9321 2397 9355 2431
rect 10701 2397 10735 2431
rect 11253 2397 11287 2431
rect 11989 2397 12023 2431
rect 12817 2397 12851 2431
rect 17049 2397 17083 2431
rect 17785 2397 17819 2431
rect 6469 2329 6503 2363
rect 8677 2329 8711 2363
<< metal1 >>
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 2501 14603 2559 14609
rect 2501 14569 2513 14603
rect 2547 14600 2559 14603
rect 2774 14600 2780 14612
rect 2547 14572 2780 14600
rect 2547 14569 2559 14572
rect 2501 14563 2559 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5040 14572 5457 14600
rect 5040 14560 5046 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1627 14436 1992 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 1964 14396 1992 14436
rect 2038 14424 2044 14476
rect 2096 14464 2102 14476
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 2096 14436 2329 14464
rect 2096 14424 2102 14436
rect 2317 14433 2329 14436
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 5166 14424 5172 14476
rect 5224 14464 5230 14476
rect 5261 14467 5319 14473
rect 5261 14464 5273 14467
rect 5224 14436 5273 14464
rect 5224 14424 5230 14436
rect 5261 14433 5273 14436
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 3050 14396 3056 14408
rect 1964 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 17678 14396 17684 14408
rect 4120 14368 17684 14396
rect 4120 14356 4126 14368
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 1670 14288 1676 14340
rect 1728 14328 1734 14340
rect 14642 14328 14648 14340
rect 1728 14300 14648 14328
rect 1728 14288 1734 14300
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 5166 14260 5172 14272
rect 5127 14232 5172 14260
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 3234 14056 3240 14068
rect 3195 14028 3240 14056
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 3476 14028 4077 14056
rect 3476 14016 3482 14028
rect 4065 14025 4077 14028
rect 4111 14025 4123 14059
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 4065 14019 4123 14025
rect 5920 14028 7941 14056
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2774 13920 2780 13932
rect 2639 13892 2780 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 5920 13920 5948 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 16206 14056 16212 14068
rect 11848 14028 16212 14056
rect 11848 14016 11854 14028
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 17589 14059 17647 14065
rect 17589 14056 17601 14059
rect 16316 14028 17601 14056
rect 16316 13988 16344 14028
rect 17589 14025 17601 14028
rect 17635 14025 17647 14059
rect 17589 14019 17647 14025
rect 17678 14016 17684 14068
rect 17736 14056 17742 14068
rect 18233 14059 18291 14065
rect 18233 14056 18245 14059
rect 17736 14028 18245 14056
rect 17736 14016 17742 14028
rect 18233 14025 18245 14028
rect 18279 14025 18291 14059
rect 18233 14019 18291 14025
rect 6196 13960 16344 13988
rect 6196 13920 6224 13960
rect 16850 13948 16856 14000
rect 16908 13988 16914 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16908 13960 17049 13988
rect 16908 13948 16914 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 6362 13920 6368 13932
rect 3896 13892 5948 13920
rect 6104 13892 6224 13920
rect 6323 13892 6368 13920
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13821 1639 13855
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1581 13815 1639 13821
rect 1596 13716 1624 13815
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 2317 13815 2375 13821
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 2332 13784 2360 13815
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3896 13861 3924 13892
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13821 3939 13855
rect 3881 13815 3939 13821
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 6104 13852 6132 13892
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 7558 13920 7564 13932
rect 7519 13892 7564 13920
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 8294 13920 8300 13932
rect 8255 13892 8300 13920
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14918 13920 14924 13932
rect 14415 13892 14924 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 4028 13824 6132 13852
rect 6181 13855 6239 13861
rect 4028 13812 4034 13824
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 7282 13852 7288 13864
rect 6227 13824 7288 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7742 13812 7748 13864
rect 7800 13852 7806 13864
rect 7929 13855 7987 13861
rect 7929 13852 7941 13855
rect 7800 13824 7941 13852
rect 7800 13812 7806 13824
rect 7929 13821 7941 13824
rect 7975 13852 7987 13855
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 7975 13824 8033 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 14103 13855 14161 13861
rect 14103 13821 14115 13855
rect 14149 13821 14161 13855
rect 14103 13815 14161 13821
rect 1728 13756 2360 13784
rect 6089 13787 6147 13793
rect 1728 13744 1734 13756
rect 6089 13753 6101 13787
rect 6135 13784 6147 13787
rect 6135 13756 7052 13784
rect 6135 13753 6147 13756
rect 6089 13747 6147 13753
rect 2222 13716 2228 13728
rect 1596 13688 2228 13716
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 7024 13725 7052 13756
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 12342 13784 12348 13796
rect 11664 13756 12348 13784
rect 11664 13744 11670 13756
rect 12342 13744 12348 13756
rect 12400 13784 12406 13796
rect 14108 13784 14136 13815
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 14700 13824 16865 13852
rect 14700 13812 14706 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 17218 13812 17224 13864
rect 17276 13852 17282 13864
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17276 13824 17417 13852
rect 17276 13812 17282 13824
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13852 18107 13855
rect 18230 13852 18236 13864
rect 18095 13824 18236 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 12400 13756 14136 13784
rect 12400 13744 12406 13756
rect 7009 13719 7067 13725
rect 7009 13685 7021 13719
rect 7055 13685 7067 13719
rect 7374 13716 7380 13728
rect 7335 13688 7380 13716
rect 7009 13679 7067 13685
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 7524 13688 7569 13716
rect 7524 13676 7530 13688
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13512 2559 13515
rect 2866 13512 2872 13524
rect 2547 13484 2872 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5718 13512 5724 13524
rect 5307 13484 5724 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6917 13515 6975 13521
rect 6917 13481 6929 13515
rect 6963 13512 6975 13515
rect 7282 13512 7288 13524
rect 6963 13484 7288 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 14642 13512 14648 13524
rect 7423 13484 14648 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 1854 13444 1860 13456
rect 1815 13416 1860 13444
rect 1854 13404 1860 13416
rect 1912 13404 1918 13456
rect 8202 13444 8208 13456
rect 5552 13416 8208 13444
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13376 1642 13388
rect 2038 13376 2044 13388
rect 1636 13348 2044 13376
rect 1636 13336 1642 13348
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2317 13379 2375 13385
rect 2317 13376 2329 13379
rect 2280 13348 2329 13376
rect 2280 13336 2286 13348
rect 2317 13345 2329 13348
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 5552 13317 5580 13416
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 6822 13376 6828 13388
rect 6319 13348 6828 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 7248 13348 7297 13376
rect 7248 13336 7254 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 8757 13379 8815 13385
rect 8757 13376 8769 13379
rect 7285 13339 7343 13345
rect 7392 13348 8769 13376
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 5368 13240 5396 13271
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 5776 13280 6377 13308
rect 5776 13268 5782 13280
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 5905 13243 5963 13249
rect 5905 13240 5917 13243
rect 5368 13212 5917 13240
rect 5905 13209 5917 13212
rect 5951 13209 5963 13243
rect 5905 13203 5963 13209
rect 6270 13200 6276 13252
rect 6328 13240 6334 13252
rect 6472 13240 6500 13271
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 7392 13308 7420 13348
rect 8757 13345 8769 13348
rect 8803 13376 8815 13379
rect 9030 13376 9036 13388
rect 8803 13348 9036 13376
rect 8803 13345 8815 13348
rect 8757 13339 8815 13345
rect 9030 13336 9036 13348
rect 9088 13336 9094 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 9824 13348 10885 13376
rect 9824 13336 9830 13348
rect 10873 13345 10885 13348
rect 10919 13376 10931 13379
rect 16206 13376 16212 13388
rect 10919 13348 16212 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 7558 13308 7564 13320
rect 6696 13280 7420 13308
rect 7519 13280 7564 13308
rect 6696 13268 6702 13280
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 8846 13308 8852 13320
rect 8807 13280 8852 13308
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 10962 13308 10968 13320
rect 10923 13280 10968 13308
rect 8941 13271 8999 13277
rect 6328 13212 6500 13240
rect 8389 13243 8447 13249
rect 6328 13200 6334 13212
rect 8389 13209 8401 13243
rect 8435 13240 8447 13243
rect 8570 13240 8576 13252
rect 8435 13212 8576 13240
rect 8435 13209 8447 13212
rect 8389 13203 8447 13209
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 8956 13240 8984 13271
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11072 13240 11100 13271
rect 8812 13212 8984 13240
rect 10980 13212 11100 13240
rect 8812 13200 8818 13212
rect 10980 13184 11008 13212
rect 4893 13175 4951 13181
rect 4893 13141 4905 13175
rect 4939 13172 4951 13175
rect 6086 13172 6092 13184
rect 4939 13144 6092 13172
rect 4939 13141 4951 13144
rect 4893 13135 4951 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 8478 13132 8484 13184
rect 8536 13172 8542 13184
rect 10505 13175 10563 13181
rect 10505 13172 10517 13175
rect 8536 13144 10517 13172
rect 8536 13132 8542 13144
rect 10505 13141 10517 13144
rect 10551 13141 10563 13175
rect 10505 13135 10563 13141
rect 10962 13132 10968 13184
rect 11020 13132 11026 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 2958 12968 2964 12980
rect 1903 12940 2964 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 6822 12968 6828 12980
rect 6783 12940 6828 12968
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 10778 12968 10784 12980
rect 7208 12940 10784 12968
rect 7208 12912 7236 12940
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 3237 12903 3295 12909
rect 3237 12869 3249 12903
rect 3283 12900 3295 12903
rect 4522 12900 4528 12912
rect 3283 12872 4528 12900
rect 3283 12869 3295 12872
rect 3237 12863 3295 12869
rect 4522 12860 4528 12872
rect 4580 12860 4586 12912
rect 7190 12900 7196 12912
rect 4724 12872 7196 12900
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2740 12804 2789 12832
rect 2740 12792 2746 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 1762 12724 1768 12776
rect 1820 12764 1826 12776
rect 3804 12764 3832 12795
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4724 12832 4752 12872
rect 7190 12860 7196 12872
rect 7248 12860 7254 12912
rect 13814 12900 13820 12912
rect 10336 12872 13820 12900
rect 10336 12844 10364 12872
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 15562 12860 15568 12912
rect 15620 12900 15626 12912
rect 15746 12900 15752 12912
rect 15620 12872 15752 12900
rect 15620 12860 15626 12872
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 4890 12832 4896 12844
rect 4120 12804 4752 12832
rect 4851 12804 4896 12832
rect 4120 12792 4126 12804
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 7282 12832 7288 12844
rect 6411 12804 7288 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 7282 12792 7288 12804
rect 7340 12832 7346 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7340 12804 7481 12832
rect 7340 12792 7346 12804
rect 7469 12801 7481 12804
rect 7515 12832 7527 12835
rect 7558 12832 7564 12844
rect 7515 12804 7564 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12832 8631 12835
rect 9122 12832 9128 12844
rect 8619 12804 9128 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 10318 12832 10324 12844
rect 10231 12804 10324 12832
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 10502 12832 10508 12844
rect 10463 12804 10508 12832
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 12066 12832 12072 12844
rect 11563 12804 12072 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12584 12804 12817 12832
rect 12584 12792 12590 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 1820 12736 3832 12764
rect 4801 12767 4859 12773
rect 1820 12724 1826 12736
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5718 12764 5724 12776
rect 4847 12736 5724 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 8846 12764 8852 12776
rect 6012 12736 8852 12764
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 6012 12696 6040 12736
rect 8846 12724 8852 12736
rect 8904 12764 8910 12776
rect 10226 12764 10232 12776
rect 8904 12736 10232 12764
rect 8904 12724 8910 12736
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12400 12736 12449 12764
rect 12400 12724 12406 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 15562 12764 15568 12776
rect 15344 12736 15568 12764
rect 15344 12724 15350 12736
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 3292 12668 6040 12696
rect 6089 12699 6147 12705
rect 3292 12656 3298 12668
rect 6089 12665 6101 12699
rect 6135 12696 6147 12699
rect 6730 12696 6736 12708
rect 6135 12668 6736 12696
rect 6135 12665 6147 12668
rect 6089 12659 6147 12665
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 7193 12699 7251 12705
rect 7193 12665 7205 12699
rect 7239 12696 7251 12699
rect 7558 12696 7564 12708
rect 7239 12668 7564 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 10134 12696 10140 12708
rect 9088 12668 10140 12696
rect 9088 12656 9094 12668
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 10410 12656 10416 12708
rect 10468 12696 10474 12708
rect 11333 12699 11391 12705
rect 11333 12696 11345 12699
rect 10468 12668 11345 12696
rect 10468 12656 10474 12668
rect 11333 12665 11345 12668
rect 11379 12665 11391 12699
rect 11333 12659 11391 12665
rect 2225 12631 2283 12637
rect 2225 12597 2237 12631
rect 2271 12628 2283 12631
rect 2314 12628 2320 12640
rect 2271 12600 2320 12628
rect 2271 12597 2283 12600
rect 2225 12591 2283 12597
rect 2314 12588 2320 12600
rect 2372 12588 2378 12640
rect 2590 12628 2596 12640
rect 2551 12600 2596 12628
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 2685 12631 2743 12637
rect 2685 12597 2697 12631
rect 2731 12628 2743 12631
rect 3050 12628 3056 12640
rect 2731 12600 3056 12628
rect 2731 12597 2743 12600
rect 2685 12591 2743 12597
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 3602 12628 3608 12640
rect 3563 12600 3608 12628
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 3694 12588 3700 12640
rect 3752 12628 3758 12640
rect 4341 12631 4399 12637
rect 3752 12600 3797 12628
rect 3752 12588 3758 12600
rect 4341 12597 4353 12631
rect 4387 12628 4399 12631
rect 4430 12628 4436 12640
rect 4387 12600 4436 12628
rect 4387 12597 4399 12600
rect 4341 12591 4399 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 4706 12628 4712 12640
rect 4667 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 6178 12588 6184 12640
rect 6236 12628 6242 12640
rect 6236 12600 6281 12628
rect 6236 12588 6242 12600
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 7285 12631 7343 12637
rect 7285 12628 7297 12631
rect 6420 12600 7297 12628
rect 6420 12588 6426 12600
rect 7285 12597 7297 12600
rect 7331 12597 7343 12631
rect 7926 12628 7932 12640
rect 7887 12600 7932 12628
rect 7285 12591 7343 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8294 12628 8300 12640
rect 8255 12600 8300 12628
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12628 8447 12631
rect 8846 12628 8852 12640
rect 8435 12600 8852 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9824 12600 9873 12628
rect 9824 12588 9830 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10229 12631 10287 12637
rect 10229 12628 10241 12631
rect 10008 12600 10241 12628
rect 10008 12588 10014 12600
rect 10229 12597 10241 12600
rect 10275 12597 10287 12631
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10229 12591 10287 12597
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11241 12631 11299 12637
rect 11241 12628 11253 12631
rect 11112 12600 11253 12628
rect 11112 12588 11118 12600
rect 11241 12597 11253 12600
rect 11287 12597 11299 12631
rect 11241 12591 11299 12597
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 17586 12628 17592 12640
rect 14700 12600 17592 12628
rect 14700 12588 14706 12600
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 1765 12427 1823 12433
rect 1765 12393 1777 12427
rect 1811 12424 1823 12427
rect 2590 12424 2596 12436
rect 1811 12396 2596 12424
rect 1811 12393 1823 12396
rect 1765 12387 1823 12393
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 2700 12396 4077 12424
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2700 12356 2728 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 4522 12424 4528 12436
rect 4483 12396 4528 12424
rect 4065 12387 4123 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5077 12427 5135 12433
rect 5077 12424 5089 12427
rect 4764 12396 5089 12424
rect 4764 12384 4770 12396
rect 5077 12393 5089 12396
rect 5123 12393 5135 12427
rect 5077 12387 5135 12393
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5316 12396 5457 12424
rect 5316 12384 5322 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 5445 12387 5503 12393
rect 6089 12427 6147 12433
rect 6089 12393 6101 12427
rect 6135 12424 6147 12427
rect 6178 12424 6184 12436
rect 6135 12396 6184 12424
rect 6135 12393 6147 12396
rect 6089 12387 6147 12393
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6454 12424 6460 12436
rect 6415 12396 6460 12424
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7432 12396 7481 12424
rect 7432 12384 7438 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 10318 12424 10324 12436
rect 7469 12387 7527 12393
rect 7944 12396 10324 12424
rect 2556 12328 2728 12356
rect 3145 12359 3203 12365
rect 2556 12316 2562 12328
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 6638 12356 6644 12368
rect 3191 12328 6644 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 2130 12288 2136 12300
rect 2091 12260 2136 12288
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 3234 12288 3240 12300
rect 3195 12260 3240 12288
rect 3234 12248 3240 12260
rect 3292 12248 3298 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 5350 12288 5356 12300
rect 4479 12260 5356 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 6546 12288 6552 12300
rect 6459 12260 6552 12288
rect 6546 12248 6552 12260
rect 6604 12288 6610 12300
rect 6604 12260 6868 12288
rect 6604 12248 6610 12260
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 2096 12192 2237 12220
rect 2096 12180 2102 12192
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2225 12183 2283 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 4614 12220 4620 12232
rect 4575 12192 4620 12220
rect 3329 12183 3387 12189
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 3344 12152 3372 12183
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 4856 12192 5549 12220
rect 4856 12180 4862 12192
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12220 5779 12223
rect 6178 12220 6184 12232
rect 5767 12192 6184 12220
rect 5767 12189 5779 12192
rect 5721 12183 5779 12189
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 6638 12220 6644 12232
rect 6599 12192 6644 12220
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6840 12220 6868 12260
rect 7944 12220 7972 12396
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 10827 12396 11345 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 11333 12393 11345 12396
rect 11379 12393 11391 12427
rect 16114 12424 16120 12436
rect 11333 12387 11391 12393
rect 11716 12396 15976 12424
rect 16075 12396 16120 12424
rect 8389 12359 8447 12365
rect 8389 12356 8401 12359
rect 6840 12192 7972 12220
rect 8312 12328 8401 12356
rect 8312 12220 8340 12328
rect 8389 12325 8401 12328
rect 8435 12325 8447 12359
rect 8389 12319 8447 12325
rect 8481 12359 8539 12365
rect 8481 12325 8493 12359
rect 8527 12356 8539 12359
rect 8570 12356 8576 12368
rect 8527 12328 8576 12356
rect 8527 12325 8539 12328
rect 8481 12319 8539 12325
rect 8570 12316 8576 12328
rect 8628 12316 8634 12368
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 11606 12356 11612 12368
rect 8996 12328 11612 12356
rect 8996 12316 9002 12328
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 9950 12288 9956 12300
rect 9088 12260 9956 12288
rect 9088 12248 9094 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10686 12288 10692 12300
rect 10647 12260 10692 12288
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 10778 12248 10784 12300
rect 10836 12288 10842 12300
rect 11716 12297 11744 12396
rect 15948 12356 15976 12396
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 17586 12424 17592 12436
rect 17547 12396 17592 12424
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 17497 12359 17555 12365
rect 17497 12356 17509 12359
rect 15212 12328 15875 12356
rect 15948 12328 17509 12356
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 10836 12260 11713 12288
rect 10836 12248 10842 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 15212 12288 15240 12328
rect 11701 12251 11759 12257
rect 12268 12260 15240 12288
rect 8386 12220 8392 12232
rect 8312 12192 8392 12220
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 9122 12220 9128 12232
rect 8711 12192 9128 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 9272 12192 10977 12220
rect 9272 12180 9278 12192
rect 10965 12189 10977 12192
rect 11011 12220 11023 12223
rect 11514 12220 11520 12232
rect 11011 12192 11520 12220
rect 11011 12189 11023 12192
rect 10965 12183 11023 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11790 12220 11796 12232
rect 11664 12192 11796 12220
rect 11664 12180 11670 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 11940 12192 11985 12220
rect 11940 12180 11946 12192
rect 12268 12152 12296 12260
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15746 12288 15752 12300
rect 15344 12260 15752 12288
rect 15344 12248 15350 12260
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 15847 12288 15875 12328
rect 17497 12325 17509 12328
rect 17543 12356 17555 12359
rect 17862 12356 17868 12368
rect 17543 12328 17868 12356
rect 17543 12325 17555 12328
rect 17497 12319 17555 12325
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 17954 12288 17960 12300
rect 15847 12260 17960 12288
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 14182 12180 14188 12232
rect 14240 12220 14246 12232
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 14240 12192 16221 12220
rect 14240 12180 14246 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12220 16359 12223
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 16347 12192 17693 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 18138 12220 18144 12232
rect 18099 12192 18144 12220
rect 17681 12183 17739 12189
rect 3200 12124 3372 12152
rect 10152 12124 12296 12152
rect 3200 12112 3206 12124
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 3326 12084 3332 12096
rect 2823 12056 3332 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 3694 12044 3700 12096
rect 3752 12084 3758 12096
rect 7834 12084 7840 12096
rect 3752 12056 7840 12084
rect 3752 12044 3758 12056
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 10152 12084 10180 12124
rect 15010 12112 15016 12164
rect 15068 12152 15074 12164
rect 16316 12152 16344 12183
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 15068 12124 16344 12152
rect 15068 12112 15074 12124
rect 10318 12084 10324 12096
rect 8628 12056 10180 12084
rect 10279 12056 10324 12084
rect 8628 12044 8634 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 12342 12044 12348 12096
rect 12400 12084 12406 12096
rect 15194 12084 15200 12096
rect 12400 12056 15200 12084
rect 12400 12044 12406 12056
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 16482 12084 16488 12096
rect 15795 12056 16488 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 17129 12087 17187 12093
rect 17129 12084 17141 12087
rect 17092 12056 17141 12084
rect 17092 12044 17098 12056
rect 17129 12053 17141 12056
rect 17175 12053 17187 12087
rect 17129 12047 17187 12053
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 6328 11852 6469 11880
rect 6328 11840 6334 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 3602 11772 3608 11824
rect 3660 11812 3666 11824
rect 3660 11784 4476 11812
rect 3660 11772 3666 11784
rect 3418 11744 3424 11756
rect 3160 11716 3424 11744
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11645 2099 11679
rect 2041 11639 2099 11645
rect 2308 11679 2366 11685
rect 2308 11645 2320 11679
rect 2354 11676 2366 11679
rect 2590 11676 2596 11688
rect 2354 11648 2596 11676
rect 2354 11645 2366 11648
rect 2308 11639 2366 11645
rect 2056 11540 2084 11639
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 2406 11568 2412 11620
rect 2464 11608 2470 11620
rect 3160 11608 3188 11716
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 4338 11744 4344 11756
rect 4299 11716 4344 11744
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 4448 11744 4476 11784
rect 6472 11744 6500 11843
rect 6822 11840 6828 11892
rect 6880 11880 6886 11892
rect 10778 11880 10784 11892
rect 6880 11852 8524 11880
rect 6880 11840 6886 11852
rect 8496 11753 8524 11852
rect 9508 11852 10784 11880
rect 8481 11747 8539 11753
rect 4448 11716 5212 11744
rect 6472 11716 6960 11744
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 4246 11676 4252 11688
rect 4203 11648 4252 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 5077 11679 5135 11685
rect 5077 11645 5089 11679
rect 5123 11645 5135 11679
rect 5184 11676 5212 11716
rect 5184 11648 5304 11676
rect 5077 11639 5135 11645
rect 4062 11608 4068 11620
rect 2464 11580 3188 11608
rect 3252 11580 4068 11608
rect 2464 11568 2470 11580
rect 3252 11540 3280 11580
rect 4062 11568 4068 11580
rect 4120 11608 4126 11620
rect 5092 11608 5120 11639
rect 4120 11580 5120 11608
rect 4120 11568 4126 11580
rect 3418 11540 3424 11552
rect 2056 11512 3280 11540
rect 3379 11512 3424 11540
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 3789 11543 3847 11549
rect 3789 11540 3801 11543
rect 3568 11512 3801 11540
rect 3568 11500 3574 11512
rect 3789 11509 3801 11512
rect 3835 11509 3847 11543
rect 3789 11503 3847 11509
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 5166 11540 5172 11552
rect 4295 11512 5172 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5276 11540 5304 11648
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 6362 11676 6368 11688
rect 5684 11648 6368 11676
rect 5684 11636 5690 11648
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 6822 11676 6828 11688
rect 6783 11648 6828 11676
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 6932 11676 6960 11716
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6932 11648 7093 11676
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 9508 11676 9536 11852
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11238 11840 11244 11892
rect 11296 11840 11302 11892
rect 11514 11880 11520 11892
rect 11475 11852 11520 11880
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 13311 11852 13369 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13357 11849 13369 11852
rect 13403 11849 13415 11883
rect 13357 11843 13415 11849
rect 11256 11812 11284 11840
rect 14366 11812 14372 11824
rect 11256 11784 14372 11812
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 12066 11744 12072 11756
rect 7081 11639 7139 11645
rect 7392 11648 9536 11676
rect 9600 11716 10272 11744
rect 5344 11611 5402 11617
rect 5344 11577 5356 11611
rect 5390 11608 5402 11611
rect 7282 11608 7288 11620
rect 5390 11580 7288 11608
rect 5390 11577 5402 11580
rect 5344 11571 5402 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 7392 11540 7420 11648
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 8748 11611 8806 11617
rect 8168 11580 8708 11608
rect 8168 11568 8174 11580
rect 8202 11540 8208 11552
rect 5276 11512 7420 11540
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8680 11540 8708 11580
rect 8748 11577 8760 11611
rect 8794 11608 8806 11611
rect 9214 11608 9220 11620
rect 8794 11580 9220 11608
rect 8794 11577 8806 11580
rect 8748 11571 8806 11577
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 9600 11540 9628 11716
rect 10134 11676 10140 11688
rect 10095 11648 10140 11676
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 10244 11676 10272 11716
rect 11164 11716 12072 11744
rect 11164 11676 11192 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13688 11716 13921 11744
rect 13688 11704 13694 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 16482 11744 16488 11756
rect 16443 11716 16488 11744
rect 13909 11707 13967 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11744 16727 11747
rect 17126 11744 17132 11756
rect 16715 11716 17132 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 10244 11648 11192 11676
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 12158 11676 12164 11688
rect 11296 11648 12164 11676
rect 11296 11636 11302 11648
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13998 11676 14004 11688
rect 13771 11648 14004 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14090 11636 14096 11688
rect 14148 11676 14154 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14148 11648 14381 11676
rect 14148 11636 14154 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 16574 11676 16580 11688
rect 14369 11639 14427 11645
rect 14476 11648 16580 11676
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10382 11611 10440 11617
rect 10382 11608 10394 11611
rect 9732 11580 10394 11608
rect 9732 11568 9738 11580
rect 10382 11577 10394 11580
rect 10428 11608 10440 11611
rect 11514 11608 11520 11620
rect 10428 11580 11520 11608
rect 10428 11577 10440 11580
rect 10382 11571 10440 11577
rect 11514 11568 11520 11580
rect 11572 11608 11578 11620
rect 11882 11608 11888 11620
rect 11572 11580 11888 11608
rect 11572 11568 11578 11580
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 13265 11611 13323 11617
rect 13265 11577 13277 11611
rect 13311 11608 13323 11611
rect 13906 11608 13912 11620
rect 13311 11580 13912 11608
rect 13311 11577 13323 11580
rect 13265 11571 13323 11577
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 14016 11608 14044 11636
rect 14476 11608 14504 11648
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16816 11648 17417 11676
rect 16816 11636 16822 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17770 11636 17776 11688
rect 17828 11676 17834 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17828 11648 18061 11676
rect 17828 11636 17834 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 14016 11580 14504 11608
rect 14636 11611 14694 11617
rect 14636 11577 14648 11611
rect 14682 11608 14694 11611
rect 14734 11608 14740 11620
rect 14682 11580 14740 11608
rect 14682 11577 14694 11580
rect 14636 11571 14694 11577
rect 14734 11568 14740 11580
rect 14792 11568 14798 11620
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 16393 11611 16451 11617
rect 16393 11608 16405 11611
rect 14884 11580 16405 11608
rect 14884 11568 14890 11580
rect 16393 11577 16405 11580
rect 16439 11577 16451 11611
rect 16393 11571 16451 11577
rect 8680 11512 9628 11540
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10134 11540 10140 11552
rect 9907 11512 10140 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11296 11512 11805 11540
rect 11296 11500 11302 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13504 11512 13829 11540
rect 13504 11500 13510 11512
rect 13817 11509 13829 11512
rect 13863 11540 13875 11543
rect 14274 11540 14280 11552
rect 13863 11512 14280 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15068 11512 15761 11540
rect 15068 11500 15074 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 15749 11503 15807 11509
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16114 11540 16120 11552
rect 16071 11512 16120 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 17589 11543 17647 11549
rect 17589 11540 17601 11543
rect 16540 11512 17601 11540
rect 16540 11500 16546 11512
rect 17589 11509 17601 11512
rect 17635 11509 17647 11543
rect 17589 11503 17647 11509
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 18322 11540 18328 11552
rect 18279 11512 18328 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2774 11336 2780 11348
rect 2455 11308 2780 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 1946 11268 1952 11280
rect 1859 11240 1952 11268
rect 1946 11228 1952 11240
rect 2004 11268 2010 11280
rect 2424 11268 2452 11299
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4396 11308 5457 11336
rect 4396 11296 4402 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5718 11336 5724 11348
rect 5679 11308 5724 11336
rect 5445 11299 5503 11305
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 5868 11308 6193 11336
rect 5868 11296 5874 11308
rect 6181 11305 6193 11308
rect 6227 11305 6239 11339
rect 6181 11299 6239 11305
rect 8021 11339 8079 11345
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8478 11336 8484 11348
rect 8067 11308 8484 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8938 11336 8944 11348
rect 8899 11308 8944 11336
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11336 10103 11339
rect 10318 11336 10324 11348
rect 10091 11308 10324 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10744 11308 10885 11336
rect 10744 11296 10750 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 10873 11299 10931 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 17681 11339 17739 11345
rect 11379 11308 14596 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 2004 11240 2452 11268
rect 2004 11228 2010 11240
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 9858 11268 9864 11280
rect 6420 11240 9864 11268
rect 6420 11228 6426 11240
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 11348 11268 11376 11299
rect 14090 11268 14096 11280
rect 10397 11240 11376 11268
rect 13096 11240 14096 11268
rect 2501 11203 2559 11209
rect 2501 11200 2513 11203
rect 1964 11172 2513 11200
rect 1964 11144 1992 11172
rect 2501 11169 2513 11172
rect 2547 11169 2559 11203
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 2501 11163 2559 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4706 11200 4712 11212
rect 4378 11172 4712 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5258 11160 5264 11212
rect 5316 11160 5322 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 1946 11092 1952 11144
rect 2004 11092 2010 11144
rect 2590 11132 2596 11144
rect 2551 11104 2596 11132
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3053 11135 3111 11141
rect 3053 11132 3065 11135
rect 2924 11104 3065 11132
rect 2924 11092 2930 11104
rect 3053 11101 3065 11104
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 4080 11132 4108 11160
rect 3660 11104 4108 11132
rect 5276 11132 5304 11160
rect 6104 11132 6132 11163
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7708 11172 7941 11200
rect 7708 11160 7714 11172
rect 7929 11169 7941 11172
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 5276 11104 6132 11132
rect 3660 11092 3666 11104
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 6236 11104 6285 11132
rect 6236 11092 6242 11104
rect 6273 11101 6285 11104
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 5316 11036 7573 11064
rect 5316 11024 5322 11036
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 7561 11027 7619 11033
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 7834 10996 7840 11008
rect 3844 10968 7840 10996
rect 3844 10956 3850 10968
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 7944 10996 7972 11163
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 10397 11200 10425 11240
rect 12250 11200 12256 11212
rect 8536 11172 10425 11200
rect 12211 11172 12256 11200
rect 8536 11160 8542 11172
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 13096 11209 13124 11240
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14568 11268 14596 11308
rect 17681 11305 17693 11339
rect 17727 11336 17739 11339
rect 18138 11336 18144 11348
rect 17727 11308 18144 11336
rect 17727 11305 17739 11308
rect 17681 11299 17739 11305
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 17773 11271 17831 11277
rect 17773 11268 17785 11271
rect 14568 11240 17785 11268
rect 17773 11237 17785 11240
rect 17819 11268 17831 11271
rect 18046 11268 18052 11280
rect 17819 11240 18052 11268
rect 17819 11237 17831 11240
rect 17773 11231 17831 11237
rect 18046 11228 18052 11240
rect 18104 11228 18110 11280
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11169 13139 11203
rect 13081 11163 13139 11169
rect 13348 11203 13406 11209
rect 13348 11169 13360 11203
rect 13394 11200 13406 11203
rect 13722 11200 13728 11212
rect 13394 11172 13728 11200
rect 13394 11169 13406 11172
rect 13348 11163 13406 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15913 11203 15971 11209
rect 15913 11200 15925 11203
rect 15068 11172 15925 11200
rect 15068 11160 15074 11172
rect 15913 11169 15925 11172
rect 15959 11200 15971 11203
rect 15959 11172 17908 11200
rect 15959 11169 15971 11172
rect 15913 11163 15971 11169
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 8220 11064 8248 11095
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 8720 11104 9045 11132
rect 8720 11092 8726 11104
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 9033 11095 9091 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 8168 11036 8248 11064
rect 8573 11067 8631 11073
rect 8168 11024 8174 11036
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 10152 11064 10180 11095
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 11514 11132 11520 11144
rect 10284 11104 10329 11132
rect 11475 11104 11520 11132
rect 10284 11092 10290 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12526 11132 12532 11144
rect 12487 11104 12532 11132
rect 12345 11095 12403 11101
rect 8619 11036 10180 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 11974 11024 11980 11076
rect 12032 11024 12038 11076
rect 12360 11064 12388 11095
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 15102 11132 15108 11144
rect 14148 11104 15108 11132
rect 14148 11092 14154 11104
rect 15102 11092 15108 11104
rect 15160 11132 15166 11144
rect 17880 11141 17908 11172
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 15160 11104 15669 11132
rect 15160 11092 15166 11104
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 12710 11064 12716 11076
rect 12360 11036 12716 11064
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 11698 10996 11704 11008
rect 7944 10968 11704 10996
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 11885 10999 11943 11005
rect 11885 10965 11897 10999
rect 11931 10996 11943 10999
rect 11992 10996 12020 11024
rect 11931 10968 12020 10996
rect 14461 10999 14519 11005
rect 11931 10965 11943 10968
rect 11885 10959 11943 10965
rect 14461 10965 14473 10999
rect 14507 10996 14519 10999
rect 14734 10996 14740 11008
rect 14507 10968 14740 10996
rect 14507 10965 14519 10968
rect 14461 10959 14519 10965
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 17037 10999 17095 11005
rect 17037 10965 17049 10999
rect 17083 10996 17095 10999
rect 17126 10996 17132 11008
rect 17083 10968 17132 10996
rect 17083 10965 17095 10968
rect 17037 10959 17095 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17310 10996 17316 11008
rect 17271 10968 17316 10996
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2130 10792 2136 10804
rect 2087 10764 2136 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 5166 10752 5172 10804
rect 5224 10792 5230 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 5224 10764 5273 10792
rect 5224 10752 5230 10764
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 5626 10752 5632 10804
rect 5684 10752 5690 10804
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6546 10792 6552 10804
rect 5776 10764 6552 10792
rect 5776 10752 5782 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 6788 10764 7113 10792
rect 6788 10752 6794 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 8754 10792 8760 10804
rect 8715 10764 8760 10792
rect 7101 10755 7159 10761
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 8996 10764 9229 10792
rect 8996 10752 9002 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 10594 10792 10600 10804
rect 9217 10755 9275 10761
rect 10244 10764 10600 10792
rect 1673 10727 1731 10733
rect 1673 10693 1685 10727
rect 1719 10724 1731 10727
rect 2774 10724 2780 10736
rect 1719 10696 2780 10724
rect 1719 10693 1731 10696
rect 1673 10687 1731 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3418 10684 3424 10736
rect 3476 10724 3482 10736
rect 3476 10696 3648 10724
rect 3476 10684 3482 10696
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2648 10628 2697 10656
rect 2648 10616 2654 10628
rect 2685 10625 2697 10628
rect 2731 10656 2743 10659
rect 3510 10656 3516 10668
rect 2731 10628 3372 10656
rect 3471 10628 3516 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 1486 10588 1492 10600
rect 1447 10560 1492 10588
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 2866 10588 2872 10600
rect 2455 10560 2872 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3344 10588 3372 10628
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3620 10665 3648 10696
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4764 10628 4813 10656
rect 4764 10616 4770 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 4338 10588 4344 10600
rect 3344 10560 4344 10588
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 5644 10588 5672 10752
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6086 10656 6092 10668
rect 5951 10628 6092 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6086 10616 6092 10628
rect 6144 10616 6150 10668
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6788 10628 7420 10656
rect 6788 10616 6794 10628
rect 4663 10560 5672 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 7392 10597 7420 10628
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9582 10656 9588 10668
rect 9364 10628 9588 10656
rect 9364 10616 9370 10628
rect 9582 10616 9588 10628
rect 9640 10656 9646 10668
rect 10244 10665 10272 10764
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11572 10764 11621 10792
rect 11572 10752 11578 10764
rect 11609 10761 11621 10764
rect 11655 10761 11667 10795
rect 11609 10755 11667 10761
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12618 10792 12624 10804
rect 11756 10764 12624 10792
rect 11756 10752 11762 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 14090 10792 14096 10804
rect 14051 10764 14096 10792
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 14826 10792 14832 10804
rect 14415 10764 14832 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 18046 10724 18052 10736
rect 13464 10696 18052 10724
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9640 10628 9781 10656
rect 9640 10616 9646 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 7285 10591 7343 10597
rect 5776 10560 5821 10588
rect 5776 10548 5782 10560
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 7644 10591 7702 10597
rect 7644 10557 7656 10591
rect 7690 10588 7702 10591
rect 8202 10588 8208 10600
rect 7690 10560 8208 10588
rect 7690 10557 7702 10560
rect 7644 10551 7702 10557
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 2547 10492 6224 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 4028 10424 4721 10452
rect 4028 10412 4034 10424
rect 4709 10421 4721 10424
rect 4755 10452 4767 10455
rect 5166 10452 5172 10464
rect 4755 10424 5172 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 5994 10452 6000 10464
rect 5675 10424 6000 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6196 10452 6224 10492
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 7300 10520 7328 10551
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 10502 10597 10508 10600
rect 10496 10588 10508 10597
rect 10463 10560 10508 10588
rect 10496 10551 10508 10560
rect 10502 10548 10508 10551
rect 10560 10548 10566 10600
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11756 10560 12449 10588
rect 11756 10548 11762 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 13464 10588 13492 10696
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14090 10656 14096 10668
rect 13872 10628 14096 10656
rect 13872 10616 13878 10628
rect 14090 10616 14096 10628
rect 14148 10656 14154 10668
rect 14458 10656 14464 10668
rect 14148 10628 14464 10656
rect 14148 10616 14154 10628
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 15010 10656 15016 10668
rect 14971 10628 15016 10656
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16298 10656 16304 10668
rect 16071 10628 16304 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 17034 10656 17040 10668
rect 16995 10628 17040 10656
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17184 10628 17229 10656
rect 17184 10616 17190 10628
rect 12437 10551 12495 10557
rect 12544 10560 13492 10588
rect 6328 10492 7328 10520
rect 6328 10480 6334 10492
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 9585 10523 9643 10529
rect 9585 10520 9597 10523
rect 7892 10492 9597 10520
rect 7892 10480 7898 10492
rect 9585 10489 9597 10492
rect 9631 10520 9643 10523
rect 9631 10492 10364 10520
rect 9631 10489 9643 10492
rect 9585 10483 9643 10489
rect 7558 10452 7564 10464
rect 6196 10424 7564 10452
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9858 10452 9864 10464
rect 9723 10424 9864 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10336 10452 10364 10492
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 12544 10520 12572 10560
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14056 10560 14289 10588
rect 14056 10548 14062 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 14918 10588 14924 10600
rect 14875 10560 14924 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15562 10588 15568 10600
rect 15344 10560 15568 10588
rect 15344 10548 15350 10560
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10588 15899 10591
rect 16114 10588 16120 10600
rect 15887 10560 16120 10588
rect 15887 10557 15899 10560
rect 15841 10551 15899 10557
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 16945 10591 17003 10597
rect 16945 10557 16957 10591
rect 16991 10588 17003 10591
rect 17310 10588 17316 10600
rect 16991 10560 17316 10588
rect 16991 10557 17003 10560
rect 16945 10551 17003 10557
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17736 10560 18061 10588
rect 17736 10548 17742 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 12710 10529 12716 10532
rect 12704 10520 12716 10529
rect 10652 10492 12572 10520
rect 12671 10492 12716 10520
rect 10652 10480 10658 10492
rect 12704 10483 12716 10492
rect 12710 10480 12716 10483
rect 12768 10480 12774 10532
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 14737 10523 14795 10529
rect 14737 10520 14749 10523
rect 13320 10492 14749 10520
rect 13320 10480 13326 10492
rect 14737 10489 14749 10492
rect 14783 10489 14795 10523
rect 14737 10483 14795 10489
rect 15749 10523 15807 10529
rect 15749 10489 15761 10523
rect 15795 10520 15807 10523
rect 15795 10492 16620 10520
rect 15795 10489 15807 10492
rect 15749 10483 15807 10489
rect 11790 10452 11796 10464
rect 10336 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13780 10424 13829 10452
rect 13780 10412 13786 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15562 10452 15568 10464
rect 15427 10424 15568 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16114 10412 16120 10464
rect 16172 10452 16178 10464
rect 16390 10452 16396 10464
rect 16172 10424 16396 10452
rect 16172 10412 16178 10424
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16592 10461 16620 10492
rect 16577 10455 16635 10461
rect 16577 10421 16589 10455
rect 16623 10421 16635 10455
rect 18230 10452 18236 10464
rect 18191 10424 18236 10452
rect 16577 10415 16635 10421
rect 18230 10412 18236 10424
rect 18288 10412 18294 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 3602 10248 3608 10260
rect 3563 10220 3608 10248
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 7101 10251 7159 10257
rect 3752 10220 6776 10248
rect 3752 10208 3758 10220
rect 1664 10183 1722 10189
rect 1664 10149 1676 10183
rect 1710 10180 1722 10183
rect 2406 10180 2412 10192
rect 1710 10152 2412 10180
rect 1710 10149 1722 10152
rect 1664 10143 1722 10149
rect 2406 10140 2412 10152
rect 2464 10140 2470 10192
rect 5810 10180 5816 10192
rect 3804 10152 5816 10180
rect 3050 10112 3056 10124
rect 3011 10084 3056 10112
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 3804 10121 3832 10152
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 5988 10183 6046 10189
rect 5988 10149 6000 10183
rect 6034 10180 6046 10183
rect 6638 10180 6644 10192
rect 6034 10152 6644 10180
rect 6034 10149 6046 10152
rect 5988 10143 6046 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 6748 10180 6776 10220
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7282 10248 7288 10260
rect 7147 10220 7288 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 9030 10248 9036 10260
rect 8352 10220 9036 10248
rect 8352 10208 8358 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9858 10248 9864 10260
rect 9819 10220 9864 10248
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10744 10220 10885 10248
rect 10744 10208 10750 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 13265 10251 13323 10257
rect 13265 10248 13277 10251
rect 10873 10211 10931 10217
rect 11072 10220 13277 10248
rect 7466 10180 7472 10192
rect 6748 10152 7472 10180
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 8185 10183 8243 10189
rect 8185 10180 8197 10183
rect 7708 10152 8197 10180
rect 7708 10140 7714 10152
rect 8185 10149 8197 10152
rect 8231 10149 8243 10183
rect 8185 10143 8243 10149
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 10042 10180 10048 10192
rect 8536 10152 10048 10180
rect 8536 10140 8542 10152
rect 10042 10140 10048 10152
rect 10100 10140 10106 10192
rect 10229 10183 10287 10189
rect 10229 10149 10241 10183
rect 10275 10180 10287 10183
rect 10275 10152 10732 10180
rect 10275 10149 10287 10152
rect 10229 10143 10287 10149
rect 3789 10115 3847 10121
rect 3789 10081 3801 10115
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 5721 10115 5779 10121
rect 4479 10084 4936 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 3510 10044 3516 10056
rect 3292 10016 3516 10044
rect 3292 10004 3298 10016
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4525 10047 4583 10053
rect 3936 10016 4108 10044
rect 3936 10004 3942 10016
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 4080 9985 4108 10016
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4525 10007 4583 10013
rect 2777 9979 2835 9985
rect 2777 9976 2789 9979
rect 2740 9948 2789 9976
rect 2740 9936 2746 9948
rect 2777 9945 2789 9948
rect 2823 9945 2835 9979
rect 2777 9939 2835 9945
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9945 4123 9979
rect 4065 9939 4123 9945
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 4540 9908 4568 10007
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4908 9976 4936 10084
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6730 10112 6736 10124
rect 5767 10084 6736 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6730 10072 6736 10084
rect 6788 10112 6794 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 6788 10084 7941 10112
rect 6788 10072 6794 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 10244 10112 10272 10143
rect 10594 10112 10600 10124
rect 7929 10075 7987 10081
rect 8036 10084 10272 10112
rect 10336 10084 10600 10112
rect 5074 10044 5080 10056
rect 5035 10016 5080 10044
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 8036 10044 8064 10084
rect 10336 10053 10364 10084
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 7944 10016 8064 10044
rect 8956 10016 10333 10044
rect 5718 9976 5724 9988
rect 4908 9948 5724 9976
rect 5718 9936 5724 9948
rect 5776 9936 5782 9988
rect 6822 9936 6828 9988
rect 6880 9976 6886 9988
rect 7944 9976 7972 10016
rect 6880 9948 7972 9976
rect 6880 9936 6886 9948
rect 4706 9908 4712 9920
rect 4540 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9908 4770 9920
rect 8956 9908 8984 10016
rect 10321 10013 10333 10016
rect 10367 10013 10379 10047
rect 10502 10044 10508 10056
rect 10463 10016 10508 10044
rect 10321 10007 10379 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 10520 9976 10548 10004
rect 9355 9948 10548 9976
rect 10704 9976 10732 10152
rect 10888 10044 10916 10211
rect 11072 10121 11100 10220
rect 13265 10217 13277 10220
rect 13311 10248 13323 10251
rect 13998 10248 14004 10260
rect 13311 10220 14004 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14182 10248 14188 10260
rect 14143 10220 14188 10248
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14516 10220 14657 10248
rect 14516 10208 14522 10220
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 14645 10211 14703 10217
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 17310 10248 17316 10260
rect 15068 10220 17316 10248
rect 15068 10208 15074 10220
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18138 10248 18144 10260
rect 18099 10220 18144 10248
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 17405 10183 17463 10189
rect 17405 10180 17417 10183
rect 12860 10152 17417 10180
rect 12860 10140 12866 10152
rect 17405 10149 17417 10152
rect 17451 10149 17463 10183
rect 17405 10143 17463 10149
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10081 11115 10115
rect 11514 10112 11520 10124
rect 11475 10084 11520 10112
rect 11057 10075 11115 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11698 10112 11704 10124
rect 11624 10084 11704 10112
rect 11624 10053 11652 10084
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11876 10115 11934 10121
rect 11876 10081 11888 10115
rect 11922 10112 11934 10115
rect 13449 10115 13507 10121
rect 11922 10084 13216 10112
rect 11922 10081 11934 10084
rect 11876 10075 11934 10081
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 10888 10016 11621 10044
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 13188 10044 13216 10084
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 13495 10084 13553 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13541 10081 13553 10084
rect 13587 10081 13599 10115
rect 13541 10075 13599 10081
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 14553 10115 14611 10121
rect 14553 10112 14565 10115
rect 14424 10084 14565 10112
rect 14424 10072 14430 10084
rect 14553 10081 14565 10084
rect 14599 10112 14611 10115
rect 14826 10112 14832 10124
rect 14599 10084 14832 10112
rect 14599 10081 14611 10084
rect 14553 10075 14611 10081
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 15102 10072 15108 10124
rect 15160 10112 15166 10124
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 15160 10084 15301 10112
rect 15160 10072 15166 10084
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 15556 10115 15614 10121
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 17126 10112 17132 10124
rect 15602 10084 17132 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 17954 10112 17960 10124
rect 17644 10084 17960 10112
rect 17644 10072 17650 10084
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 13630 10044 13636 10056
rect 13188 10016 13636 10044
rect 11609 10007 11667 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14458 10044 14464 10056
rect 13771 10016 14464 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 14792 10016 14837 10044
rect 14792 10004 14798 10016
rect 16390 10004 16396 10056
rect 16448 10044 16454 10056
rect 16758 10044 16764 10056
rect 16448 10016 16764 10044
rect 16448 10004 16454 10016
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17494 10044 17500 10056
rect 17455 10016 17500 10044
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 11146 9976 11152 9988
rect 10704 9948 11152 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 13538 9976 13544 9988
rect 12636 9948 13544 9976
rect 4764 9880 8984 9908
rect 4764 9868 4770 9880
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 11238 9908 11244 9920
rect 9088 9880 11244 9908
rect 9088 9868 9094 9880
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11333 9911 11391 9917
rect 11333 9877 11345 9911
rect 11379 9908 11391 9911
rect 12636 9908 12664 9948
rect 13538 9936 13544 9948
rect 13596 9936 13602 9988
rect 11379 9880 12664 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12986 9908 12992 9920
rect 12768 9880 12992 9908
rect 12768 9868 12774 9880
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 13998 9908 14004 9920
rect 13320 9880 14004 9908
rect 13320 9868 13326 9880
rect 13998 9868 14004 9880
rect 14056 9868 14062 9920
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 16356 9880 16681 9908
rect 16356 9868 16362 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16669 9871 16727 9877
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3605 9707 3663 9713
rect 3605 9704 3617 9707
rect 3476 9676 3617 9704
rect 3476 9664 3482 9676
rect 3605 9673 3617 9676
rect 3651 9673 3663 9707
rect 3605 9667 3663 9673
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 6178 9704 6184 9716
rect 4488 9676 6184 9704
rect 4488 9664 4494 9676
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 10686 9704 10692 9716
rect 9692 9676 10692 9704
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6270 9636 6276 9648
rect 5868 9608 6276 9636
rect 5868 9596 5874 9608
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 8662 9636 8668 9648
rect 8623 9608 8668 9636
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3844 9540 4077 9568
rect 3844 9528 3850 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 4338 9568 4344 9580
rect 4295 9540 4344 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 6638 9568 6644 9580
rect 6012 9540 6644 9568
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1452 9472 1777 9500
rect 1452 9460 1458 9472
rect 1765 9469 1777 9472
rect 1811 9500 1823 9503
rect 2406 9500 2412 9512
rect 1811 9472 2412 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 3602 9500 3608 9512
rect 2464 9472 3608 9500
rect 2464 9460 2470 9472
rect 3602 9460 3608 9472
rect 3660 9500 3666 9512
rect 4890 9509 4896 9512
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 3660 9472 4629 9500
rect 3660 9460 3666 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 4884 9500 4896 9509
rect 4851 9472 4896 9500
rect 4617 9463 4675 9469
rect 4884 9463 4896 9472
rect 4890 9460 4896 9463
rect 4948 9460 4954 9512
rect 2032 9435 2090 9441
rect 2032 9401 2044 9435
rect 2078 9432 2090 9435
rect 2682 9432 2688 9444
rect 2078 9404 2688 9432
rect 2078 9401 2090 9404
rect 2032 9395 2090 9401
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 3050 9392 3056 9444
rect 3108 9432 3114 9444
rect 3970 9432 3976 9444
rect 3108 9404 3976 9432
rect 3108 9392 3114 9404
rect 3970 9392 3976 9404
rect 4028 9392 4034 9444
rect 3142 9364 3148 9376
rect 3055 9336 3148 9364
rect 3142 9324 3148 9336
rect 3200 9364 3206 9376
rect 3694 9364 3700 9376
rect 3200 9336 3700 9364
rect 3200 9324 3206 9336
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 6012 9373 6040 9540
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6788 9540 6837 9568
rect 6788 9528 6794 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 6825 9531 6883 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 9692 9577 9720 9676
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 12526 9704 12532 9716
rect 12308 9676 12532 9704
rect 12308 9664 12314 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 16666 9704 16672 9716
rect 13872 9676 16672 9704
rect 13872 9664 13878 9676
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 16945 9707 17003 9713
rect 16945 9704 16957 9707
rect 16816 9676 16957 9704
rect 16816 9664 16822 9676
rect 16945 9673 16957 9676
rect 16991 9704 17003 9707
rect 17494 9704 17500 9716
rect 16991 9676 17500 9704
rect 16991 9673 17003 9676
rect 16945 9667 17003 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 11057 9639 11115 9645
rect 11057 9636 11069 9639
rect 11020 9608 11069 9636
rect 11020 9596 11026 9608
rect 11057 9605 11069 9608
rect 11103 9605 11115 9639
rect 11057 9599 11115 9605
rect 11333 9639 11391 9645
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 11379 9608 12940 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 12912 9577 12940 9608
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13044 9608 14044 9636
rect 13044 9596 13050 9608
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9537 9735 9571
rect 9677 9531 9735 9537
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12897 9571 12955 9577
rect 12023 9540 12848 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 6236 9472 6469 9500
rect 6236 9460 6242 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 9030 9500 9036 9512
rect 6604 9472 9036 9500
rect 6604 9460 6610 9472
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9950 9509 9956 9512
rect 9944 9463 9956 9509
rect 10008 9500 10014 9512
rect 12526 9500 12532 9512
rect 10008 9472 10044 9500
rect 10152 9472 12532 9500
rect 9950 9460 9956 9463
rect 10008 9460 10014 9472
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6638 9432 6644 9444
rect 6420 9404 6644 9432
rect 6420 9392 6426 9404
rect 6638 9392 6644 9404
rect 6696 9432 6702 9444
rect 7092 9435 7150 9441
rect 7092 9432 7104 9435
rect 6696 9404 7104 9432
rect 6696 9392 6702 9404
rect 7092 9401 7104 9404
rect 7138 9432 7150 9435
rect 7374 9432 7380 9444
rect 7138 9404 7380 9432
rect 7138 9401 7150 9404
rect 7092 9395 7150 9401
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 9766 9432 9772 9444
rect 9171 9404 9772 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 9858 9392 9864 9444
rect 9916 9432 9922 9444
rect 10152 9432 10180 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12710 9500 12716 9512
rect 12636 9472 12716 9500
rect 11882 9432 11888 9444
rect 9916 9404 10180 9432
rect 10428 9404 11888 9432
rect 9916 9392 9922 9404
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9333 6055 9367
rect 5997 9327 6055 9333
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7708 9336 8217 9364
rect 7708 9324 7714 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 9033 9367 9091 9373
rect 9033 9333 9045 9367
rect 9079 9364 9091 9367
rect 10428 9364 10456 9404
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 11698 9364 11704 9376
rect 9079 9336 10456 9364
rect 11659 9336 11704 9364
rect 9079 9333 9091 9336
rect 9033 9327 9091 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 12158 9364 12164 9376
rect 11839 9336 12164 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12636 9364 12664 9472
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 12820 9500 12848 9540
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13004 9500 13032 9596
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13722 9568 13728 9580
rect 13127 9540 13728 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 13906 9568 13912 9580
rect 13867 9540 13912 9568
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14016 9577 14044 9608
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 15378 9636 15384 9648
rect 14792 9608 15384 9636
rect 14792 9596 14798 9608
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14918 9568 14924 9580
rect 14001 9531 14059 9537
rect 14108 9540 14924 9568
rect 12820 9472 13032 9500
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 14108 9500 14136 9540
rect 14918 9528 14924 9540
rect 14976 9568 14982 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14976 9540 15025 9568
rect 14976 9528 14982 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15160 9540 15577 9568
rect 15160 9528 15166 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 13688 9472 14136 9500
rect 13688 9460 13694 9472
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14516 9472 14841 9500
rect 14516 9460 14522 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 15832 9503 15890 9509
rect 15832 9469 15844 9503
rect 15878 9500 15890 9503
rect 16298 9500 16304 9512
rect 15878 9472 16304 9500
rect 15878 9469 15890 9472
rect 15832 9463 15890 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16632 9472 17417 9500
rect 16632 9460 16638 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17920 9472 18061 9500
rect 17920 9460 17926 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 13817 9435 13875 9441
rect 12851 9404 13492 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 13464 9373 13492 9404
rect 13817 9401 13829 9435
rect 13863 9432 13875 9435
rect 13863 9404 14504 9432
rect 13863 9401 13875 9404
rect 13817 9395 13875 9401
rect 14476 9373 14504 9404
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 14608 9404 14933 9432
rect 14608 9392 14614 9404
rect 14921 9401 14933 9404
rect 14967 9432 14979 9435
rect 15654 9432 15660 9444
rect 14967 9404 15660 9432
rect 14967 9401 14979 9404
rect 14921 9395 14979 9401
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 12483 9336 12664 9364
rect 13449 9367 13507 9373
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 13449 9333 13461 9367
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 14461 9367 14519 9373
rect 14461 9333 14473 9367
rect 14507 9333 14519 9367
rect 17586 9364 17592 9376
rect 17547 9336 17592 9364
rect 14461 9327 14519 9333
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 18230 9364 18236 9376
rect 18191 9336 18236 9364
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 3142 9160 3148 9172
rect 1679 9132 3148 9160
rect 1679 9101 1707 9132
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 4948 9132 5457 9160
rect 4948 9120 4954 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 7374 9160 7380 9172
rect 5445 9123 5503 9129
rect 5552 9132 6868 9160
rect 7335 9132 7380 9160
rect 1664 9095 1722 9101
rect 1664 9061 1676 9095
rect 1710 9061 1722 9095
rect 3418 9092 3424 9104
rect 1664 9055 1722 9061
rect 3068 9064 3424 9092
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 1946 8984 1952 9036
rect 2004 9024 2010 9036
rect 3068 9033 3096 9064
rect 3418 9052 3424 9064
rect 3476 9092 3482 9104
rect 5552 9092 5580 9132
rect 6840 9092 6868 9132
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7484 9132 8892 9160
rect 7484 9092 7512 9132
rect 3476 9064 5580 9092
rect 6012 9064 6776 9092
rect 6840 9064 7512 9092
rect 8196 9095 8254 9101
rect 3476 9052 3482 9064
rect 3053 9027 3111 9033
rect 2004 8996 3004 9024
rect 2004 8984 2010 8996
rect 2976 8956 3004 8996
rect 3053 8993 3065 9027
rect 3099 8993 3111 9027
rect 3053 8987 3111 8993
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 4338 9033 4344 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3660 8996 4077 9024
rect 3660 8984 3666 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4332 9024 4344 9033
rect 4299 8996 4344 9024
rect 4065 8987 4123 8993
rect 4332 8987 4344 8996
rect 4338 8984 4344 8987
rect 4396 8984 4402 9036
rect 6012 9033 6040 9064
rect 6748 9036 6776 9064
rect 8196 9061 8208 9095
rect 8242 9092 8254 9095
rect 8754 9092 8760 9104
rect 8242 9064 8760 9092
rect 8242 9061 8254 9064
rect 8196 9055 8254 9061
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 8864 9092 8892 9132
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 9180 9132 9321 9160
rect 9180 9120 9186 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 10410 9160 10416 9172
rect 9723 9132 10416 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 12529 9163 12587 9169
rect 12529 9160 12541 9163
rect 12216 9132 12541 9160
rect 12216 9120 12222 9132
rect 12529 9129 12541 9132
rect 12575 9129 12587 9163
rect 14918 9160 14924 9172
rect 14879 9132 14924 9160
rect 12529 9123 12587 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 10962 9101 10968 9104
rect 10505 9095 10563 9101
rect 8864 9064 10180 9092
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 8993 6055 9027
rect 6264 9027 6322 9033
rect 6264 9024 6276 9027
rect 5997 8987 6055 8993
rect 6104 8996 6276 9024
rect 3142 8956 3148 8968
rect 2976 8928 3148 8956
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 6104 8956 6132 8996
rect 6264 8993 6276 8996
rect 6310 9024 6322 9027
rect 6546 9024 6552 9036
rect 6310 8996 6552 9024
rect 6310 8993 6322 8996
rect 6264 8987 6322 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7834 9024 7840 9036
rect 6788 8996 7840 9024
rect 6788 8984 6794 8996
rect 7834 8984 7840 8996
rect 7892 9024 7898 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7892 8996 7941 9024
rect 7892 8984 7898 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 9858 9024 9864 9036
rect 7929 8987 7987 8993
rect 8036 8996 9864 9024
rect 5592 8928 6132 8956
rect 5592 8916 5598 8928
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 8036 8956 8064 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10152 9024 10180 9064
rect 10505 9061 10517 9095
rect 10551 9092 10563 9095
rect 10956 9092 10968 9101
rect 10551 9064 10968 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 10956 9055 10968 9064
rect 10962 9052 10968 9055
rect 11020 9052 11026 9104
rect 13446 9092 13452 9104
rect 11072 9064 13452 9092
rect 11072 9024 11100 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 14826 9092 14832 9104
rect 13556 9064 14832 9092
rect 12894 9024 12900 9036
rect 10152 8996 11100 9024
rect 12855 8996 12900 9024
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13556 9033 13584 9064
rect 14826 9052 14832 9064
rect 14884 9092 14890 9104
rect 15102 9092 15108 9104
rect 14884 9064 15108 9092
rect 14884 9052 14890 9064
rect 15102 9052 15108 9064
rect 15160 9092 15166 9104
rect 16758 9101 16764 9104
rect 16752 9092 16764 9101
rect 15160 9064 16528 9092
rect 16719 9064 16764 9092
rect 15160 9052 15166 9064
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 13808 9027 13866 9033
rect 13808 8993 13820 9027
rect 13854 9024 13866 9027
rect 14366 9024 14372 9036
rect 13854 8996 14372 9024
rect 13854 8993 13866 8996
rect 13808 8987 13866 8993
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 15841 9027 15899 9033
rect 15841 9024 15853 9027
rect 15712 8996 15853 9024
rect 15712 8984 15718 8996
rect 15841 8993 15853 8996
rect 15887 8993 15899 9027
rect 15841 8987 15899 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16298 9024 16304 9036
rect 15979 8996 16304 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 16500 9033 16528 9064
rect 16752 9055 16764 9064
rect 16758 9052 16764 9055
rect 16816 9052 16822 9104
rect 16485 9027 16543 9033
rect 16485 8993 16497 9027
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 7064 8928 8064 8956
rect 10137 8959 10195 8965
rect 7064 8916 7070 8928
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10226 8956 10232 8968
rect 10183 8928 10232 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10367 8928 10517 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10686 8956 10692 8968
rect 10647 8928 10692 8956
rect 10505 8919 10563 8925
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 8996 8860 9444 8888
rect 8996 8848 9002 8860
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 2777 8823 2835 8829
rect 2777 8820 2789 8823
rect 2740 8792 2789 8820
rect 2740 8780 2746 8792
rect 2777 8789 2789 8792
rect 2823 8789 2835 8823
rect 2777 8783 2835 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3108 8792 3249 8820
rect 3108 8780 3114 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 4798 8820 4804 8832
rect 3660 8792 4804 8820
rect 3660 8780 3666 8792
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 7926 8820 7932 8832
rect 6052 8792 7932 8820
rect 6052 8780 6058 8792
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 9416 8820 9444 8860
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 10336 8888 10364 8919
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 11848 8928 13001 8956
rect 11848 8916 11854 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13262 8956 13268 8968
rect 13219 8928 13268 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13262 8916 13268 8928
rect 13320 8956 13326 8968
rect 13648 8956 13676 8984
rect 16114 8956 16120 8968
rect 13320 8928 13676 8956
rect 16075 8928 16120 8956
rect 13320 8916 13326 8928
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 9824 8860 10364 8888
rect 15304 8860 16528 8888
rect 9824 8848 9830 8860
rect 11054 8820 11060 8832
rect 9416 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 15304 8820 15332 8860
rect 15470 8820 15476 8832
rect 12584 8792 15332 8820
rect 15431 8792 15476 8820
rect 12584 8780 12590 8792
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 16500 8820 16528 8860
rect 17678 8820 17684 8832
rect 16500 8792 17684 8820
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 17862 8820 17868 8832
rect 17823 8792 17868 8820
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 1397 8619 1455 8625
rect 1397 8585 1409 8619
rect 1443 8616 1455 8619
rect 3602 8616 3608 8628
rect 1443 8588 3608 8616
rect 1443 8585 1455 8588
rect 1397 8579 1455 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 4338 8616 4344 8628
rect 3835 8588 4344 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 6730 8616 6736 8628
rect 4755 8588 6736 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7009 8619 7067 8625
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 7282 8616 7288 8628
rect 7055 8588 7288 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8938 8616 8944 8628
rect 8343 8588 8944 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9766 8616 9772 8628
rect 9232 8588 9772 8616
rect 5721 8551 5779 8557
rect 5721 8517 5733 8551
rect 5767 8548 5779 8551
rect 5767 8520 7512 8548
rect 5767 8517 5779 8520
rect 5721 8511 5779 8517
rect 1486 8440 1492 8492
rect 1544 8480 1550 8492
rect 1854 8480 1860 8492
rect 1544 8452 1860 8480
rect 1544 8440 1550 8452
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2222 8480 2228 8492
rect 2087 8452 2228 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 2406 8480 2412 8492
rect 2367 8452 2412 8480
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 4706 8480 4712 8492
rect 3896 8452 4712 8480
rect 1302 8372 1308 8424
rect 1360 8412 1366 8424
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 1360 8384 1777 8412
rect 1360 8372 1366 8384
rect 1765 8381 1777 8384
rect 1811 8412 1823 8415
rect 3896 8412 3924 8452
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 4948 8452 5181 8480
rect 4948 8440 4954 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5534 8480 5540 8492
rect 5399 8452 5540 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 6362 8480 6368 8492
rect 6323 8452 6368 8480
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 7006 8480 7012 8492
rect 6595 8452 7012 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7484 8489 7512 8520
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7650 8480 7656 8492
rect 7611 8452 7656 8480
rect 7469 8443 7527 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8480 8999 8483
rect 9232 8480 9260 8588
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 11756 8588 12633 8616
rect 11756 8576 11762 8588
rect 12621 8585 12633 8588
rect 12667 8585 12679 8619
rect 12621 8579 12679 8585
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16485 8619 16543 8625
rect 16485 8616 16497 8619
rect 16356 8588 16497 8616
rect 16356 8576 16362 8588
rect 16485 8585 16497 8588
rect 16531 8585 16543 8619
rect 16485 8579 16543 8585
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 9582 8548 9588 8560
rect 9355 8520 9588 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 10137 8551 10195 8557
rect 10137 8548 10149 8551
rect 9876 8520 10149 8548
rect 9876 8480 9904 8520
rect 10137 8517 10149 8520
rect 10183 8517 10195 8551
rect 10137 8511 10195 8517
rect 10321 8551 10379 8557
rect 10321 8517 10333 8551
rect 10367 8548 10379 8551
rect 10502 8548 10508 8560
rect 10367 8520 10508 8548
rect 10367 8517 10379 8520
rect 10321 8511 10379 8517
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 18233 8551 18291 8557
rect 11379 8520 13124 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 8987 8452 9260 8480
rect 9324 8452 9904 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 4062 8412 4068 8424
rect 1811 8384 3924 8412
rect 3975 8384 4068 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2682 8353 2688 8356
rect 2654 8347 2688 8353
rect 2654 8344 2666 8347
rect 2280 8316 2666 8344
rect 2280 8304 2286 8316
rect 2654 8313 2666 8316
rect 2740 8344 2746 8356
rect 2740 8316 2802 8344
rect 2654 8307 2688 8313
rect 2682 8304 2688 8307
rect 2740 8304 2746 8316
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 3988 8344 4016 8384
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4856 8384 5089 8412
rect 4856 8372 4862 8384
rect 5077 8381 5089 8384
rect 5123 8412 5135 8415
rect 5123 8384 5396 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 3200 8316 4016 8344
rect 4080 8316 4384 8344
rect 3200 8304 3206 8316
rect 1854 8236 1860 8288
rect 1912 8276 1918 8288
rect 4080 8276 4108 8316
rect 4246 8276 4252 8288
rect 1912 8248 4108 8276
rect 4207 8248 4252 8276
rect 1912 8236 1918 8248
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4356 8276 4384 8316
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 5368 8344 5396 8384
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 6052 8384 6101 8412
rect 6052 8372 6058 8384
rect 6089 8381 6101 8384
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 8018 8412 8024 8424
rect 6227 8384 8024 8412
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8754 8412 8760 8424
rect 8444 8384 8760 8412
rect 8444 8372 8450 8384
rect 8754 8372 8760 8384
rect 8812 8412 8818 8424
rect 9324 8412 9352 8452
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10008 8452 10053 8480
rect 10612 8452 10793 8480
rect 10008 8440 10014 8452
rect 8812 8384 9352 8412
rect 9769 8415 9827 8421
rect 8812 8372 8818 8384
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10134 8412 10140 8424
rect 9815 8384 10140 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8412 10287 8415
rect 10612 8412 10640 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10962 8480 10968 8492
rect 10875 8452 10968 8480
rect 10781 8443 10839 8449
rect 10962 8440 10968 8452
rect 11020 8480 11026 8492
rect 13096 8489 13124 8520
rect 18233 8517 18245 8551
rect 18279 8548 18291 8551
rect 18322 8548 18328 8560
rect 18279 8520 18328 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18322 8508 18328 8520
rect 18380 8508 18386 8560
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11020 8452 11989 8480
rect 11020 8440 11026 8452
rect 11977 8449 11989 8452
rect 12023 8480 12035 8483
rect 13081 8483 13139 8489
rect 12023 8452 12388 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 10275 8384 10640 8412
rect 10689 8415 10747 8421
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 11146 8412 11152 8424
rect 10735 8384 11152 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 11146 8372 11152 8384
rect 11204 8372 11210 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11296 8384 11805 8412
rect 11296 8372 11302 8384
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 4488 8316 5120 8344
rect 5368 8316 6561 8344
rect 4488 8304 4494 8316
rect 4982 8276 4988 8288
rect 4356 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 5092 8276 5120 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 6880 8316 7389 8344
rect 6880 8304 6886 8316
rect 7377 8313 7389 8316
rect 7423 8313 7435 8347
rect 7377 8307 7435 8313
rect 9677 8347 9735 8353
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 11054 8344 11060 8356
rect 9723 8316 11060 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 12360 8344 12388 8452
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13262 8480 13268 8492
rect 13223 8452 13268 8480
rect 13081 8443 13139 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14550 8480 14556 8492
rect 14507 8452 14556 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14826 8480 14832 8492
rect 14787 8452 14832 8480
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17862 8480 17868 8492
rect 17083 8452 17868 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12676 8384 13001 8412
rect 12676 8372 12682 8384
rect 12989 8381 13001 8384
rect 13035 8381 13047 8415
rect 14274 8412 14280 8424
rect 14187 8384 14280 8412
rect 12989 8375 13047 8381
rect 14274 8372 14280 8384
rect 14332 8412 14338 8424
rect 15096 8415 15154 8421
rect 14332 8384 14780 8412
rect 14332 8372 14338 8384
rect 14366 8344 14372 8356
rect 11624 8316 11928 8344
rect 12360 8316 14372 8344
rect 8110 8276 8116 8288
rect 5092 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8352 8248 8677 8276
rect 8352 8236 8358 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 11238 8276 11244 8288
rect 8904 8248 11244 8276
rect 8904 8236 8910 8248
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 11624 8276 11652 8316
rect 11388 8248 11652 8276
rect 11388 8236 11394 8248
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 11900 8276 11928 8316
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 14752 8344 14780 8384
rect 15096 8381 15108 8415
rect 15142 8412 15154 8415
rect 17052 8412 17080 8443
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18046 8412 18052 8424
rect 15142 8384 17080 8412
rect 18007 8384 18052 8412
rect 15142 8381 15154 8384
rect 15096 8375 15154 8381
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 17954 8344 17960 8356
rect 14752 8316 17960 8344
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 12158 8276 12164 8288
rect 11756 8248 11801 8276
rect 11900 8248 12164 8276
rect 11756 8236 11762 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13814 8276 13820 8288
rect 13775 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 14185 8279 14243 8285
rect 14185 8245 14197 8279
rect 14231 8276 14243 8279
rect 14734 8276 14740 8288
rect 14231 8248 14740 8276
rect 14231 8245 14243 8248
rect 14185 8239 14243 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 16172 8248 16221 8276
rect 16172 8236 16178 8248
rect 16209 8245 16221 8248
rect 16255 8245 16267 8279
rect 16209 8239 16267 8245
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8276 16911 8279
rect 17034 8276 17040 8288
rect 16899 8248 17040 8276
rect 16899 8245 16911 8248
rect 16853 8239 16911 8245
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 17494 8276 17500 8288
rect 17455 8248 17500 8276
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 3142 8072 3148 8084
rect 1627 8044 3148 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 3418 8072 3424 8084
rect 3379 8044 3424 8072
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 5166 8072 5172 8084
rect 3927 8044 5172 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 5307 8044 6653 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 6788 8044 6833 8072
rect 6788 8032 6794 8044
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 10321 8075 10379 8081
rect 7616 8044 10272 8072
rect 7616 8032 7622 8044
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 8004 2375 8007
rect 5074 8004 5080 8016
rect 2363 7976 5080 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 5629 8007 5687 8013
rect 5629 7973 5641 8007
rect 5675 8004 5687 8007
rect 9677 8007 9735 8013
rect 9677 8004 9689 8007
rect 5675 7976 9689 8004
rect 5675 7973 5687 7976
rect 5629 7967 5687 7973
rect 9677 7973 9689 7976
rect 9723 7973 9735 8007
rect 9677 7967 9735 7973
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3510 7936 3516 7948
rect 3375 7908 3516 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 5258 7936 5264 7948
rect 4663 7908 5264 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 7285 7939 7343 7945
rect 5592 7908 5948 7936
rect 5592 7896 5598 7908
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2222 7760 2228 7812
rect 2280 7800 2286 7812
rect 2516 7800 2544 7831
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3605 7871 3663 7877
rect 3605 7868 3617 7871
rect 3476 7840 3617 7868
rect 3476 7828 3482 7840
rect 3605 7837 3617 7840
rect 3651 7868 3663 7871
rect 4430 7868 4436 7880
rect 3651 7840 4436 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7868 4951 7871
rect 4939 7840 5672 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 3881 7803 3939 7809
rect 3881 7800 3893 7803
rect 2280 7772 2544 7800
rect 2884 7772 3893 7800
rect 2280 7760 2286 7772
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2884 7732 2912 7772
rect 3881 7769 3893 7772
rect 3927 7769 3939 7803
rect 3881 7763 3939 7769
rect 4338 7760 4344 7812
rect 4396 7800 4402 7812
rect 4908 7800 4936 7831
rect 4396 7772 4936 7800
rect 4396 7760 4402 7772
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 5442 7800 5448 7812
rect 5132 7772 5448 7800
rect 5132 7760 5138 7772
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 1995 7704 2912 7732
rect 2961 7735 3019 7741
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 3786 7732 3792 7744
rect 3007 7704 3792 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 5534 7732 5540 7744
rect 4295 7704 5540 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 5644 7732 5672 7840
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 5920 7877 5948 7908
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7558 7936 7564 7948
rect 7331 7908 7564 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7834 7936 7840 7948
rect 7795 7908 7840 7936
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8110 7945 8116 7948
rect 8104 7936 8116 7945
rect 8071 7908 8116 7936
rect 8104 7899 8116 7908
rect 8110 7896 8116 7899
rect 8168 7896 8174 7948
rect 5905 7871 5963 7877
rect 5776 7840 5821 7868
rect 5776 7828 5782 7840
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 6546 7868 6552 7880
rect 5905 7831 5963 7837
rect 6288 7840 6552 7868
rect 6288 7809 6316 7840
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6696 7840 6837 7868
rect 6696 7828 6702 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7742 7868 7748 7880
rect 7432 7840 7748 7868
rect 7432 7828 7438 7840
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 6273 7803 6331 7809
rect 6273 7769 6285 7803
rect 6319 7769 6331 7803
rect 6273 7763 6331 7769
rect 6380 7772 7604 7800
rect 6380 7732 6408 7772
rect 5644 7704 6408 7732
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 6696 7704 7481 7732
rect 6696 7692 6702 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 7576 7732 7604 7772
rect 9214 7732 9220 7744
rect 7576 7704 9220 7732
rect 7469 7695 7527 7701
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 10244 7732 10272 8044
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 11790 8072 11796 8084
rect 10367 8044 11796 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 14182 8072 14188 8084
rect 11900 8044 14188 8072
rect 10778 7964 10784 8016
rect 10836 8004 10842 8016
rect 10836 7976 11376 8004
rect 10836 7964 10842 7976
rect 10502 7896 10508 7948
rect 10560 7936 10566 7948
rect 11348 7945 11376 7976
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 11900 8004 11928 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15194 8072 15200 8084
rect 14875 8044 15200 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 15528 8044 15853 8072
rect 15528 8032 15534 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 15841 8035 15899 8041
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 16807 8044 17417 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17405 8041 17417 8044
rect 17451 8041 17463 8075
rect 17405 8035 17463 8041
rect 11480 7976 11928 8004
rect 11480 7964 11486 7976
rect 12158 7964 12164 8016
rect 12216 8004 12222 8016
rect 15749 8007 15807 8013
rect 12216 7976 14688 8004
rect 12216 7964 12222 7976
rect 10689 7939 10747 7945
rect 10689 7936 10701 7939
rect 10560 7908 10701 7936
rect 10560 7896 10566 7908
rect 10689 7905 10701 7908
rect 10735 7905 10747 7939
rect 10689 7899 10747 7905
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11600 7939 11658 7945
rect 11600 7905 11612 7939
rect 11646 7936 11658 7939
rect 12066 7936 12072 7948
rect 11646 7908 12072 7936
rect 11646 7905 11658 7908
rect 11600 7899 11658 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 14660 7945 14688 7976
rect 15749 7973 15761 8007
rect 15795 8004 15807 8007
rect 16408 8004 16436 8035
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17552 8044 17785 8072
rect 17552 8032 17558 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 15795 7976 16436 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 17862 7964 17868 8016
rect 17920 7964 17926 8016
rect 13245 7939 13303 7945
rect 13245 7936 13257 7939
rect 12728 7908 13257 7936
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10778 7868 10784 7880
rect 10376 7840 10784 7868
rect 10376 7828 10382 7840
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 11256 7800 11284 7828
rect 10928 7772 11284 7800
rect 10928 7760 10934 7772
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12728 7809 12756 7908
rect 13245 7905 13257 7908
rect 13291 7905 13303 7939
rect 13245 7899 13303 7905
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 17880 7936 17908 7964
rect 14645 7899 14703 7905
rect 15304 7908 17080 7936
rect 17880 7908 18000 7936
rect 12986 7868 12992 7880
rect 12947 7840 12992 7868
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 15194 7868 15200 7880
rect 14148 7840 15200 7868
rect 14148 7828 14154 7840
rect 15194 7828 15200 7840
rect 15252 7868 15258 7880
rect 15304 7868 15332 7908
rect 15252 7840 15332 7868
rect 16025 7871 16083 7877
rect 15252 7828 15258 7840
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 16206 7868 16212 7880
rect 16071 7840 16212 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16850 7868 16856 7880
rect 16811 7840 16856 7868
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 17052 7868 17080 7908
rect 17972 7877 18000 7908
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17052 7840 17877 7868
rect 16945 7831 17003 7837
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 12713 7803 12771 7809
rect 12713 7800 12725 7803
rect 12400 7772 12725 7800
rect 12400 7760 12406 7772
rect 12713 7769 12725 7772
rect 12759 7769 12771 7803
rect 15470 7800 15476 7812
rect 12713 7763 12771 7769
rect 13924 7772 15476 7800
rect 12250 7732 12256 7744
rect 10244 7704 12256 7732
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 12802 7732 12808 7744
rect 12676 7704 12808 7732
rect 12676 7692 12682 7704
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13924 7732 13952 7772
rect 15470 7760 15476 7772
rect 15528 7760 15534 7812
rect 16114 7760 16120 7812
rect 16172 7800 16178 7812
rect 16960 7800 16988 7831
rect 16172 7772 16988 7800
rect 16172 7760 16178 7772
rect 13044 7704 13952 7732
rect 13044 7692 13050 7704
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15381 7735 15439 7741
rect 15381 7732 15393 7735
rect 15252 7704 15393 7732
rect 15252 7692 15258 7704
rect 15381 7701 15393 7704
rect 15427 7701 15439 7735
rect 15381 7695 15439 7701
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 1854 7528 1860 7540
rect 1719 7500 1860 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 5810 7528 5816 7540
rect 3743 7500 5816 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6086 7528 6092 7540
rect 6047 7500 6092 7528
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 9030 7528 9036 7540
rect 8864 7500 9036 7528
rect 5718 7420 5724 7472
rect 5776 7460 5782 7472
rect 8864 7460 8892 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10502 7528 10508 7540
rect 10284 7500 10508 7528
rect 10284 7488 10290 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 12069 7531 12127 7537
rect 12069 7497 12081 7531
rect 12115 7528 12127 7531
rect 15562 7528 15568 7540
rect 12115 7500 15568 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 16206 7528 16212 7540
rect 16167 7500 16212 7528
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 16908 7500 16957 7528
rect 16908 7488 16914 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 16945 7491 17003 7497
rect 5776 7432 8892 7460
rect 5776 7420 5782 7432
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 12434 7460 12440 7472
rect 8996 7432 12440 7460
rect 8996 7420 9002 7432
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 12618 7420 12624 7472
rect 12676 7460 12682 7472
rect 12676 7432 13952 7460
rect 12676 7420 12682 7432
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7392 3387 7395
rect 3418 7392 3424 7404
rect 3375 7364 3424 7392
rect 3375 7361 3387 7364
rect 3329 7355 3387 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3844 7364 4169 7392
rect 3844 7352 3850 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 4157 7355 4215 7361
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 4430 7352 4436 7404
rect 4488 7392 4494 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4488 7364 4721 7392
rect 4488 7352 4494 7364
rect 4709 7361 4721 7364
rect 4755 7361 4767 7395
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 4709 7355 4767 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 7760 7364 10701 7392
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 2130 7324 2136 7336
rect 2087 7296 2136 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2130 7284 2136 7296
rect 2188 7284 2194 7336
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 3878 7324 3884 7336
rect 3099 7296 3884 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7760 7324 7788 7364
rect 10689 7361 10701 7364
rect 10735 7392 10747 7395
rect 11514 7392 11520 7404
rect 10735 7364 11520 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11698 7392 11704 7404
rect 11659 7364 11704 7392
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 13170 7392 13176 7404
rect 12452 7364 13176 7392
rect 6687 7296 7788 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7834 7284 7840 7336
rect 7892 7324 7898 7336
rect 8202 7324 8208 7336
rect 7892 7296 8208 7324
rect 7892 7284 7898 7296
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8938 7324 8944 7336
rect 8899 7296 8944 7324
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 11808 7324 11836 7352
rect 12452 7336 12480 7364
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7361 13875 7395
rect 13924 7392 13952 7432
rect 13924 7364 14964 7392
rect 13817 7355 13875 7361
rect 9088 7296 11836 7324
rect 9088 7284 9094 7296
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 11940 7296 11985 7324
rect 11940 7284 11946 7296
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 12802 7324 12808 7336
rect 12759 7296 12808 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 13044 7296 13093 7324
rect 13044 7284 13050 7296
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 13630 7324 13636 7336
rect 13591 7296 13636 7324
rect 13081 7287 13139 7293
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13832 7324 13860 7355
rect 14090 7324 14096 7336
rect 13832 7296 14096 7324
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14826 7324 14832 7336
rect 14787 7296 14832 7324
rect 14277 7287 14335 7293
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 2700 7228 4077 7256
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2590 7188 2596 7200
rect 2179 7160 2596 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 2700 7197 2728 7228
rect 4065 7225 4077 7228
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 4976 7259 5034 7265
rect 4976 7225 4988 7259
rect 5022 7256 5034 7259
rect 5442 7256 5448 7268
rect 5022 7228 5448 7256
rect 5022 7225 5034 7228
rect 4976 7219 5034 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 6328 7228 7205 7256
rect 6328 7216 6334 7228
rect 7193 7225 7205 7228
rect 7239 7256 7251 7259
rect 8846 7256 8852 7268
rect 7239 7228 8852 7256
rect 7239 7225 7251 7228
rect 7193 7219 7251 7225
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 9766 7216 9772 7268
rect 9824 7256 9830 7268
rect 11238 7256 11244 7268
rect 9824 7228 11244 7256
rect 9824 7216 9830 7228
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 11425 7259 11483 7265
rect 11425 7225 11437 7259
rect 11471 7256 11483 7259
rect 12618 7256 12624 7268
rect 11471 7228 12624 7256
rect 11471 7225 11483 7228
rect 11425 7219 11483 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 13725 7259 13783 7265
rect 12820 7228 13400 7256
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7157 2743 7191
rect 2685 7151 2743 7157
rect 3145 7191 3203 7197
rect 3145 7157 3157 7191
rect 3191 7188 3203 7191
rect 5718 7188 5724 7200
rect 3191 7160 5724 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 6178 7148 6184 7200
rect 6236 7188 6242 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 6236 7160 6469 7188
rect 6236 7148 6242 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6604 7160 6837 7188
rect 6604 7148 6610 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7926 7188 7932 7200
rect 7331 7160 7932 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 8076 7160 8121 7188
rect 8076 7148 8082 7160
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 11330 7188 11336 7200
rect 8260 7160 11336 7188
rect 8260 7148 8266 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11974 7188 11980 7200
rect 11563 7160 11980 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12820 7188 12848 7228
rect 12216 7160 12848 7188
rect 12897 7191 12955 7197
rect 12216 7148 12222 7160
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 13081 7191 13139 7197
rect 13081 7188 13093 7191
rect 12943 7160 13093 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13081 7157 13093 7160
rect 13127 7157 13139 7191
rect 13262 7188 13268 7200
rect 13223 7160 13268 7188
rect 13081 7151 13139 7157
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 13372 7188 13400 7228
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 13814 7256 13820 7268
rect 13771 7228 13820 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14292 7188 14320 7287
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 14936 7324 14964 7364
rect 16574 7352 16580 7404
rect 16632 7352 16638 7404
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 17589 7395 17647 7401
rect 17589 7392 17601 7395
rect 16724 7364 17601 7392
rect 16724 7352 16730 7364
rect 17589 7361 17601 7364
rect 17635 7392 17647 7395
rect 17862 7392 17868 7404
rect 17635 7364 17868 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 16485 7327 16543 7333
rect 16485 7324 16497 7327
rect 14936 7296 16497 7324
rect 16485 7293 16497 7296
rect 16531 7293 16543 7327
rect 16485 7287 16543 7293
rect 15096 7259 15154 7265
rect 15096 7225 15108 7259
rect 15142 7256 15154 7259
rect 16114 7256 16120 7268
rect 15142 7228 16120 7256
rect 15142 7225 15154 7228
rect 15096 7219 15154 7225
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 16592 7256 16620 7352
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 17678 7324 17684 7336
rect 17359 7296 17684 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 18012 7296 18061 7324
rect 18012 7284 18018 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 16592 7228 17417 7256
rect 17405 7225 17417 7228
rect 17451 7225 17463 7259
rect 17405 7219 17463 7225
rect 13372 7160 14320 7188
rect 14461 7191 14519 7197
rect 14461 7157 14473 7191
rect 14507 7188 14519 7191
rect 15378 7188 15384 7200
rect 14507 7160 15384 7188
rect 14507 7157 14519 7160
rect 14461 7151 14519 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 18230 7188 18236 7200
rect 18191 7160 18236 7188
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 7926 6984 7932 6996
rect 5592 6956 7932 6984
rect 5592 6944 5598 6956
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 9766 6984 9772 6996
rect 8628 6956 9772 6984
rect 8628 6944 8634 6956
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 9916 6956 10241 6984
rect 9916 6944 9922 6956
rect 10229 6953 10241 6956
rect 10275 6953 10287 6987
rect 11698 6984 11704 6996
rect 10229 6947 10287 6953
rect 11155 6956 11704 6984
rect 3510 6916 3516 6928
rect 3344 6888 3516 6916
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 3344 6857 3372 6888
rect 3510 6876 3516 6888
rect 3568 6916 3574 6928
rect 8380 6919 8438 6925
rect 3568 6888 7512 6916
rect 3568 6876 3574 6888
rect 1929 6851 1987 6857
rect 1929 6848 1941 6851
rect 1820 6820 1941 6848
rect 1820 6808 1826 6820
rect 1929 6817 1941 6820
rect 1975 6817 1987 6851
rect 1929 6811 1987 6817
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6817 3387 6851
rect 4614 6848 4620 6860
rect 3329 6811 3387 6817
rect 3436 6820 4620 6848
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1452 6752 1685 6780
rect 1452 6740 1458 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 3436 6724 3464 6820
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 4792 6851 4850 6857
rect 4792 6817 4804 6851
rect 4838 6848 4850 6851
rect 6540 6851 6598 6857
rect 4838 6820 6224 6848
rect 4838 6817 4850 6820
rect 4792 6811 4850 6817
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 3418 6712 3424 6724
rect 3099 6684 3424 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 3513 6647 3571 6653
rect 3513 6613 3525 6647
rect 3559 6644 3571 6647
rect 3602 6644 3608 6656
rect 3559 6616 3608 6644
rect 3559 6613 3571 6616
rect 3513 6607 3571 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 4080 6644 4108 6743
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4488 6752 4537 6780
rect 4488 6740 4494 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 5626 6644 5632 6656
rect 4080 6616 5632 6644
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6196 6644 6224 6820
rect 6540 6817 6552 6851
rect 6586 6848 6598 6851
rect 7374 6848 7380 6860
rect 6586 6820 7380 6848
rect 6586 6817 6598 6820
rect 6540 6811 6598 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 7484 6848 7512 6888
rect 8380 6885 8392 6919
rect 8426 6916 8438 6919
rect 9214 6916 9220 6928
rect 8426 6888 9220 6916
rect 8426 6885 8438 6888
rect 8380 6879 8438 6885
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 11155 6925 11183 6956
rect 11698 6944 11704 6956
rect 11756 6984 11762 6996
rect 11756 6956 13216 6984
rect 11756 6944 11762 6956
rect 11140 6919 11198 6925
rect 11140 6885 11152 6919
rect 11186 6885 11198 6919
rect 11140 6879 11198 6885
rect 13188 6916 13216 6956
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 13814 6984 13820 6996
rect 13320 6956 13820 6984
rect 13320 6944 13326 6956
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 14148 6956 14933 6984
rect 14148 6944 14154 6956
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 17770 6984 17776 6996
rect 16632 6956 17776 6984
rect 16632 6944 16638 6956
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 14108 6916 14136 6944
rect 13188 6888 14136 6916
rect 10410 6848 10416 6860
rect 7484 6820 10416 6848
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 12342 6848 12348 6860
rect 10520 6820 12348 6848
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 8110 6780 8116 6792
rect 6328 6752 6373 6780
rect 8071 6752 8116 6780
rect 6328 6740 6334 6752
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10520 6789 10548 6820
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12894 6848 12900 6860
rect 12855 6820 12900 6848
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13188 6789 13216 6888
rect 14826 6876 14832 6928
rect 14884 6916 14890 6928
rect 16016 6919 16074 6925
rect 14884 6888 15056 6916
rect 14884 6876 14890 6888
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 13797 6851 13855 6857
rect 13797 6848 13809 6851
rect 13504 6820 13809 6848
rect 13504 6808 13510 6820
rect 13797 6817 13809 6820
rect 13843 6817 13855 6851
rect 15028 6848 15056 6888
rect 16016 6885 16028 6919
rect 16062 6916 16074 6919
rect 16206 6916 16212 6928
rect 16062 6888 16212 6916
rect 16062 6885 16074 6888
rect 16016 6879 16074 6885
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 15028 6820 15761 6848
rect 13797 6811 13855 6817
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 17678 6848 17684 6860
rect 15749 6811 15807 6817
rect 15856 6820 17684 6848
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 9766 6672 9772 6724
rect 9824 6712 9830 6724
rect 10888 6712 10916 6743
rect 9824 6684 10916 6712
rect 9824 6672 9830 6684
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 12253 6715 12311 6721
rect 12253 6712 12265 6715
rect 12124 6684 12265 6712
rect 12124 6672 12130 6684
rect 12253 6681 12265 6684
rect 12299 6681 12311 6715
rect 12253 6675 12311 6681
rect 6454 6644 6460 6656
rect 6196 6616 6460 6644
rect 6454 6604 6460 6616
rect 6512 6644 6518 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 6512 6616 7665 6644
rect 6512 6604 6518 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 7653 6607 7711 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 12158 6644 12164 6656
rect 9907 6616 12164 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 13004 6644 13032 6743
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13412 6752 13553 6780
rect 13412 6740 13418 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15160 6752 15301 6780
rect 15160 6740 15166 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15856 6780 15884 6820
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 17862 6780 17868 6792
rect 15289 6743 15347 6749
rect 15764 6752 15884 6780
rect 17823 6752 17868 6780
rect 13906 6644 13912 6656
rect 13004 6616 13912 6644
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 15764 6644 15792 6752
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 16684 6684 17417 6712
rect 14332 6616 15792 6644
rect 14332 6604 14338 6616
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 16684 6644 16712 6684
rect 17405 6681 17417 6684
rect 17451 6681 17463 6715
rect 17405 6675 17463 6681
rect 17770 6672 17776 6724
rect 17828 6712 17834 6724
rect 17972 6712 18000 6743
rect 17828 6684 18000 6712
rect 17828 6672 17834 6684
rect 17126 6644 17132 6656
rect 16448 6616 16712 6644
rect 17087 6616 17132 6644
rect 16448 6604 16454 6616
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 1946 6440 1952 6452
rect 1820 6412 1952 6440
rect 1820 6400 1826 6412
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 4338 6440 4344 6452
rect 2700 6412 4344 6440
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 1452 6344 2636 6372
rect 1452 6332 1458 6344
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2314 6304 2320 6316
rect 2188 6276 2320 6304
rect 2188 6264 2194 6276
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6236 1547 6239
rect 1762 6236 1768 6248
rect 1535 6208 1768 6236
rect 1535 6205 1547 6208
rect 1489 6199 1547 6205
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2498 6236 2504 6248
rect 2455 6208 2504 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 2608 6236 2636 6344
rect 2700 6313 2728 6412
rect 4338 6400 4344 6412
rect 4396 6440 4402 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4396 6412 4445 6440
rect 4396 6400 4402 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 8110 6440 8116 6452
rect 6788 6412 8116 6440
rect 6788 6400 6794 6412
rect 8110 6400 8116 6412
rect 8168 6440 8174 6452
rect 8757 6443 8815 6449
rect 8168 6412 8616 6440
rect 8168 6400 8174 6412
rect 7929 6375 7987 6381
rect 7929 6372 7941 6375
rect 4632 6344 6316 6372
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 2608 6208 3065 6236
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 2958 6168 2964 6180
rect 1780 6140 2964 6168
rect 1673 6103 1731 6109
rect 1673 6069 1685 6103
rect 1719 6100 1731 6103
rect 1780 6100 1808 6140
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 2038 6100 2044 6112
rect 1719 6072 1808 6100
rect 1999 6072 2044 6100
rect 1719 6069 1731 6072
rect 1673 6063 1731 6069
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 2280 6072 2513 6100
rect 2280 6060 2286 6072
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 3068 6100 3096 6199
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 4632 6236 4660 6344
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5500 6276 5641 6304
rect 5500 6264 5506 6276
rect 5629 6273 5641 6276
rect 5675 6304 5687 6307
rect 5902 6304 5908 6316
rect 5675 6276 5908 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 4120 6208 4660 6236
rect 4985 6239 5043 6245
rect 4120 6196 4126 6208
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 6178 6236 6184 6248
rect 5031 6208 6184 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 6288 6236 6316 6344
rect 6380 6344 7941 6372
rect 6380 6313 6408 6344
rect 7929 6341 7941 6344
rect 7975 6341 7987 6375
rect 7929 6335 7987 6341
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6512 6276 6557 6304
rect 6512 6264 6518 6276
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7432 6276 7665 6304
rect 7432 6264 7438 6276
rect 7653 6273 7665 6276
rect 7699 6304 7711 6307
rect 8202 6304 8208 6316
rect 7699 6276 8208 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 8202 6264 8208 6276
rect 8260 6304 8266 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8260 6276 8493 6304
rect 8260 6264 8266 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8588 6304 8616 6412
rect 8757 6409 8769 6443
rect 8803 6440 8815 6443
rect 10962 6440 10968 6452
rect 8803 6412 10968 6440
rect 8803 6409 8815 6412
rect 8757 6403 8815 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 11146 6440 11152 6452
rect 11107 6412 11152 6440
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 12250 6440 12256 6452
rect 11296 6412 12256 6440
rect 11296 6400 11302 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 12894 6440 12900 6452
rect 12851 6412 12900 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 14642 6440 14648 6452
rect 13412 6412 14648 6440
rect 13412 6400 13418 6412
rect 14642 6400 14648 6412
rect 14700 6440 14706 6452
rect 14826 6440 14832 6452
rect 14700 6412 14832 6440
rect 14700 6400 14706 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 15712 6412 15853 6440
rect 15712 6400 15718 6412
rect 15841 6409 15853 6412
rect 15887 6409 15899 6443
rect 15841 6403 15899 6409
rect 10318 6332 10324 6384
rect 10376 6372 10382 6384
rect 13630 6372 13636 6384
rect 10376 6344 13636 6372
rect 10376 6332 10382 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6372 13875 6375
rect 17862 6372 17868 6384
rect 13863 6344 17868 6372
rect 13863 6341 13875 6344
rect 13817 6335 13875 6341
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8588 6276 8861 6304
rect 8481 6267 8539 6273
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 8849 6267 8907 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13265 6307 13323 6313
rect 13265 6304 13277 6307
rect 13228 6276 13277 6304
rect 13228 6264 13234 6276
rect 13265 6273 13277 6276
rect 13311 6273 13323 6307
rect 13446 6304 13452 6316
rect 13359 6276 13452 6304
rect 13265 6267 13323 6273
rect 13446 6264 13452 6276
rect 13504 6304 13510 6316
rect 13504 6276 14228 6304
rect 13504 6264 13510 6276
rect 7466 6236 7472 6248
rect 6288 6208 7236 6236
rect 7427 6208 7472 6236
rect 3320 6171 3378 6177
rect 3320 6137 3332 6171
rect 3366 6168 3378 6171
rect 3418 6168 3424 6180
rect 3366 6140 3424 6168
rect 3366 6137 3378 6140
rect 3320 6131 3378 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 7208 6168 7236 6208
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 8110 6236 8116 6248
rect 7616 6208 8116 6236
rect 7616 6196 7622 6208
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6236 8355 6239
rect 8570 6236 8576 6248
rect 8343 6208 8576 6236
rect 8343 6205 8355 6208
rect 8297 6199 8355 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9116 6239 9174 6245
rect 9116 6205 9128 6239
rect 9162 6236 9174 6239
rect 9490 6236 9496 6248
rect 9162 6208 9496 6236
rect 9162 6205 9174 6208
rect 9116 6199 9174 6205
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9640 6208 10517 6236
rect 9640 6196 9646 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 11020 6208 12480 6236
rect 11020 6196 11026 6208
rect 8478 6168 8484 6180
rect 5491 6140 5948 6168
rect 7208 6140 8484 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 4062 6100 4068 6112
rect 3068 6072 4068 6100
rect 2501 6063 2559 6069
rect 4062 6060 4068 6072
rect 4120 6100 4126 6112
rect 4430 6100 4436 6112
rect 4120 6072 4436 6100
rect 4120 6060 4126 6072
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 4948 6072 5089 6100
rect 4948 6060 4954 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5537 6103 5595 6109
rect 5537 6069 5549 6103
rect 5583 6100 5595 6103
rect 5718 6100 5724 6112
rect 5583 6072 5724 6100
rect 5583 6069 5595 6072
rect 5537 6063 5595 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5920 6109 5948 6140
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 10318 6128 10324 6180
rect 10376 6168 10382 6180
rect 11606 6168 11612 6180
rect 10376 6140 11612 6168
rect 10376 6128 10382 6140
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 12452 6168 12480 6208
rect 12526 6196 12532 6248
rect 12584 6236 12590 6248
rect 14090 6236 14096 6248
rect 12584 6208 14096 6236
rect 12584 6196 12590 6208
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14200 6236 14228 6276
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14461 6307 14519 6313
rect 14332 6276 14377 6304
rect 14332 6264 14338 6276
rect 14461 6273 14473 6307
rect 14507 6304 14519 6307
rect 14918 6304 14924 6316
rect 14507 6276 14924 6304
rect 14507 6273 14519 6276
rect 14461 6267 14519 6273
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 15286 6304 15292 6316
rect 15247 6276 15292 6304
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16390 6304 16396 6316
rect 16347 6276 16396 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 14550 6236 14556 6248
rect 14200 6208 14556 6236
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15488 6236 15516 6267
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16666 6304 16672 6316
rect 16531 6276 16672 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 17313 6307 17371 6313
rect 17313 6273 17325 6307
rect 17359 6304 17371 6307
rect 17402 6304 17408 6316
rect 17359 6276 17408 6304
rect 17359 6273 17371 6276
rect 17313 6267 17371 6273
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 17770 6304 17776 6316
rect 17543 6276 17776 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 17512 6236 17540 6267
rect 17770 6264 17776 6276
rect 17828 6264 17834 6316
rect 15488 6208 17540 6236
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17736 6208 18061 6236
rect 17736 6196 17742 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 15197 6171 15255 6177
rect 12452 6140 13400 6168
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6273 6103 6331 6109
rect 6273 6069 6285 6103
rect 6319 6100 6331 6103
rect 7101 6103 7159 6109
rect 7101 6100 7113 6103
rect 6319 6072 7113 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 7101 6069 7113 6072
rect 7147 6069 7159 6103
rect 8386 6100 8392 6112
rect 8347 6072 8392 6100
rect 7101 6063 7159 6069
rect 8386 6060 8392 6072
rect 8444 6100 8450 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8444 6072 8769 6100
rect 8444 6060 8450 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 10008 6072 10241 6100
rect 10008 6060 10014 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10229 6063 10287 6069
rect 11517 6103 11575 6109
rect 11517 6069 11529 6103
rect 11563 6100 11575 6103
rect 11790 6100 11796 6112
rect 11563 6072 11796 6100
rect 11563 6069 11575 6072
rect 11517 6063 11575 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13372 6100 13400 6140
rect 13832 6140 14964 6168
rect 13832 6100 13860 6140
rect 13372 6072 13860 6100
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 14056 6072 14197 6100
rect 14056 6060 14062 6072
rect 14185 6069 14197 6072
rect 14231 6100 14243 6103
rect 14458 6100 14464 6112
rect 14231 6072 14464 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14826 6100 14832 6112
rect 14787 6072 14832 6100
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 14936 6100 14964 6140
rect 15197 6137 15209 6171
rect 15243 6168 15255 6171
rect 18138 6168 18144 6180
rect 15243 6140 18144 6168
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 16114 6100 16120 6112
rect 14936 6072 16120 6100
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16482 6100 16488 6112
rect 16255 6072 16488 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 16850 6100 16856 6112
rect 16811 6072 16856 6100
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 17221 6103 17279 6109
rect 17221 6069 17233 6103
rect 17267 6100 17279 6103
rect 17586 6100 17592 6112
rect 17267 6072 17592 6100
rect 17267 6069 17279 6072
rect 17221 6063 17279 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 17920 6072 18245 6100
rect 17920 6060 17926 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 18233 6063 18291 6069
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 2222 5896 2228 5908
rect 2183 5868 2228 5896
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 5718 5896 5724 5908
rect 5679 5868 5724 5896
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6546 5896 6552 5908
rect 6135 5868 6552 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 7742 5896 7748 5908
rect 7616 5868 7748 5896
rect 7616 5856 7622 5868
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 8260 5868 8401 5896
rect 8260 5856 8266 5868
rect 8389 5865 8401 5868
rect 8435 5865 8447 5899
rect 8389 5859 8447 5865
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8536 5868 9137 5896
rect 8536 5856 8542 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 9272 5868 11069 5896
rect 9272 5856 9278 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11882 5896 11888 5908
rect 11843 5868 11888 5896
rect 11057 5859 11115 5865
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 12943 5868 14780 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 4154 5828 4160 5840
rect 1688 5800 4160 5828
rect 1688 5769 1716 5800
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 4338 5837 4344 5840
rect 4332 5828 4344 5837
rect 4299 5800 4344 5828
rect 4332 5791 4344 5800
rect 4338 5788 4344 5791
rect 4396 5788 4402 5840
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 5902 5828 5908 5840
rect 4856 5800 5908 5828
rect 4856 5788 4862 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 13532 5831 13590 5837
rect 6472 5800 13492 5828
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1762 5720 1768 5772
rect 1820 5760 1826 5772
rect 2593 5763 2651 5769
rect 2593 5760 2605 5763
rect 1820 5732 2605 5760
rect 1820 5720 1826 5732
rect 2593 5729 2605 5732
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 6472 5760 6500 5800
rect 3283 5732 6500 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 7276 5763 7334 5769
rect 6604 5732 6649 5760
rect 6604 5720 6610 5732
rect 7276 5729 7288 5763
rect 7322 5760 7334 5763
rect 7322 5732 8064 5760
rect 7322 5729 7334 5732
rect 7276 5723 7334 5729
rect 2682 5692 2688 5704
rect 2643 5664 2688 5692
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 3418 5692 3424 5704
rect 2915 5664 3424 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 6178 5692 6184 5704
rect 6139 5664 6184 5692
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6454 5692 6460 5704
rect 6411 5664 6460 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6788 5664 7021 5692
rect 6788 5652 6794 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 8036 5624 8064 5732
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8168 5732 8493 5760
rect 8168 5720 8174 5732
rect 8481 5729 8493 5732
rect 8527 5760 8539 5763
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 8527 5732 8585 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8573 5729 8585 5732
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9030 5760 9036 5772
rect 8987 5732 9036 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9950 5769 9956 5772
rect 9933 5763 9956 5769
rect 9933 5760 9945 5763
rect 9416 5732 9945 5760
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 9416 5692 9444 5732
rect 9933 5729 9945 5732
rect 10008 5760 10014 5772
rect 10008 5732 10081 5760
rect 9933 5723 9956 5729
rect 9950 5720 9956 5723
rect 10008 5720 10014 5732
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 10744 5732 12725 5760
rect 10744 5720 10750 5732
rect 12713 5729 12725 5732
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5760 13323 5763
rect 13354 5760 13360 5772
rect 13311 5732 13360 5760
rect 13311 5729 13323 5732
rect 13265 5723 13323 5729
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 13464 5760 13492 5800
rect 13532 5797 13544 5831
rect 13578 5828 13590 5831
rect 13722 5828 13728 5840
rect 13578 5800 13728 5828
rect 13578 5797 13590 5800
rect 13532 5791 13590 5797
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 14752 5828 14780 5868
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 14884 5868 15669 5896
rect 14884 5856 14890 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 16850 5896 16856 5908
rect 15795 5868 16856 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 16206 5828 16212 5840
rect 14752 5800 16212 5828
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 13998 5760 14004 5772
rect 13464 5732 14004 5760
rect 13998 5720 14004 5732
rect 14056 5720 14062 5772
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14292 5732 15117 5760
rect 8260 5664 9444 5692
rect 8260 5652 8266 5664
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 11974 5692 11980 5704
rect 9732 5664 9777 5692
rect 11935 5664 11980 5692
rect 9732 5652 9738 5664
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12158 5692 12164 5704
rect 12119 5664 12164 5692
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 8110 5624 8116 5636
rect 5000 5596 6868 5624
rect 8023 5596 8116 5624
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5556 1915 5559
rect 2866 5556 2872 5568
rect 1903 5528 2872 5556
rect 1903 5525 1915 5528
rect 1857 5519 1915 5525
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 5000 5556 5028 5596
rect 5442 5556 5448 5568
rect 4304 5528 5028 5556
rect 5403 5528 5448 5556
rect 4304 5516 4310 5528
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6052 5528 6745 5556
rect 6052 5516 6058 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6840 5556 6868 5596
rect 8110 5584 8116 5596
rect 8168 5624 8174 5636
rect 8386 5624 8392 5636
rect 8168 5596 8392 5624
rect 8168 5584 8174 5596
rect 8386 5584 8392 5596
rect 8444 5584 8450 5636
rect 8481 5627 8539 5633
rect 8481 5593 8493 5627
rect 8527 5624 8539 5627
rect 9582 5624 9588 5636
rect 8527 5596 9588 5624
rect 8527 5593 8539 5596
rect 8481 5587 8539 5593
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 10686 5584 10692 5636
rect 10744 5624 10750 5636
rect 12434 5624 12440 5636
rect 10744 5596 12440 5624
rect 10744 5584 10750 5596
rect 12434 5584 12440 5596
rect 12492 5624 12498 5636
rect 13170 5624 13176 5636
rect 12492 5596 13176 5624
rect 12492 5584 12498 5596
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 6840 5528 8769 5556
rect 6733 5519 6791 5525
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 11514 5556 11520 5568
rect 11475 5528 11520 5556
rect 8757 5519 8815 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 14292 5556 14320 5732
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 16741 5763 16799 5769
rect 16741 5760 16753 5763
rect 15105 5723 15163 5729
rect 15856 5732 16753 5760
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 15856 5692 15884 5732
rect 16741 5729 16753 5732
rect 16787 5760 16799 5763
rect 17126 5760 17132 5772
rect 16787 5732 17132 5760
rect 16787 5729 16799 5732
rect 16741 5723 16799 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 14976 5664 15884 5692
rect 15933 5695 15991 5701
rect 14976 5652 14982 5664
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16390 5692 16396 5704
rect 15979 5664 16396 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 14660 5624 14688 5652
rect 16500 5624 16528 5655
rect 14660 5596 16528 5624
rect 13596 5528 14320 5556
rect 13596 5516 13602 5528
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14645 5559 14703 5565
rect 14645 5556 14657 5559
rect 14608 5528 14657 5556
rect 14608 5516 14614 5528
rect 14645 5525 14657 5528
rect 14691 5525 14703 5559
rect 14918 5556 14924 5568
rect 14879 5528 14924 5556
rect 14645 5519 14703 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 17865 5559 17923 5565
rect 17865 5556 17877 5559
rect 17828 5528 17877 5556
rect 17828 5516 17834 5528
rect 17865 5525 17877 5528
rect 17911 5525 17923 5559
rect 17865 5519 17923 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3510 5312 3516 5364
rect 3568 5312 3574 5364
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 3752 5324 5856 5352
rect 3752 5312 3758 5324
rect 3528 5284 3556 5312
rect 3344 5256 3556 5284
rect 5828 5284 5856 5324
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6236 5324 6837 5352
rect 6236 5312 6242 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 7653 5355 7711 5361
rect 6825 5315 6883 5321
rect 6932 5324 7604 5352
rect 6932 5284 6960 5324
rect 5828 5256 6960 5284
rect 7576 5284 7604 5324
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 10137 5355 10195 5361
rect 7699 5324 8340 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 8018 5284 8024 5296
rect 7576 5256 8024 5284
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 1452 5188 2329 5216
rect 1452 5176 1458 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 2038 5148 2044 5160
rect 1627 5120 2044 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5080 1915 5083
rect 2130 5080 2136 5092
rect 1903 5052 2136 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 2130 5040 2136 5052
rect 2188 5040 2194 5092
rect 2584 5083 2642 5089
rect 2584 5049 2596 5083
rect 2630 5080 2642 5083
rect 2774 5080 2780 5092
rect 2630 5052 2780 5080
rect 2630 5049 2642 5052
rect 2584 5043 2642 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 3234 5040 3240 5092
rect 3292 5080 3298 5092
rect 3344 5080 3372 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 4338 5216 4344 5228
rect 3568 5188 4344 5216
rect 3568 5176 3574 5188
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4488 5188 4905 5216
rect 4488 5176 4494 5188
rect 4893 5185 4905 5188
rect 4939 5185 4951 5219
rect 7374 5216 7380 5228
rect 7335 5188 7380 5216
rect 4893 5179 4951 5185
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4798 5148 4804 5160
rect 4203 5120 4804 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 4430 5080 4436 5092
rect 3292 5052 3372 5080
rect 4391 5052 4436 5080
rect 3292 5040 3298 5052
rect 4430 5040 4436 5052
rect 4488 5040 4494 5092
rect 4908 5080 4936 5179
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 8312 5225 8340 5324
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 11882 5352 11888 5364
rect 10183 5324 11888 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 13722 5352 13728 5364
rect 13096 5324 13728 5352
rect 8941 5287 8999 5293
rect 8941 5253 8953 5287
rect 8987 5284 8999 5287
rect 10410 5284 10416 5296
rect 8987 5256 10416 5284
rect 8987 5253 8999 5256
rect 8941 5247 8999 5253
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 12526 5284 12532 5296
rect 10520 5256 12532 5284
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 9490 5216 9496 5228
rect 8444 5188 8489 5216
rect 9451 5188 9496 5216
rect 8444 5176 8450 5188
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 5160 5151 5218 5157
rect 5160 5117 5172 5151
rect 5206 5148 5218 5151
rect 5442 5148 5448 5160
rect 5206 5120 5448 5148
rect 5206 5117 5218 5120
rect 5160 5111 5218 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 6144 5120 7665 5148
rect 6144 5108 6150 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 10520 5157 10548 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11330 5216 11336 5228
rect 10827 5188 11336 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 13096 5216 13124 5324
rect 13722 5312 13728 5324
rect 13780 5352 13786 5364
rect 14461 5355 14519 5361
rect 14461 5352 14473 5355
rect 13780 5324 14473 5352
rect 13780 5312 13786 5324
rect 14461 5321 14473 5324
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14737 5355 14795 5361
rect 14737 5352 14749 5355
rect 14700 5324 14749 5352
rect 14700 5312 14706 5324
rect 14737 5321 14749 5324
rect 14783 5321 14795 5355
rect 14737 5315 14795 5321
rect 11839 5188 13124 5216
rect 14752 5216 14780 5315
rect 15010 5312 15016 5364
rect 15068 5352 15074 5364
rect 17310 5352 17316 5364
rect 15068 5324 17316 5352
rect 15068 5312 15074 5324
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 14752 5188 15025 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 15013 5185 15025 5188
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17184 5188 17509 5216
rect 17184 5176 17190 5188
rect 17497 5185 17509 5188
rect 17543 5216 17555 5219
rect 17586 5216 17592 5228
rect 17543 5188 17592 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 7984 5120 9413 5148
rect 7984 5108 7990 5120
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5117 10563 5151
rect 10962 5148 10968 5160
rect 10505 5111 10563 5117
rect 10612 5120 10968 5148
rect 5258 5080 5264 5092
rect 4908 5052 5264 5080
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 5810 5040 5816 5092
rect 5868 5080 5874 5092
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 5868 5052 9321 5080
rect 5868 5040 5874 5052
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9309 5043 9367 5049
rect 9674 5040 9680 5092
rect 9732 5080 9738 5092
rect 10612 5089 10640 5120
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11514 5148 11520 5160
rect 11475 5120 11520 5148
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12492 5120 13093 5148
rect 12492 5108 12498 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 14918 5148 14924 5160
rect 14879 5120 14924 5148
rect 13081 5111 13139 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15280 5151 15338 5157
rect 15280 5117 15292 5151
rect 15326 5148 15338 5151
rect 17770 5148 17776 5160
rect 15326 5120 17776 5148
rect 15326 5117 15338 5120
rect 15280 5111 15338 5117
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 10597 5083 10655 5089
rect 10597 5080 10609 5083
rect 9732 5052 10609 5080
rect 9732 5040 9738 5052
rect 10597 5049 10609 5052
rect 10643 5049 10655 5083
rect 11238 5080 11244 5092
rect 10597 5043 10655 5049
rect 10980 5052 11244 5080
rect 1946 4972 1952 5024
rect 2004 5012 2010 5024
rect 2222 5012 2228 5024
rect 2004 4984 2228 5012
rect 2004 4972 2010 4984
rect 2222 4972 2228 4984
rect 2280 5012 2286 5024
rect 3697 5015 3755 5021
rect 3697 5012 3709 5015
rect 2280 4984 3709 5012
rect 2280 4972 2286 4984
rect 3697 4981 3709 4984
rect 3743 4981 3755 5015
rect 3697 4975 3755 4981
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 5534 5012 5540 5024
rect 4396 4984 5540 5012
rect 4396 4972 4402 4984
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6512 4984 7205 5012
rect 6512 4972 6518 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7331 4984 7849 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 7837 4975 7895 4981
rect 8205 5015 8263 5021
rect 8205 4981 8217 5015
rect 8251 5012 8263 5015
rect 8478 5012 8484 5024
rect 8251 4984 8484 5012
rect 8251 4981 8263 4984
rect 8205 4975 8263 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 10980 5012 11008 5052
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 12158 5040 12164 5092
rect 12216 5080 12222 5092
rect 13348 5083 13406 5089
rect 13348 5080 13360 5083
rect 12216 5052 13360 5080
rect 12216 5040 12222 5052
rect 13348 5049 13360 5052
rect 13394 5080 13406 5083
rect 13998 5080 14004 5092
rect 13394 5052 14004 5080
rect 13394 5049 13406 5052
rect 13348 5043 13406 5049
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 17034 5040 17040 5092
rect 17092 5080 17098 5092
rect 18064 5080 18092 5111
rect 17092 5052 18092 5080
rect 17092 5040 17098 5052
rect 11146 5012 11152 5024
rect 8812 4984 11008 5012
rect 11107 4984 11152 5012
rect 8812 4972 8818 4984
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 11572 4984 11621 5012
rect 11572 4972 11578 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 11609 4975 11667 4981
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 11756 4984 12449 5012
rect 11756 4972 11762 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12437 4975 12495 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 14366 5012 14372 5024
rect 12584 4984 14372 5012
rect 12584 4972 12590 4984
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16942 5012 16948 5024
rect 16903 4984 16948 5012
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 18233 5015 18291 5021
rect 17460 4984 17505 5012
rect 17460 4972 17466 4984
rect 18233 4981 18245 5015
rect 18279 5012 18291 5015
rect 18322 5012 18328 5024
rect 18279 4984 18328 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 18322 4972 18328 4984
rect 18380 4972 18386 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 2590 4768 2596 4820
rect 2648 4808 2654 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2648 4780 2973 4808
rect 2648 4768 2654 4780
rect 2961 4777 2973 4780
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 3326 4768 3332 4820
rect 3384 4768 3390 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 4571 4780 5089 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 5077 4771 5135 4777
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 5316 4780 6101 4808
rect 5316 4768 5322 4780
rect 6089 4777 6101 4780
rect 6135 4777 6147 4811
rect 6089 4771 6147 4777
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 8754 4808 8760 4820
rect 6512 4780 8760 4808
rect 6512 4768 6518 4780
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9030 4808 9036 4820
rect 8991 4780 9036 4808
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9861 4811 9919 4817
rect 9861 4777 9873 4811
rect 9907 4777 9919 4811
rect 9861 4771 9919 4777
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 10183 4780 10977 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 10965 4771 11023 4777
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 3344 4740 3372 4768
rect 4246 4740 4252 4752
rect 2455 4712 3372 4740
rect 3436 4712 4252 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1486 4672 1492 4684
rect 1443 4644 1492 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2424 4644 3188 4672
rect 1210 4564 1216 4616
rect 1268 4604 1274 4616
rect 2424 4604 2452 4644
rect 1268 4576 2452 4604
rect 1268 4564 1274 4576
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 3160 4604 3188 4644
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 3292 4644 3341 4672
rect 3292 4632 3298 4644
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3436 4613 3464 4712
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 5810 4700 5816 4752
rect 5868 4740 5874 4752
rect 9876 4740 9904 4771
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 15102 4808 15108 4820
rect 14424 4780 15108 4808
rect 14424 4768 14430 4780
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 16482 4768 16488 4820
rect 16540 4808 16546 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16540 4780 16681 4808
rect 16540 4768 16546 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 16669 4771 16727 4777
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 17678 4808 17684 4820
rect 17543 4780 17684 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 5868 4712 9904 4740
rect 5868 4700 5874 4712
rect 10318 4700 10324 4752
rect 10376 4700 10382 4752
rect 11885 4743 11943 4749
rect 11885 4740 11897 4743
rect 10704 4712 11897 4740
rect 4338 4672 4344 4684
rect 3528 4644 4344 4672
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 2556 4576 2601 4604
rect 3160 4576 3433 4604
rect 2556 4564 2562 4576
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 1949 4539 2007 4545
rect 1949 4505 1961 4539
rect 1995 4536 2007 4539
rect 3528 4536 3556 4644
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 5718 4672 5724 4684
rect 5491 4644 5724 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 3786 4604 3792 4616
rect 3651 4576 3792 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 1995 4508 3556 4536
rect 1995 4505 2007 4508
rect 1949 4499 2007 4505
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2498 4428 2504 4480
rect 2556 4468 2562 4480
rect 3620 4468 3648 4567
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4448 4604 4476 4635
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6273 4675 6331 4681
rect 6273 4672 6285 4675
rect 5960 4644 6285 4672
rect 5960 4632 5966 4644
rect 6273 4641 6285 4644
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6621 4675 6679 4681
rect 6621 4672 6633 4675
rect 6512 4644 6633 4672
rect 6512 4632 6518 4644
rect 6621 4641 6633 4644
rect 6667 4641 6679 4675
rect 6621 4635 6679 4641
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7432 4644 8033 4672
rect 7432 4632 7438 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8938 4672 8944 4684
rect 8899 4644 8944 4672
rect 8021 4635 8079 4641
rect 4614 4604 4620 4616
rect 4212 4576 4476 4604
rect 4575 4576 4620 4604
rect 4212 4564 4218 4576
rect 4448 4536 4476 4576
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 5629 4567 5687 4573
rect 6288 4576 6377 4604
rect 4798 4536 4804 4548
rect 4448 4508 4804 4536
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 5644 4536 5672 4567
rect 5500 4508 5672 4536
rect 5500 4496 5506 4508
rect 2556 4440 3648 4468
rect 4065 4471 4123 4477
rect 2556 4428 2562 4440
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 5074 4468 5080 4480
rect 4111 4440 5080 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 6288 4468 6316 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 7926 4604 7932 4616
rect 6365 4567 6423 4573
rect 7760 4576 7932 4604
rect 7760 4545 7788 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 7745 4539 7803 4545
rect 7745 4505 7757 4539
rect 7791 4505 7803 4539
rect 8036 4536 8064 4635
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4672 9735 4675
rect 10336 4672 10364 4700
rect 9723 4644 10364 4672
rect 10413 4675 10471 4681
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 10413 4641 10425 4675
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9306 4604 9312 4616
rect 9263 4576 9312 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9416 4576 10149 4604
rect 8294 4536 8300 4548
rect 8036 4508 8300 4536
rect 7745 4499 7803 4505
rect 8294 4496 8300 4508
rect 8352 4536 8358 4548
rect 9416 4536 9444 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 8352 4508 9444 4536
rect 8352 4496 8358 4508
rect 9582 4496 9588 4548
rect 9640 4536 9646 4548
rect 10042 4536 10048 4548
rect 9640 4508 10048 4536
rect 9640 4496 9646 4508
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 6730 4468 6736 4480
rect 5592 4440 6736 4468
rect 5592 4428 5598 4440
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 8076 4440 8217 4468
rect 8076 4428 8082 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 9674 4468 9680 4480
rect 8619 4440 9680 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10229 4471 10287 4477
rect 10229 4468 10241 4471
rect 9824 4440 10241 4468
rect 9824 4428 9830 4440
rect 10229 4437 10241 4440
rect 10275 4468 10287 4471
rect 10318 4468 10324 4480
rect 10275 4440 10324 4468
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 10428 4468 10456 4635
rect 10505 4539 10563 4545
rect 10505 4505 10517 4539
rect 10551 4536 10563 4539
rect 10704 4536 10732 4712
rect 11885 4709 11897 4712
rect 11931 4709 11943 4743
rect 11885 4703 11943 4709
rect 13170 4700 13176 4752
rect 13228 4740 13234 4752
rect 17405 4743 17463 4749
rect 17405 4740 17417 4743
rect 13228 4712 17417 4740
rect 13228 4700 13234 4712
rect 17405 4709 17417 4712
rect 17451 4709 17463 4743
rect 17405 4703 17463 4709
rect 10870 4672 10876 4684
rect 10783 4644 10876 4672
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11330 4672 11336 4684
rect 11164 4644 11336 4672
rect 10551 4508 10732 4536
rect 10888 4536 10916 4632
rect 11164 4613 11192 4644
rect 11330 4632 11336 4644
rect 11388 4672 11394 4684
rect 12877 4675 12935 4681
rect 12877 4672 12889 4675
rect 11388 4644 12889 4672
rect 11388 4632 11394 4644
rect 12877 4641 12889 4644
rect 12923 4672 12935 4675
rect 13722 4672 13728 4684
rect 12923 4644 13728 4672
rect 12923 4641 12935 4644
rect 12877 4635 12935 4641
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14332 4644 14657 4672
rect 14332 4632 14338 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 16482 4632 16488 4684
rect 16540 4672 16546 4684
rect 16540 4644 16585 4672
rect 16540 4632 16546 4644
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 18049 4675 18107 4681
rect 18049 4672 18061 4675
rect 17552 4644 18061 4672
rect 17552 4632 17558 4644
rect 18049 4641 18061 4644
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11572 4576 11989 4604
rect 11572 4564 11578 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 12158 4604 12164 4616
rect 12119 4576 12164 4604
rect 11977 4567 12035 4573
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12492 4576 12633 4604
rect 12492 4564 12498 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15712 4576 15761 4604
rect 15712 4564 15718 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 15841 4567 15899 4573
rect 11606 4536 11612 4548
rect 10888 4508 11612 4536
rect 10551 4505 10563 4508
rect 10505 4499 10563 4505
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 14829 4539 14887 4545
rect 14829 4505 14841 4539
rect 14875 4536 14887 4539
rect 15378 4536 15384 4548
rect 14875 4508 15384 4536
rect 14875 4505 14887 4508
rect 14829 4499 14887 4505
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 15562 4496 15568 4548
rect 15620 4536 15626 4548
rect 15856 4536 15884 4567
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 15620 4508 15884 4536
rect 15620 4496 15626 4508
rect 14918 4468 14924 4480
rect 10428 4440 14924 4468
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 17034 4468 17040 4480
rect 16995 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 18230 4468 18236 4480
rect 18191 4440 18236 4468
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 2832 4236 2877 4264
rect 2832 4224 2838 4236
rect 6638 4224 6644 4276
rect 6696 4264 6702 4276
rect 8018 4264 8024 4276
rect 6696 4236 8024 4264
rect 6696 4224 6702 4236
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8570 4224 8576 4276
rect 8628 4264 8634 4276
rect 9766 4264 9772 4276
rect 8628 4236 9772 4264
rect 8628 4224 8634 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10520 4236 11560 4264
rect 6288 4168 7420 4196
rect 6288 4140 6316 4168
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3068 4100 3985 4128
rect 1412 4060 1440 4088
rect 3068 4060 3096 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 3973 4091 4031 4097
rect 5920 4100 6193 4128
rect 3234 4060 3240 4072
rect 1412 4032 3096 4060
rect 3195 4032 3240 4060
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 5810 4060 5816 4072
rect 3559 4032 5816 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 382 3952 388 4004
rect 440 3992 446 4004
rect 1642 3995 1700 4001
rect 1642 3992 1654 3995
rect 440 3964 1654 3992
rect 440 3952 446 3964
rect 1642 3961 1654 3964
rect 1688 3961 1700 3995
rect 1642 3955 1700 3961
rect 4240 3995 4298 4001
rect 4240 3961 4252 3995
rect 4286 3992 4298 3995
rect 4614 3992 4620 4004
rect 4286 3964 4620 3992
rect 4286 3961 4298 3964
rect 4240 3955 4298 3961
rect 4614 3952 4620 3964
rect 4672 3992 4678 4004
rect 5920 3992 5948 4100
rect 6181 4097 6193 4100
rect 6227 4128 6239 4131
rect 6270 4128 6276 4140
rect 6227 4100 6276 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 7392 4137 7420 4168
rect 7377 4131 7435 4137
rect 6696 4100 7144 4128
rect 6696 4088 6702 4100
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 7006 4060 7012 4072
rect 6135 4032 7012 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7116 4060 7144 4100
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10520 4137 10548 4236
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10376 4100 10517 4128
rect 10376 4088 10382 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 11532 4128 11560 4236
rect 13722 4224 13728 4276
rect 13780 4264 13786 4276
rect 13817 4267 13875 4273
rect 13817 4264 13829 4267
rect 13780 4236 13829 4264
rect 13780 4224 13786 4236
rect 13817 4233 13829 4236
rect 13863 4233 13875 4267
rect 14642 4264 14648 4276
rect 13817 4227 13875 4233
rect 14292 4236 14648 4264
rect 12434 4128 12440 4140
rect 11532 4100 12440 4128
rect 10505 4091 10563 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 14292 4137 14320 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15654 4224 15660 4276
rect 15712 4264 15718 4276
rect 15933 4267 15991 4273
rect 15933 4264 15945 4267
rect 15712 4236 15945 4264
rect 15712 4224 15718 4236
rect 15933 4233 15945 4236
rect 15979 4233 15991 4267
rect 15933 4227 15991 4233
rect 17770 4196 17776 4208
rect 17604 4168 17776 4196
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4097 16543 4131
rect 16485 4091 16543 4097
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7116 4032 7297 4060
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 8294 4060 8300 4072
rect 7883 4032 8300 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8444 4032 8489 4060
rect 8444 4020 8450 4032
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 14544 4063 14602 4069
rect 9272 4032 14504 4060
rect 9272 4020 9278 4032
rect 4672 3964 5948 3992
rect 5997 3995 6055 4001
rect 4672 3952 4678 3964
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6546 3992 6552 4004
rect 6043 3964 6552 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 8656 3995 8714 4001
rect 6696 3964 8064 3992
rect 6696 3952 6702 3964
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4430 3924 4436 3936
rect 3844 3896 4436 3924
rect 3844 3884 3850 3896
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 5316 3896 5365 3924
rect 5316 3884 5322 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5626 3924 5632 3936
rect 5587 3896 5632 3924
rect 5353 3887 5411 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 6178 3884 6184 3936
rect 6236 3924 6242 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6236 3896 6837 3924
rect 6236 3884 6242 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 6825 3887 6883 3893
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7558 3924 7564 3936
rect 7239 3896 7564 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 8036 3933 8064 3964
rect 8656 3961 8668 3995
rect 8702 3992 8714 3995
rect 9306 3992 9312 4004
rect 8702 3964 9312 3992
rect 8702 3961 8714 3964
rect 8656 3955 8714 3961
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 10134 3992 10140 4004
rect 9784 3964 10140 3992
rect 9784 3933 9812 3964
rect 10134 3952 10140 3964
rect 10192 3992 10198 4004
rect 12710 4001 12716 4004
rect 10750 3995 10808 4001
rect 10750 3992 10762 3995
rect 10192 3964 10762 3992
rect 10192 3952 10198 3964
rect 10750 3961 10762 3964
rect 10796 3961 10808 3995
rect 12704 3992 12716 4001
rect 10750 3955 10808 3961
rect 11900 3964 12716 3992
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3893 9827 3927
rect 9769 3887 9827 3893
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10962 3924 10968 3936
rect 10091 3896 10968 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11900 3933 11928 3964
rect 12704 3955 12716 3964
rect 12710 3952 12716 3955
rect 12768 3952 12774 4004
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 14366 3924 14372 3936
rect 12216 3896 14372 3924
rect 12216 3884 12222 3896
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14476 3924 14504 4032
rect 14544 4029 14556 4063
rect 14590 4060 14602 4063
rect 16390 4060 16396 4072
rect 14590 4032 16396 4060
rect 14590 4029 14602 4032
rect 14544 4023 14602 4029
rect 16390 4020 16396 4032
rect 16448 4060 16454 4072
rect 16500 4060 16528 4091
rect 16942 4088 16948 4140
rect 17000 4128 17006 4140
rect 17604 4137 17632 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 17000 4100 17417 4128
rect 17000 4088 17006 4100
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 17589 4131 17647 4137
rect 17589 4097 17601 4131
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 16448 4032 16528 4060
rect 16448 4020 16454 4032
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 17092 4032 17325 4060
rect 17092 4020 17098 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17552 4032 18061 4060
rect 17552 4020 17558 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 16298 3992 16304 4004
rect 16259 3964 16304 3992
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 16758 3952 16764 4004
rect 16816 3992 16822 4004
rect 17586 3992 17592 4004
rect 16816 3964 17592 3992
rect 16816 3952 16822 3964
rect 17586 3952 17592 3964
rect 17644 3952 17650 4004
rect 15562 3924 15568 3936
rect 14476 3896 15568 3924
rect 15562 3884 15568 3896
rect 15620 3924 15626 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15620 3896 15669 3924
rect 15620 3884 15626 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16439 3896 16957 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 16945 3887 17003 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 1394 3680 1400 3732
rect 1452 3680 1458 3732
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2314 3720 2320 3732
rect 2179 3692 2320 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2464 3692 3188 3720
rect 2464 3680 2470 3692
rect 1412 3652 1440 3680
rect 1673 3655 1731 3661
rect 1412 3624 1624 3652
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1412 3380 1440 3547
rect 1596 3516 1624 3624
rect 1673 3621 1685 3655
rect 1719 3652 1731 3655
rect 3050 3652 3056 3664
rect 1719 3624 3056 3652
rect 1719 3621 1731 3624
rect 1673 3615 1731 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 2406 3544 2412 3596
rect 2464 3584 2470 3596
rect 3160 3593 3188 3692
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 4522 3720 4528 3732
rect 3292 3692 4528 3720
rect 3292 3680 3298 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 4985 3723 5043 3729
rect 4985 3689 4997 3723
rect 5031 3720 5043 3723
rect 5626 3720 5632 3732
rect 5031 3692 5632 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 6788 3692 7389 3720
rect 6788 3680 6794 3692
rect 7377 3689 7389 3692
rect 7423 3720 7435 3723
rect 8386 3720 8392 3732
rect 7423 3692 8392 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 5074 3652 5080 3664
rect 3752 3624 4200 3652
rect 5035 3624 5080 3652
rect 3752 3612 3758 3624
rect 2501 3587 2559 3593
rect 2501 3584 2513 3587
rect 2464 3556 2513 3584
rect 2464 3544 2470 3556
rect 2501 3553 2513 3556
rect 2547 3553 2559 3587
rect 2501 3547 2559 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3553 3203 3587
rect 4062 3584 4068 3596
rect 4023 3556 4068 3584
rect 3145 3547 3203 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4172 3584 4200 3624
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 5184 3624 6776 3652
rect 5184 3584 5212 3624
rect 5977 3587 6035 3593
rect 5977 3584 5989 3587
rect 4172 3556 5212 3584
rect 5276 3556 5989 3584
rect 5276 3528 5304 3556
rect 5977 3553 5989 3556
rect 6023 3553 6035 3587
rect 5977 3547 6035 3553
rect 2590 3516 2596 3528
rect 1596 3488 2596 3516
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 4890 3516 4896 3528
rect 3467 3488 4896 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 2700 3448 2728 3479
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5258 3516 5264 3528
rect 5219 3488 5264 3516
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5592 3488 5733 3516
rect 5592 3476 5598 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 6748 3516 6776 3624
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7668 3593 7696 3692
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 9732 3692 10149 3720
rect 9732 3680 9738 3692
rect 10137 3689 10149 3692
rect 10183 3689 10195 3723
rect 10137 3683 10195 3689
rect 10965 3723 11023 3729
rect 10965 3689 10977 3723
rect 11011 3720 11023 3723
rect 11514 3720 11520 3732
rect 11011 3692 11520 3720
rect 11011 3689 11023 3692
rect 10965 3683 11023 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 11974 3720 11980 3732
rect 11935 3692 11980 3720
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 12308 3692 12357 3720
rect 12308 3680 12314 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12345 3683 12403 3689
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 12526 3720 12532 3732
rect 12483 3692 12532 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13906 3720 13912 3732
rect 13867 3692 13912 3720
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 14458 3720 14464 3732
rect 14415 3692 14464 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 17402 3720 17408 3732
rect 17276 3692 17408 3720
rect 17276 3680 17282 3692
rect 17402 3680 17408 3692
rect 17460 3720 17466 3732
rect 17460 3692 17816 3720
rect 17460 3680 17466 3692
rect 7920 3655 7978 3661
rect 7920 3621 7932 3655
rect 7966 3652 7978 3655
rect 9122 3652 9128 3664
rect 7966 3624 9128 3652
rect 7966 3621 7978 3624
rect 7920 3615 7978 3621
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 10594 3652 10600 3664
rect 9232 3624 10600 3652
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7524 3556 7573 3584
rect 7524 3544 7530 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 7653 3587 7711 3593
rect 7653 3553 7665 3587
rect 7699 3553 7711 3587
rect 9232 3584 9260 3624
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 14277 3655 14335 3661
rect 14277 3621 14289 3655
rect 14323 3652 14335 3655
rect 15010 3652 15016 3664
rect 14323 3624 15016 3652
rect 14323 3621 14335 3624
rect 14277 3615 14335 3621
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 15120 3624 16344 3652
rect 7653 3547 7711 3553
rect 7760 3556 9260 3584
rect 7760 3516 7788 3556
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9640 3556 10057 3584
rect 9640 3544 9646 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 11330 3584 11336 3596
rect 10192 3556 10272 3584
rect 11291 3556 11336 3584
rect 10192 3544 10198 3556
rect 10244 3525 10272 3556
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 12989 3587 13047 3593
rect 12989 3584 13001 3587
rect 12676 3556 13001 3584
rect 12676 3544 12682 3556
rect 12989 3553 13001 3556
rect 13035 3553 13047 3587
rect 12989 3547 13047 3553
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 15120 3584 15148 3624
rect 16316 3596 16344 3624
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 17313 3655 17371 3661
rect 17313 3652 17325 3655
rect 16540 3624 17325 3652
rect 16540 3612 16546 3624
rect 17313 3621 17325 3624
rect 17359 3621 17371 3655
rect 17313 3615 17371 3621
rect 15286 3584 15292 3596
rect 14424 3556 15148 3584
rect 15247 3556 15292 3584
rect 14424 3544 14430 3556
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 16298 3584 16304 3596
rect 16259 3556 16304 3584
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 17034 3584 17040 3596
rect 16995 3556 17040 3584
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 17788 3593 17816 3692
rect 17773 3587 17831 3593
rect 17773 3553 17785 3587
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 6748 3488 7788 3516
rect 10229 3519 10287 3525
rect 5721 3479 5779 3485
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 11238 3516 11244 3528
rect 10468 3488 11244 3516
rect 10468 3476 10474 3488
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11422 3516 11428 3528
rect 11383 3488 11428 3516
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 11572 3488 12541 3516
rect 11572 3476 11578 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 12529 3479 12587 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 14550 3516 14556 3528
rect 14511 3488 14556 3516
rect 14550 3476 14556 3488
rect 14608 3476 14614 3528
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3516 15623 3519
rect 15654 3516 15660 3528
rect 15611 3488 15660 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3485 16635 3519
rect 18046 3516 18052 3528
rect 18007 3488 18052 3516
rect 16577 3479 16635 3485
rect 2556 3420 2728 3448
rect 2556 3408 2562 3420
rect 3510 3408 3516 3460
rect 3568 3448 3574 3460
rect 4249 3451 4307 3457
rect 4249 3448 4261 3451
rect 3568 3420 4261 3448
rect 3568 3408 3574 3420
rect 4249 3417 4261 3420
rect 4295 3417 4307 3451
rect 11698 3448 11704 3460
rect 4249 3411 4307 3417
rect 8588 3420 11704 3448
rect 4338 3380 4344 3392
rect 1412 3352 4344 3380
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4614 3380 4620 3392
rect 4575 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 6454 3380 6460 3392
rect 5592 3352 6460 3380
rect 5592 3340 5598 3352
rect 6454 3340 6460 3352
rect 6512 3380 6518 3392
rect 7101 3383 7159 3389
rect 7101 3380 7113 3383
rect 6512 3352 7113 3380
rect 6512 3340 6518 3352
rect 7101 3349 7113 3352
rect 7147 3349 7159 3383
rect 7101 3343 7159 3349
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 8588 3380 8616 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 16592 3448 16620 3479
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18506 3448 18512 3460
rect 16592 3420 18512 3448
rect 18506 3408 18512 3420
rect 18564 3408 18570 3460
rect 7248 3352 8616 3380
rect 9033 3383 9091 3389
rect 7248 3340 7254 3352
rect 9033 3349 9045 3383
rect 9079 3380 9091 3383
rect 9306 3380 9312 3392
rect 9079 3352 9312 3380
rect 9079 3349 9091 3352
rect 9033 3343 9091 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 11054 3380 11060 3392
rect 9723 3352 11060 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 17310 3380 17316 3392
rect 11664 3352 17316 3380
rect 11664 3340 11670 3352
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 2682 3176 2688 3188
rect 1719 3148 2688 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 3513 3179 3571 3185
rect 3513 3145 3525 3179
rect 3559 3176 3571 3179
rect 6086 3176 6092 3188
rect 3559 3148 6092 3176
rect 3559 3145 3571 3148
rect 3513 3139 3571 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 7190 3176 7196 3188
rect 6595 3148 7196 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 8573 3179 8631 3185
rect 8573 3145 8585 3179
rect 8619 3176 8631 3179
rect 8938 3176 8944 3188
rect 8619 3148 8944 3176
rect 8619 3145 8631 3148
rect 8573 3139 8631 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9582 3176 9588 3188
rect 9543 3148 9588 3176
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10502 3176 10508 3188
rect 9824 3148 10508 3176
rect 9824 3136 9830 3148
rect 10502 3136 10508 3148
rect 10560 3176 10566 3188
rect 10560 3148 10824 3176
rect 10560 3136 10566 3148
rect 3605 3111 3663 3117
rect 3605 3077 3617 3111
rect 3651 3108 3663 3111
rect 4982 3108 4988 3120
rect 3651 3080 4988 3108
rect 3651 3077 3663 3080
rect 3605 3071 3663 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 7374 3108 7380 3120
rect 5500 3080 7380 3108
rect 5500 3068 5506 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 7561 3111 7619 3117
rect 7561 3077 7573 3111
rect 7607 3108 7619 3111
rect 8754 3108 8760 3120
rect 7607 3080 8760 3108
rect 7607 3077 7619 3080
rect 7561 3071 7619 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 10686 3108 10692 3120
rect 9048 3080 10692 3108
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3234 3040 3240 3052
rect 2832 3012 3240 3040
rect 2832 3000 2838 3012
rect 3234 3000 3240 3012
rect 3292 3040 3298 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 3292 3012 4261 3040
rect 3292 3000 3298 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 5258 3040 5264 3052
rect 5219 3012 5264 3040
rect 4249 3003 4307 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 6178 3040 6184 3052
rect 5644 3012 6184 3040
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3384 2944 4077 2972
rect 3384 2932 3390 2944
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5644 2972 5672 3012
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6328 3012 6373 3040
rect 6328 3000 6334 3012
rect 6546 3000 6552 3052
rect 6604 3040 6610 3052
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6604 3012 7481 3040
rect 6604 3000 6610 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7800 3012 8033 3040
rect 7800 3000 7806 3012
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8202 3040 8208 3052
rect 8163 3012 8208 3040
rect 8021 3003 8079 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 9048 3049 9076 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 10796 3108 10824 3148
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 11480 3148 12449 3176
rect 11480 3136 11486 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 13449 3179 13507 3185
rect 13449 3145 13461 3179
rect 13495 3176 13507 3179
rect 13630 3176 13636 3188
rect 13495 3148 13636 3176
rect 13495 3145 13507 3148
rect 13449 3139 13507 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18414 3176 18420 3188
rect 18279 3148 18420 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 10796 3080 11744 3108
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8352 3012 9045 3040
rect 8352 3000 8358 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9180 3012 9225 3040
rect 9180 3000 9186 3012
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 10137 3043 10195 3049
rect 10137 3040 10149 3043
rect 9364 3012 10149 3040
rect 9364 3000 9370 3012
rect 10137 3009 10149 3012
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 10928 3012 11069 3040
rect 10928 3000 10934 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 11238 3040 11244 3052
rect 11199 3012 11244 3040
rect 11057 3003 11115 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 5215 2944 5672 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6512 2944 6837 2972
rect 6512 2932 6518 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 7926 2972 7932 2984
rect 7887 2944 7932 2972
rect 6825 2935 6883 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 2406 2864 2412 2916
rect 2464 2904 2470 2916
rect 2774 2904 2780 2916
rect 2464 2876 2780 2904
rect 2464 2864 2470 2876
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 3145 2907 3203 2913
rect 3145 2873 3157 2907
rect 3191 2904 3203 2907
rect 3513 2907 3571 2913
rect 3513 2904 3525 2907
rect 3191 2876 3525 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 3513 2873 3525 2876
rect 3559 2873 3571 2907
rect 3513 2867 3571 2873
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 4246 2904 4252 2916
rect 4203 2876 4252 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 6086 2904 6092 2916
rect 5123 2876 5672 2904
rect 6047 2876 6092 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 2133 2839 2191 2845
rect 2133 2805 2145 2839
rect 2179 2836 2191 2839
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2179 2808 2697 2836
rect 2179 2805 2191 2808
rect 2133 2799 2191 2805
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 3099 2808 3617 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3605 2805 3617 2808
rect 3651 2805 3663 2839
rect 3605 2799 3663 2805
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 4706 2836 4712 2848
rect 3752 2808 3797 2836
rect 4667 2808 4712 2836
rect 3752 2796 3758 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 5644 2836 5672 2876
rect 6086 2864 6092 2876
rect 6144 2864 6150 2916
rect 6270 2864 6276 2916
rect 6328 2904 6334 2916
rect 6549 2907 6607 2913
rect 6549 2904 6561 2907
rect 6328 2876 6561 2904
rect 6328 2864 6334 2876
rect 6549 2873 6561 2876
rect 6595 2873 6607 2907
rect 6549 2867 6607 2873
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 7101 2907 7159 2913
rect 7101 2904 7113 2907
rect 6788 2876 7113 2904
rect 6788 2864 6794 2876
rect 7101 2873 7113 2876
rect 7147 2873 7159 2907
rect 7101 2867 7159 2873
rect 7469 2907 7527 2913
rect 7469 2873 7481 2907
rect 7515 2904 7527 2907
rect 8941 2907 8999 2913
rect 8941 2904 8953 2907
rect 7515 2876 8953 2904
rect 7515 2873 7527 2876
rect 7469 2867 7527 2873
rect 8941 2873 8953 2876
rect 8987 2873 8999 2907
rect 9140 2904 9168 3000
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 10962 2972 10968 2984
rect 9456 2944 10732 2972
rect 10923 2944 10968 2972
rect 9456 2932 9462 2944
rect 9490 2904 9496 2916
rect 9140 2876 9496 2904
rect 8941 2867 8999 2873
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 9953 2907 10011 2913
rect 9953 2873 9965 2907
rect 9999 2904 10011 2907
rect 10704 2904 10732 2944
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 11388 2944 11621 2972
rect 11388 2932 11394 2944
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11716 2972 11744 3080
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 12124 3080 13840 3108
rect 12124 3068 12130 3080
rect 12710 3000 12716 3052
rect 12768 3040 12774 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12768 3012 13001 3040
rect 12768 3000 12774 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 13812 3040 13840 3080
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 13964 3080 14688 3108
rect 13964 3068 13970 3080
rect 14660 3049 14688 3080
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13812 3012 14013 3040
rect 12989 3003 13047 3009
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 15470 3040 15476 3052
rect 14645 3003 14703 3009
rect 14936 3012 15476 3040
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 11716 2944 12817 2972
rect 11609 2935 11667 2941
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 13814 2972 13820 2984
rect 13775 2944 13820 2972
rect 12805 2935 12863 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 14936 2972 14964 3012
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 17402 3040 17408 3052
rect 17236 3012 17408 3040
rect 15194 2972 15200 2984
rect 14507 2944 14964 2972
rect 15155 2944 15200 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 16172 2944 16497 2972
rect 16172 2932 16178 2944
rect 16485 2941 16497 2944
rect 16531 2972 16543 2975
rect 16574 2972 16580 2984
rect 16531 2944 16580 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 17236 2981 17264 3012
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 19426 3040 19432 3052
rect 17543 3012 19432 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17368 2944 18061 2972
rect 17368 2932 17374 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 9999 2876 10640 2904
rect 10704 2876 11897 2904
rect 9999 2873 10011 2876
rect 9953 2867 10011 2873
rect 5721 2839 5779 2845
rect 5721 2836 5733 2839
rect 5644 2808 5733 2836
rect 5721 2805 5733 2808
rect 5767 2805 5779 2839
rect 5721 2799 5779 2805
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6362 2836 6368 2848
rect 6227 2808 6368 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 9858 2836 9864 2848
rect 8076 2808 9864 2836
rect 8076 2796 8082 2808
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10612 2845 10640 2876
rect 11885 2873 11897 2876
rect 11931 2873 11943 2907
rect 11885 2867 11943 2873
rect 13909 2907 13967 2913
rect 13909 2873 13921 2907
rect 13955 2904 13967 2907
rect 14090 2904 14096 2916
rect 13955 2876 14096 2904
rect 13955 2873 13967 2876
rect 13909 2867 13967 2873
rect 14090 2864 14096 2876
rect 14148 2864 14154 2916
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 14884 2876 15485 2904
rect 14884 2864 14890 2876
rect 15473 2873 15485 2876
rect 15519 2873 15531 2907
rect 16758 2904 16764 2916
rect 16719 2876 16764 2904
rect 15473 2867 15531 2873
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 10597 2839 10655 2845
rect 10100 2808 10145 2836
rect 10100 2796 10106 2808
rect 10597 2805 10609 2839
rect 10643 2805 10655 2839
rect 10597 2799 10655 2805
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 10836 2808 12909 2836
rect 10836 2796 10842 2808
rect 12897 2805 12909 2808
rect 12943 2836 12955 2839
rect 17494 2836 17500 2848
rect 12943 2808 17500 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1762 2632 1768 2644
rect 1719 2604 1768 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2096 2604 2697 2632
rect 2096 2592 2102 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 2685 2595 2743 2601
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 2832 2604 3065 2632
rect 2832 2592 2838 2604
rect 3053 2601 3065 2604
rect 3099 2632 3111 2635
rect 4249 2635 4307 2641
rect 3099 2604 4200 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 3694 2564 3700 2576
rect 2179 2536 3700 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 4172 2564 4200 2604
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 4338 2632 4344 2644
rect 4295 2604 4344 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4706 2632 4712 2644
rect 4663 2604 4712 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5350 2632 5356 2644
rect 5307 2604 5356 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 5718 2632 5724 2644
rect 5675 2604 5724 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 7834 2632 7840 2644
rect 6380 2604 7840 2632
rect 5442 2564 5448 2576
rect 4172 2536 5448 2564
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 6380 2564 6408 2604
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8754 2592 8760 2644
rect 8812 2632 8818 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8812 2604 9137 2632
rect 8812 2592 8818 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 9125 2595 9183 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10502 2632 10508 2644
rect 10459 2604 10508 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 16577 2635 16635 2641
rect 16577 2632 16589 2635
rect 12492 2604 16589 2632
rect 12492 2592 12498 2604
rect 16577 2601 16589 2604
rect 16623 2632 16635 2635
rect 16850 2632 16856 2644
rect 16623 2604 16856 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 5736 2536 6408 2564
rect 2041 2499 2099 2505
rect 2041 2465 2053 2499
rect 2087 2496 2099 2499
rect 3418 2496 3424 2508
rect 2087 2468 3424 2496
rect 2087 2465 2099 2468
rect 2041 2459 2099 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 4614 2456 4620 2508
rect 4672 2496 4678 2508
rect 5736 2505 5764 2536
rect 7282 2524 7288 2576
rect 7340 2524 7346 2576
rect 7944 2536 9628 2564
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 4672 2468 4721 2496
rect 4672 2456 4678 2468
rect 4709 2465 4721 2468
rect 4755 2465 4767 2499
rect 5721 2499 5779 2505
rect 4709 2459 4767 2465
rect 4816 2468 5672 2496
rect 2314 2428 2320 2440
rect 2227 2400 2320 2428
rect 2314 2388 2320 2400
rect 2372 2428 2378 2440
rect 2372 2400 2728 2428
rect 2372 2388 2378 2400
rect 2700 2292 2728 2400
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3145 2431 3203 2437
rect 3145 2428 3157 2431
rect 2832 2400 3157 2428
rect 2832 2388 2838 2400
rect 3145 2397 3157 2400
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 4816 2428 4844 2468
rect 3292 2400 3337 2428
rect 3988 2400 4844 2428
rect 4893 2431 4951 2437
rect 3292 2388 3298 2400
rect 3988 2292 4016 2400
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5534 2428 5540 2440
rect 4939 2400 5540 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5644 2428 5672 2468
rect 5721 2465 5733 2499
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5960 2468 6285 2496
rect 5960 2456 5966 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 7101 2499 7159 2505
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 7300 2496 7328 2524
rect 7944 2505 7972 2536
rect 7147 2468 7328 2496
rect 7929 2499 7987 2505
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 7929 2465 7941 2499
rect 7975 2465 7987 2499
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 7929 2459 7987 2465
rect 8036 2468 9045 2496
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5644 2400 5825 2428
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2428 7435 2431
rect 7558 2428 7564 2440
rect 7423 2400 7564 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 6457 2363 6515 2369
rect 6457 2360 6469 2363
rect 4120 2332 6469 2360
rect 4120 2320 4126 2332
rect 6457 2329 6469 2332
rect 6503 2329 6515 2363
rect 6457 2323 6515 2329
rect 2700 2264 4016 2292
rect 4798 2252 4804 2304
rect 4856 2292 4862 2304
rect 8036 2292 8064 2468
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9600 2496 9628 2536
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 11238 2564 11244 2576
rect 9916 2536 10548 2564
rect 9916 2524 9922 2536
rect 10226 2496 10232 2508
rect 9600 2468 10232 2496
rect 9033 2459 9091 2465
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 10520 2505 10548 2536
rect 10796 2536 11244 2564
rect 10505 2499 10563 2505
rect 10505 2465 10517 2499
rect 10551 2496 10563 2499
rect 10594 2496 10600 2508
rect 10551 2468 10600 2496
rect 10551 2465 10563 2468
rect 10505 2459 10563 2465
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2428 8263 2431
rect 8478 2428 8484 2440
rect 8251 2400 8484 2428
rect 8251 2397 8263 2400
rect 8205 2391 8263 2397
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9490 2428 9496 2440
rect 9355 2400 9496 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9490 2388 9496 2400
rect 9548 2428 9554 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 9548 2400 10701 2428
rect 9548 2388 9554 2400
rect 10689 2397 10701 2400
rect 10735 2428 10747 2431
rect 10796 2428 10824 2536
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 11054 2496 11060 2508
rect 11015 2468 11060 2496
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11146 2456 11152 2508
rect 11204 2496 11210 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11204 2468 11805 2496
rect 11204 2456 11210 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12400 2468 12633 2496
rect 12400 2456 12406 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 16592 2496 16620 2595
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 16761 2499 16819 2505
rect 16761 2496 16773 2499
rect 16592 2468 16773 2496
rect 12621 2459 12679 2465
rect 16761 2465 16773 2468
rect 16807 2465 16819 2499
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 16761 2459 16819 2465
rect 16868 2468 17509 2496
rect 10735 2400 10824 2428
rect 11241 2431 11299 2437
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 11241 2397 11253 2431
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9030 2360 9036 2372
rect 8711 2332 9036 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 10318 2320 10324 2372
rect 10376 2360 10382 2372
rect 11256 2360 11284 2391
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11388 2400 11989 2428
rect 11388 2388 11394 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12216 2400 12817 2428
rect 12216 2388 12222 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 16390 2388 16396 2440
rect 16448 2428 16454 2440
rect 16868 2428 16896 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 17034 2428 17040 2440
rect 16448 2400 16896 2428
rect 16995 2400 17040 2428
rect 16448 2388 16454 2400
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 17770 2428 17776 2440
rect 17731 2400 17776 2428
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 10376 2332 11284 2360
rect 10376 2320 10382 2332
rect 4856 2264 8064 2292
rect 4856 2252 4862 2264
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 1854 2048 1860 2100
rect 1912 2088 1918 2100
rect 16390 2088 16396 2100
rect 1912 2060 16396 2088
rect 1912 2048 1918 2060
rect 16390 2048 16396 2060
rect 16448 2048 16454 2100
rect 1210 1980 1216 2032
rect 1268 2020 1274 2032
rect 9214 2020 9220 2032
rect 1268 1992 9220 2020
rect 1268 1980 1274 1992
rect 9214 1980 9220 1992
rect 9272 1980 9278 2032
rect 3510 1300 3516 1352
rect 3568 1340 3574 1352
rect 6638 1340 6644 1352
rect 3568 1312 6644 1340
rect 3568 1300 3574 1312
rect 6638 1300 6644 1312
rect 6696 1300 6702 1352
rect 3418 552 3424 604
rect 3476 592 3482 604
rect 5994 592 6000 604
rect 3476 564 6000 592
rect 3476 552 3482 564
rect 5994 552 6000 564
rect 6052 552 6058 604
<< via1 >>
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 2780 14560 2832 14612
rect 4988 14560 5040 14612
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 2044 14424 2096 14476
rect 5172 14424 5224 14476
rect 3056 14356 3108 14408
rect 4068 14356 4120 14408
rect 17684 14356 17736 14408
rect 1676 14288 1728 14340
rect 14648 14288 14700 14340
rect 5172 14263 5224 14272
rect 5172 14229 5181 14263
rect 5181 14229 5215 14263
rect 5215 14229 5224 14263
rect 5172 14220 5224 14229
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 3424 14016 3476 14068
rect 2780 13880 2832 13932
rect 11796 14016 11848 14068
rect 16212 14016 16264 14068
rect 17684 14016 17736 14068
rect 16856 13948 16908 14000
rect 6368 13923 6420 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 3056 13855 3108 13864
rect 1676 13744 1728 13796
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3976 13812 4028 13864
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 7564 13923 7616 13932
rect 7564 13889 7573 13923
rect 7573 13889 7607 13923
rect 7607 13889 7616 13923
rect 7564 13880 7616 13889
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 14924 13880 14976 13932
rect 7288 13812 7340 13864
rect 7748 13812 7800 13864
rect 2228 13676 2280 13728
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 11612 13744 11664 13796
rect 12348 13744 12400 13796
rect 14648 13812 14700 13864
rect 17224 13812 17276 13864
rect 18236 13812 18288 13864
rect 7380 13719 7432 13728
rect 7380 13685 7389 13719
rect 7389 13685 7423 13719
rect 7423 13685 7432 13719
rect 7380 13676 7432 13685
rect 7472 13719 7524 13728
rect 7472 13685 7481 13719
rect 7481 13685 7515 13719
rect 7515 13685 7524 13719
rect 7472 13676 7524 13685
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 2872 13472 2924 13524
rect 5724 13472 5776 13524
rect 7288 13472 7340 13524
rect 14648 13472 14700 13524
rect 1860 13447 1912 13456
rect 1860 13413 1869 13447
rect 1869 13413 1903 13447
rect 1903 13413 1912 13447
rect 1860 13404 1912 13413
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2044 13336 2096 13388
rect 2228 13336 2280 13388
rect 8208 13404 8260 13456
rect 6828 13336 6880 13388
rect 7196 13336 7248 13388
rect 5724 13268 5776 13320
rect 6276 13200 6328 13252
rect 6644 13268 6696 13320
rect 9036 13336 9088 13388
rect 9772 13336 9824 13388
rect 16212 13336 16264 13388
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 8852 13311 8904 13320
rect 8852 13277 8861 13311
rect 8861 13277 8895 13311
rect 8895 13277 8904 13311
rect 8852 13268 8904 13277
rect 10968 13311 11020 13320
rect 8576 13200 8628 13252
rect 8760 13200 8812 13252
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 6092 13132 6144 13184
rect 8484 13132 8536 13184
rect 10968 13132 11020 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 2964 12928 3016 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 10784 12928 10836 12980
rect 4528 12860 4580 12912
rect 2688 12792 2740 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 1768 12724 1820 12776
rect 4068 12792 4120 12844
rect 7196 12860 7248 12912
rect 13820 12860 13872 12912
rect 15568 12860 15620 12912
rect 15752 12860 15804 12912
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 7288 12792 7340 12844
rect 7564 12792 7616 12844
rect 9128 12792 9180 12844
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 12072 12792 12124 12844
rect 12532 12792 12584 12844
rect 5724 12724 5776 12776
rect 3240 12656 3292 12708
rect 8852 12724 8904 12776
rect 10232 12724 10284 12776
rect 12348 12724 12400 12776
rect 15292 12724 15344 12776
rect 15568 12724 15620 12776
rect 6736 12656 6788 12708
rect 7564 12656 7616 12708
rect 9036 12656 9088 12708
rect 10140 12656 10192 12708
rect 10416 12656 10468 12708
rect 2320 12588 2372 12640
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 3056 12588 3108 12640
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 4436 12588 4488 12640
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 6368 12588 6420 12640
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 8300 12631 8352 12640
rect 8300 12597 8309 12631
rect 8309 12597 8343 12631
rect 8343 12597 8352 12631
rect 8300 12588 8352 12597
rect 8852 12588 8904 12640
rect 9772 12588 9824 12640
rect 9956 12588 10008 12640
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 11060 12588 11112 12640
rect 14648 12588 14700 12640
rect 17592 12588 17644 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 2596 12384 2648 12436
rect 2504 12316 2556 12368
rect 4528 12427 4580 12436
rect 4528 12393 4537 12427
rect 4537 12393 4571 12427
rect 4571 12393 4580 12427
rect 4528 12384 4580 12393
rect 4712 12384 4764 12436
rect 5264 12384 5316 12436
rect 6184 12384 6236 12436
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 7380 12384 7432 12436
rect 6644 12316 6696 12368
rect 2136 12291 2188 12300
rect 2136 12257 2145 12291
rect 2145 12257 2179 12291
rect 2179 12257 2188 12291
rect 2136 12248 2188 12257
rect 3240 12291 3292 12300
rect 3240 12257 3249 12291
rect 3249 12257 3283 12291
rect 3283 12257 3292 12291
rect 3240 12248 3292 12257
rect 5356 12248 5408 12300
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 2044 12180 2096 12232
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 4620 12223 4672 12232
rect 3148 12112 3200 12164
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 4804 12180 4856 12232
rect 6184 12180 6236 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 10324 12384 10376 12436
rect 16120 12427 16172 12436
rect 8576 12316 8628 12368
rect 8944 12316 8996 12368
rect 11612 12316 11664 12368
rect 9036 12248 9088 12300
rect 9956 12248 10008 12300
rect 10692 12291 10744 12300
rect 10692 12257 10701 12291
rect 10701 12257 10735 12291
rect 10735 12257 10744 12291
rect 10692 12248 10744 12257
rect 10784 12248 10836 12300
rect 16120 12393 16129 12427
rect 16129 12393 16163 12427
rect 16163 12393 16172 12427
rect 16120 12384 16172 12393
rect 17592 12427 17644 12436
rect 17592 12393 17601 12427
rect 17601 12393 17635 12427
rect 17635 12393 17644 12427
rect 17592 12384 17644 12393
rect 8392 12180 8444 12232
rect 9128 12180 9180 12232
rect 9220 12180 9272 12232
rect 11520 12180 11572 12232
rect 11612 12180 11664 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 15292 12248 15344 12300
rect 15752 12248 15804 12300
rect 17868 12316 17920 12368
rect 17960 12248 18012 12300
rect 14188 12180 14240 12232
rect 18144 12223 18196 12232
rect 3332 12044 3384 12096
rect 3700 12044 3752 12096
rect 7840 12044 7892 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 8576 12044 8628 12096
rect 15016 12112 15068 12164
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 10324 12044 10376 12053
rect 12348 12044 12400 12096
rect 15200 12044 15252 12096
rect 16488 12044 16540 12096
rect 17040 12044 17092 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 6276 11840 6328 11892
rect 3608 11772 3660 11824
rect 2596 11636 2648 11688
rect 2412 11568 2464 11620
rect 3424 11704 3476 11756
rect 4344 11747 4396 11756
rect 4344 11713 4353 11747
rect 4353 11713 4387 11747
rect 4387 11713 4396 11747
rect 4344 11704 4396 11713
rect 6828 11840 6880 11892
rect 4252 11636 4304 11688
rect 4068 11568 4120 11620
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 3516 11500 3568 11552
rect 5172 11500 5224 11552
rect 5632 11636 5684 11688
rect 6368 11636 6420 11688
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 10784 11840 10836 11892
rect 11244 11840 11296 11892
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 14372 11772 14424 11824
rect 7288 11568 7340 11620
rect 8116 11568 8168 11620
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 9220 11568 9272 11620
rect 10140 11679 10192 11688
rect 10140 11645 10149 11679
rect 10149 11645 10183 11679
rect 10183 11645 10192 11679
rect 10140 11636 10192 11645
rect 12072 11704 12124 11756
rect 13636 11704 13688 11756
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 17132 11704 17184 11756
rect 11244 11636 11296 11688
rect 12164 11636 12216 11688
rect 14004 11636 14056 11688
rect 14096 11636 14148 11688
rect 9680 11568 9732 11620
rect 11520 11568 11572 11620
rect 11888 11568 11940 11620
rect 13912 11568 13964 11620
rect 16580 11636 16632 11688
rect 16764 11636 16816 11688
rect 17776 11636 17828 11688
rect 14740 11568 14792 11620
rect 14832 11568 14884 11620
rect 10140 11500 10192 11552
rect 11244 11500 11296 11552
rect 13452 11500 13504 11552
rect 14280 11500 14332 11552
rect 15016 11500 15068 11552
rect 16120 11500 16172 11552
rect 16488 11500 16540 11552
rect 18328 11500 18380 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 1952 11271 2004 11280
rect 1952 11237 1961 11271
rect 1961 11237 1995 11271
rect 1995 11237 2004 11271
rect 2780 11296 2832 11348
rect 4344 11296 4396 11348
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 5816 11296 5868 11348
rect 8484 11296 8536 11348
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 10324 11296 10376 11348
rect 10692 11296 10744 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 1952 11228 2004 11237
rect 6368 11228 6420 11280
rect 9864 11228 9916 11280
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4712 11160 4764 11212
rect 5264 11160 5316 11212
rect 1952 11092 2004 11144
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 2872 11092 2924 11144
rect 3608 11092 3660 11144
rect 7656 11160 7708 11212
rect 6184 11092 6236 11144
rect 5264 11024 5316 11076
rect 3792 10956 3844 11008
rect 7840 10956 7892 11008
rect 8484 11160 8536 11212
rect 12256 11203 12308 11212
rect 12256 11169 12265 11203
rect 12265 11169 12299 11203
rect 12299 11169 12308 11203
rect 12256 11160 12308 11169
rect 14096 11228 14148 11280
rect 18144 11296 18196 11348
rect 18052 11228 18104 11280
rect 13728 11160 13780 11212
rect 15016 11160 15068 11212
rect 8116 11024 8168 11076
rect 8668 11092 8720 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 11520 11135 11572 11144
rect 10232 11092 10284 11101
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 12532 11135 12584 11144
rect 11980 11024 12032 11076
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 14096 11092 14148 11144
rect 15108 11092 15160 11144
rect 12716 11024 12768 11076
rect 11704 10956 11756 11008
rect 14740 10956 14792 11008
rect 17132 10956 17184 11008
rect 17316 10999 17368 11008
rect 17316 10965 17325 10999
rect 17325 10965 17359 10999
rect 17359 10965 17368 10999
rect 17316 10956 17368 10965
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2136 10752 2188 10804
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 5172 10752 5224 10804
rect 5632 10752 5684 10804
rect 5724 10752 5776 10804
rect 6552 10752 6604 10804
rect 6736 10752 6788 10804
rect 8760 10795 8812 10804
rect 8760 10761 8769 10795
rect 8769 10761 8803 10795
rect 8803 10761 8812 10795
rect 8760 10752 8812 10761
rect 8944 10752 8996 10804
rect 2780 10684 2832 10736
rect 3424 10684 3476 10736
rect 2596 10616 2648 10668
rect 3516 10659 3568 10668
rect 1492 10591 1544 10600
rect 1492 10557 1501 10591
rect 1501 10557 1535 10591
rect 1535 10557 1544 10591
rect 1492 10548 1544 10557
rect 2872 10548 2924 10600
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 4712 10616 4764 10668
rect 4344 10548 4396 10600
rect 6092 10616 6144 10668
rect 6736 10616 6788 10668
rect 5724 10591 5776 10600
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 9312 10616 9364 10668
rect 9588 10616 9640 10668
rect 10600 10752 10652 10804
rect 11520 10752 11572 10804
rect 11704 10752 11756 10804
rect 12624 10752 12676 10804
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14832 10752 14884 10804
rect 5724 10548 5776 10557
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3976 10412 4028 10464
rect 5172 10412 5224 10464
rect 6000 10412 6052 10464
rect 6276 10480 6328 10532
rect 8208 10548 8260 10600
rect 10508 10591 10560 10600
rect 10508 10557 10542 10591
rect 10542 10557 10560 10591
rect 10508 10548 10560 10557
rect 11704 10548 11756 10600
rect 18052 10684 18104 10736
rect 13820 10616 13872 10668
rect 14096 10616 14148 10668
rect 14464 10616 14516 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 16304 10616 16356 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 7840 10480 7892 10532
rect 7564 10412 7616 10464
rect 9864 10412 9916 10464
rect 10600 10480 10652 10532
rect 14004 10548 14056 10600
rect 14924 10548 14976 10600
rect 15292 10548 15344 10600
rect 15568 10548 15620 10600
rect 16120 10548 16172 10600
rect 17316 10548 17368 10600
rect 17684 10548 17736 10600
rect 12716 10523 12768 10532
rect 12716 10489 12750 10523
rect 12750 10489 12768 10523
rect 12716 10480 12768 10489
rect 13268 10480 13320 10532
rect 11796 10412 11848 10464
rect 13728 10412 13780 10464
rect 15568 10412 15620 10464
rect 16120 10412 16172 10464
rect 16396 10412 16448 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 3700 10208 3752 10260
rect 2412 10140 2464 10192
rect 3056 10115 3108 10124
rect 3056 10081 3065 10115
rect 3065 10081 3099 10115
rect 3099 10081 3108 10115
rect 3056 10072 3108 10081
rect 5816 10140 5868 10192
rect 6644 10140 6696 10192
rect 7288 10208 7340 10260
rect 8300 10208 8352 10260
rect 9036 10208 9088 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10692 10208 10744 10260
rect 7472 10140 7524 10192
rect 7656 10140 7708 10192
rect 8484 10140 8536 10192
rect 10048 10140 10100 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3240 10004 3292 10056
rect 3516 10004 3568 10056
rect 3884 10004 3936 10056
rect 2688 9936 2740 9988
rect 4712 10047 4764 10056
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 6736 10072 6788 10124
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 10600 10072 10652 10124
rect 5724 9936 5776 9988
rect 6828 9936 6880 9988
rect 4712 9868 4764 9920
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 14004 10208 14056 10260
rect 14188 10251 14240 10260
rect 14188 10217 14197 10251
rect 14197 10217 14231 10251
rect 14231 10217 14240 10251
rect 14188 10208 14240 10217
rect 14464 10208 14516 10260
rect 15016 10208 15068 10260
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 12808 10140 12860 10192
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 11704 10072 11756 10124
rect 14372 10072 14424 10124
rect 14832 10072 14884 10124
rect 15108 10072 15160 10124
rect 17132 10072 17184 10124
rect 17592 10072 17644 10124
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 13636 10004 13688 10056
rect 14464 10004 14516 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 16396 10004 16448 10056
rect 16764 10004 16816 10056
rect 17500 10047 17552 10056
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 17500 10004 17552 10013
rect 11152 9936 11204 9988
rect 13544 9979 13596 9988
rect 9036 9868 9088 9920
rect 11244 9868 11296 9920
rect 13544 9945 13553 9979
rect 13553 9945 13587 9979
rect 13587 9945 13596 9979
rect 13544 9936 13596 9945
rect 12716 9868 12768 9920
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 13268 9868 13320 9920
rect 14004 9868 14056 9920
rect 16304 9868 16356 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3424 9664 3476 9716
rect 4436 9664 4488 9716
rect 6184 9664 6236 9716
rect 5816 9596 5868 9648
rect 6276 9639 6328 9648
rect 6276 9605 6285 9639
rect 6285 9605 6319 9639
rect 6319 9605 6328 9639
rect 6276 9596 6328 9605
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 3792 9528 3844 9580
rect 4344 9528 4396 9580
rect 1400 9460 1452 9512
rect 2412 9460 2464 9512
rect 3608 9460 3660 9512
rect 4896 9503 4948 9512
rect 4896 9469 4930 9503
rect 4930 9469 4948 9503
rect 4896 9460 4948 9469
rect 2688 9392 2740 9444
rect 3056 9392 3108 9444
rect 3976 9435 4028 9444
rect 3976 9401 3985 9435
rect 3985 9401 4019 9435
rect 4019 9401 4028 9435
rect 3976 9392 4028 9401
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 3700 9324 3752 9376
rect 6644 9528 6696 9580
rect 6736 9528 6788 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10692 9664 10744 9716
rect 12256 9664 12308 9716
rect 12532 9664 12584 9716
rect 13820 9664 13872 9716
rect 16672 9664 16724 9716
rect 16764 9664 16816 9716
rect 17500 9664 17552 9716
rect 10968 9596 11020 9648
rect 12992 9596 13044 9648
rect 6184 9460 6236 9512
rect 6552 9460 6604 9512
rect 9036 9460 9088 9512
rect 9956 9503 10008 9512
rect 9956 9469 9990 9503
rect 9990 9469 10008 9503
rect 9956 9460 10008 9469
rect 6368 9392 6420 9444
rect 6644 9392 6696 9444
rect 7380 9392 7432 9444
rect 9772 9392 9824 9444
rect 9864 9392 9916 9444
rect 12532 9460 12584 9512
rect 7656 9324 7708 9376
rect 11888 9392 11940 9444
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 12164 9324 12216 9376
rect 12716 9460 12768 9512
rect 13728 9528 13780 9580
rect 13912 9571 13964 9580
rect 13912 9537 13921 9571
rect 13921 9537 13955 9571
rect 13955 9537 13964 9571
rect 13912 9528 13964 9537
rect 14740 9596 14792 9648
rect 15384 9596 15436 9648
rect 13636 9460 13688 9512
rect 14924 9528 14976 9580
rect 15108 9528 15160 9580
rect 14464 9460 14516 9512
rect 16304 9460 16356 9512
rect 16580 9460 16632 9512
rect 17868 9460 17920 9512
rect 14556 9392 14608 9444
rect 15660 9392 15712 9444
rect 17592 9367 17644 9376
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 17592 9324 17644 9333
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 3148 9120 3200 9172
rect 4896 9120 4948 9172
rect 7380 9163 7432 9172
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1952 8984 2004 9036
rect 3424 9052 3476 9104
rect 7380 9129 7389 9163
rect 7389 9129 7423 9163
rect 7423 9129 7432 9163
rect 7380 9120 7432 9129
rect 3608 8984 3660 9036
rect 4344 9027 4396 9036
rect 4344 8993 4378 9027
rect 4378 8993 4396 9027
rect 4344 8984 4396 8993
rect 8760 9052 8812 9104
rect 9128 9120 9180 9172
rect 10416 9120 10468 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 12164 9120 12216 9172
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 3148 8916 3200 8968
rect 5540 8916 5592 8968
rect 6552 8984 6604 9036
rect 6736 8984 6788 9036
rect 7840 8984 7892 9036
rect 7012 8916 7064 8968
rect 9864 8984 9916 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10968 9095 11020 9104
rect 10968 9061 11002 9095
rect 11002 9061 11020 9095
rect 10968 9052 11020 9061
rect 13452 9052 13504 9104
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 14832 9052 14884 9104
rect 15108 9052 15160 9104
rect 16764 9095 16816 9104
rect 13636 8984 13688 9036
rect 14372 8984 14424 9036
rect 15660 8984 15712 9036
rect 16304 8984 16356 9036
rect 16764 9061 16798 9095
rect 16798 9061 16816 9095
rect 16764 9052 16816 9061
rect 10232 8916 10284 8968
rect 10692 8959 10744 8968
rect 8944 8848 8996 8900
rect 2688 8780 2740 8832
rect 3056 8780 3108 8832
rect 3608 8780 3660 8832
rect 4804 8780 4856 8832
rect 6000 8780 6052 8832
rect 7932 8780 7984 8832
rect 9772 8848 9824 8900
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 11796 8916 11848 8968
rect 13268 8916 13320 8968
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 11060 8780 11112 8832
rect 12532 8780 12584 8832
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 17684 8780 17736 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 3608 8576 3660 8628
rect 4344 8576 4396 8628
rect 6736 8576 6788 8628
rect 7288 8576 7340 8628
rect 8944 8576 8996 8628
rect 1492 8440 1544 8492
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 2228 8440 2280 8492
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 1308 8372 1360 8424
rect 4712 8440 4764 8492
rect 4896 8440 4948 8492
rect 5540 8440 5592 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 7012 8440 7064 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 9772 8576 9824 8628
rect 11704 8576 11756 8628
rect 16304 8576 16356 8628
rect 9588 8508 9640 8560
rect 10508 8508 10560 8560
rect 4068 8415 4120 8424
rect 2228 8304 2280 8356
rect 2688 8347 2740 8356
rect 2688 8313 2700 8347
rect 2700 8313 2740 8347
rect 2688 8304 2740 8313
rect 3148 8304 3200 8356
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4804 8372 4856 8424
rect 1860 8236 1912 8288
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 4436 8304 4488 8356
rect 6000 8372 6052 8424
rect 8024 8372 8076 8424
rect 8392 8372 8444 8424
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 8760 8372 8812 8381
rect 10140 8372 10192 8424
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 18328 8508 18380 8560
rect 10968 8440 11020 8449
rect 11152 8372 11204 8424
rect 11244 8372 11296 8424
rect 4988 8236 5040 8288
rect 6828 8304 6880 8356
rect 11060 8304 11112 8356
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 14556 8440 14608 8492
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 12624 8372 12676 8424
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 8116 8236 8168 8288
rect 8300 8236 8352 8288
rect 8852 8236 8904 8288
rect 11244 8236 11296 8288
rect 11336 8236 11388 8288
rect 11704 8279 11756 8288
rect 11704 8245 11713 8279
rect 11713 8245 11747 8279
rect 11747 8245 11756 8279
rect 14372 8304 14424 8356
rect 17868 8440 17920 8492
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 17960 8304 18012 8356
rect 11704 8236 11756 8245
rect 12164 8236 12216 8288
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 14740 8236 14792 8288
rect 16120 8236 16172 8288
rect 17040 8236 17092 8288
rect 17500 8279 17552 8288
rect 17500 8245 17509 8279
rect 17509 8245 17543 8279
rect 17543 8245 17552 8279
rect 17500 8236 17552 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3148 8032 3200 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 5172 8032 5224 8084
rect 6736 8075 6788 8084
rect 6736 8041 6745 8075
rect 6745 8041 6779 8075
rect 6779 8041 6788 8075
rect 6736 8032 6788 8041
rect 7564 8032 7616 8084
rect 5080 7964 5132 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 3516 7896 3568 7948
rect 5264 7896 5316 7948
rect 5540 7896 5592 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2228 7760 2280 7812
rect 3424 7828 3476 7880
rect 4436 7828 4488 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 4344 7760 4396 7812
rect 5080 7760 5132 7812
rect 5448 7760 5500 7812
rect 3792 7692 3844 7744
rect 5540 7692 5592 7744
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 7564 7896 7616 7948
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 8116 7939 8168 7948
rect 8116 7905 8150 7939
rect 8150 7905 8168 7939
rect 8116 7896 8168 7905
rect 5724 7828 5776 7837
rect 6552 7828 6604 7880
rect 6644 7828 6696 7880
rect 7380 7828 7432 7880
rect 7748 7828 7800 7880
rect 6644 7692 6696 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 11796 8032 11848 8084
rect 10784 7964 10836 8016
rect 10508 7896 10560 7948
rect 11428 7964 11480 8016
rect 14188 8032 14240 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 15200 8032 15252 8084
rect 15476 8032 15528 8084
rect 12164 7964 12216 8016
rect 12072 7896 12124 7948
rect 17500 8032 17552 8084
rect 17868 7964 17920 8016
rect 10324 7828 10376 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11244 7828 11296 7880
rect 10876 7760 10928 7812
rect 12348 7760 12400 7812
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 14096 7828 14148 7880
rect 15200 7828 15252 7880
rect 16212 7828 16264 7880
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 12256 7692 12308 7744
rect 12624 7692 12676 7744
rect 12808 7692 12860 7744
rect 12992 7692 13044 7744
rect 15476 7760 15528 7812
rect 16120 7760 16172 7812
rect 15200 7692 15252 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 1860 7488 1912 7540
rect 5816 7488 5868 7540
rect 6092 7531 6144 7540
rect 6092 7497 6101 7531
rect 6101 7497 6135 7531
rect 6135 7497 6144 7531
rect 6092 7488 6144 7497
rect 5724 7420 5776 7472
rect 9036 7488 9088 7540
rect 10232 7488 10284 7540
rect 10508 7488 10560 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 15568 7488 15620 7540
rect 16212 7531 16264 7540
rect 16212 7497 16221 7531
rect 16221 7497 16255 7531
rect 16255 7497 16264 7531
rect 16212 7488 16264 7497
rect 16856 7488 16908 7540
rect 8944 7420 8996 7472
rect 12440 7420 12492 7472
rect 12624 7420 12676 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 3424 7352 3476 7404
rect 3792 7352 3844 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 4436 7352 4488 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 2136 7284 2188 7336
rect 3884 7284 3936 7336
rect 11520 7352 11572 7404
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 11796 7352 11848 7404
rect 7840 7327 7892 7336
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 8208 7284 8260 7336
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 9036 7284 9088 7336
rect 13176 7352 13228 7404
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 12440 7284 12492 7336
rect 12808 7284 12860 7336
rect 12992 7284 13044 7336
rect 13636 7327 13688 7336
rect 13636 7293 13645 7327
rect 13645 7293 13679 7327
rect 13679 7293 13688 7327
rect 13636 7284 13688 7293
rect 14096 7284 14148 7336
rect 14832 7327 14884 7336
rect 2596 7148 2648 7200
rect 5448 7216 5500 7268
rect 6276 7216 6328 7268
rect 8852 7216 8904 7268
rect 9772 7216 9824 7268
rect 11244 7216 11296 7268
rect 12624 7216 12676 7268
rect 5724 7148 5776 7200
rect 6184 7148 6236 7200
rect 6552 7148 6604 7200
rect 7932 7148 7984 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 8208 7148 8260 7200
rect 11336 7148 11388 7200
rect 11980 7148 12032 7200
rect 12164 7148 12216 7200
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 13820 7216 13872 7268
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 16580 7352 16632 7404
rect 16672 7352 16724 7404
rect 17868 7352 17920 7404
rect 16120 7216 16172 7268
rect 17684 7284 17736 7336
rect 17960 7284 18012 7336
rect 15384 7148 15436 7200
rect 18236 7191 18288 7200
rect 18236 7157 18245 7191
rect 18245 7157 18279 7191
rect 18279 7157 18288 7191
rect 18236 7148 18288 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 5540 6944 5592 6996
rect 7932 6944 7984 6996
rect 8576 6944 8628 6996
rect 9772 6944 9824 6996
rect 9864 6944 9916 6996
rect 1768 6808 1820 6860
rect 3516 6876 3568 6928
rect 1400 6740 1452 6792
rect 4620 6808 4672 6860
rect 3424 6672 3476 6724
rect 3608 6604 3660 6656
rect 4436 6740 4488 6792
rect 5632 6604 5684 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 7380 6808 7432 6860
rect 9220 6876 9272 6928
rect 11704 6944 11756 6996
rect 13268 6944 13320 6996
rect 13820 6944 13872 6996
rect 14096 6944 14148 6996
rect 16580 6944 16632 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 10416 6808 10468 6860
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 8116 6783 8168 6792
rect 6276 6740 6328 6749
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 12348 6808 12400 6860
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 14832 6876 14884 6928
rect 13452 6808 13504 6860
rect 16212 6876 16264 6928
rect 9772 6672 9824 6724
rect 12072 6672 12124 6724
rect 6460 6604 6512 6656
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 12164 6604 12216 6656
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 13360 6740 13412 6792
rect 15108 6740 15160 6792
rect 17684 6808 17736 6860
rect 17868 6783 17920 6792
rect 13912 6604 13964 6656
rect 14280 6604 14332 6656
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 16396 6604 16448 6656
rect 17776 6672 17828 6724
rect 17132 6647 17184 6656
rect 17132 6613 17141 6647
rect 17141 6613 17175 6647
rect 17175 6613 17184 6647
rect 17132 6604 17184 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 1768 6400 1820 6452
rect 1952 6400 2004 6452
rect 1400 6332 1452 6384
rect 2136 6264 2188 6316
rect 2320 6264 2372 6316
rect 1768 6196 1820 6248
rect 2504 6196 2556 6248
rect 4344 6400 4396 6452
rect 6736 6400 6788 6452
rect 8116 6400 8168 6452
rect 2964 6128 3016 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 2228 6060 2280 6112
rect 4068 6196 4120 6248
rect 5448 6264 5500 6316
rect 5908 6264 5960 6316
rect 6184 6196 6236 6248
rect 6460 6307 6512 6316
rect 6460 6273 6469 6307
rect 6469 6273 6503 6307
rect 6503 6273 6512 6307
rect 6460 6264 6512 6273
rect 7380 6264 7432 6316
rect 8208 6264 8260 6316
rect 10968 6400 11020 6452
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 11244 6400 11296 6452
rect 12256 6400 12308 6452
rect 12900 6400 12952 6452
rect 13360 6400 13412 6452
rect 14648 6400 14700 6452
rect 14832 6400 14884 6452
rect 15660 6400 15712 6452
rect 10324 6332 10376 6384
rect 13636 6332 13688 6384
rect 17868 6332 17920 6384
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 13176 6264 13228 6316
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 7472 6239 7524 6248
rect 3424 6128 3476 6180
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 8116 6196 8168 6248
rect 8576 6196 8628 6248
rect 9496 6196 9548 6248
rect 9588 6196 9640 6248
rect 10968 6196 11020 6248
rect 4068 6060 4120 6112
rect 4436 6060 4488 6112
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 4896 6060 4948 6112
rect 5724 6060 5776 6112
rect 8484 6128 8536 6180
rect 10324 6128 10376 6180
rect 11612 6171 11664 6180
rect 11612 6137 11621 6171
rect 11621 6137 11655 6171
rect 11655 6137 11664 6171
rect 11612 6128 11664 6137
rect 12532 6196 12584 6248
rect 14096 6196 14148 6248
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 14924 6264 14976 6316
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 14556 6196 14608 6248
rect 16396 6264 16448 6316
rect 16672 6264 16724 6316
rect 17408 6264 17460 6316
rect 17776 6264 17828 6316
rect 17684 6196 17736 6248
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 9956 6060 10008 6112
rect 11796 6060 11848 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 14004 6060 14056 6112
rect 14464 6060 14516 6112
rect 14832 6103 14884 6112
rect 14832 6069 14841 6103
rect 14841 6069 14875 6103
rect 14875 6069 14884 6103
rect 14832 6060 14884 6069
rect 18144 6128 18196 6180
rect 16120 6060 16172 6112
rect 16488 6060 16540 6112
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 17592 6060 17644 6112
rect 17868 6060 17920 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 5724 5899 5776 5908
rect 5724 5865 5733 5899
rect 5733 5865 5767 5899
rect 5767 5865 5776 5899
rect 5724 5856 5776 5865
rect 6552 5856 6604 5908
rect 7564 5856 7616 5908
rect 7748 5856 7800 5908
rect 8208 5856 8260 5908
rect 8484 5856 8536 5908
rect 9220 5856 9272 5908
rect 11888 5899 11940 5908
rect 11888 5865 11897 5899
rect 11897 5865 11931 5899
rect 11931 5865 11940 5899
rect 11888 5856 11940 5865
rect 4160 5788 4212 5840
rect 4344 5831 4396 5840
rect 4344 5797 4378 5831
rect 4378 5797 4396 5831
rect 4344 5788 4396 5797
rect 4804 5788 4856 5840
rect 5908 5788 5960 5840
rect 1768 5720 1820 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 3424 5652 3476 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 6460 5652 6512 5704
rect 6736 5652 6788 5704
rect 8116 5720 8168 5772
rect 9036 5720 9088 5772
rect 9956 5763 10008 5772
rect 8208 5652 8260 5704
rect 9956 5729 9979 5763
rect 9979 5729 10008 5763
rect 9956 5720 10008 5729
rect 10692 5720 10744 5772
rect 13360 5720 13412 5772
rect 13728 5788 13780 5840
rect 14832 5856 14884 5908
rect 16856 5856 16908 5908
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 16212 5788 16264 5840
rect 14004 5720 14056 5772
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 11980 5695 12032 5704
rect 9680 5652 9732 5661
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 2872 5516 2924 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 4252 5516 4304 5568
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 6000 5516 6052 5568
rect 8116 5584 8168 5636
rect 8392 5584 8444 5636
rect 9588 5584 9640 5636
rect 10692 5584 10744 5636
rect 12440 5584 12492 5636
rect 13176 5584 13228 5636
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 13544 5516 13596 5568
rect 14648 5652 14700 5704
rect 14924 5652 14976 5704
rect 17132 5720 17184 5772
rect 16396 5652 16448 5704
rect 14556 5516 14608 5568
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 17776 5516 17828 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3516 5312 3568 5364
rect 3700 5312 3752 5364
rect 6184 5312 6236 5364
rect 1400 5176 1452 5228
rect 2044 5108 2096 5160
rect 2136 5040 2188 5092
rect 2780 5040 2832 5092
rect 3240 5040 3292 5092
rect 8024 5244 8076 5296
rect 3516 5176 3568 5228
rect 4344 5176 4396 5228
rect 4436 5176 4488 5228
rect 7380 5219 7432 5228
rect 4804 5108 4856 5160
rect 4436 5083 4488 5092
rect 4436 5049 4445 5083
rect 4445 5049 4479 5083
rect 4479 5049 4488 5083
rect 4436 5040 4488 5049
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 11888 5312 11940 5364
rect 10416 5244 10468 5296
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 9496 5219 9548 5228
rect 8392 5176 8444 5185
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 5448 5108 5500 5160
rect 6092 5108 6144 5160
rect 7932 5108 7984 5160
rect 12532 5244 12584 5296
rect 11336 5176 11388 5228
rect 13728 5312 13780 5364
rect 14648 5312 14700 5364
rect 15016 5312 15068 5364
rect 17316 5312 17368 5364
rect 17132 5176 17184 5228
rect 17592 5176 17644 5228
rect 5264 5040 5316 5092
rect 5816 5040 5868 5092
rect 9680 5040 9732 5092
rect 10968 5108 11020 5160
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 12440 5108 12492 5160
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 14924 5108 14976 5117
rect 17776 5108 17828 5160
rect 1952 4972 2004 5024
rect 2228 4972 2280 5024
rect 4344 4972 4396 5024
rect 5540 4972 5592 5024
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6460 4972 6512 5024
rect 8484 4972 8536 5024
rect 8760 4972 8812 5024
rect 11244 5040 11296 5092
rect 12164 5040 12216 5092
rect 14004 5040 14056 5092
rect 17040 5040 17092 5092
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 11520 4972 11572 5024
rect 11704 4972 11756 5024
rect 12532 4972 12584 5024
rect 14372 4972 14424 5024
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 17408 5015 17460 5024
rect 17408 4981 17417 5015
rect 17417 4981 17451 5015
rect 17451 4981 17460 5015
rect 17408 4972 17460 4981
rect 18328 4972 18380 5024
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 2596 4768 2648 4820
rect 3332 4768 3384 4820
rect 5264 4768 5316 4820
rect 6460 4768 6512 4820
rect 8760 4768 8812 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 11520 4811 11572 4820
rect 1492 4632 1544 4684
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 1216 4564 1268 4616
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 3240 4632 3292 4684
rect 4252 4700 4304 4752
rect 5816 4700 5868 4752
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14372 4768 14424 4820
rect 15108 4768 15160 4820
rect 15292 4768 15344 4820
rect 16488 4768 16540 4820
rect 17684 4768 17736 4820
rect 10324 4700 10376 4752
rect 2504 4564 2556 4573
rect 4344 4632 4396 4684
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2504 4428 2556 4480
rect 3792 4564 3844 4616
rect 4160 4564 4212 4616
rect 5724 4632 5776 4684
rect 5908 4632 5960 4684
rect 6460 4632 6512 4684
rect 7380 4632 7432 4684
rect 8944 4675 8996 4684
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 4804 4496 4856 4548
rect 5448 4496 5500 4548
rect 5080 4428 5132 4480
rect 5540 4428 5592 4480
rect 7932 4564 7984 4616
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9312 4564 9364 4616
rect 8300 4496 8352 4548
rect 9588 4496 9640 4548
rect 10048 4496 10100 4548
rect 6736 4428 6788 4480
rect 8024 4428 8076 4480
rect 9680 4428 9732 4480
rect 9772 4428 9824 4480
rect 10324 4428 10376 4480
rect 13176 4700 13228 4752
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 11336 4632 11388 4684
rect 13728 4632 13780 4684
rect 14280 4632 14332 4684
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 17500 4632 17552 4684
rect 11520 4564 11572 4616
rect 12164 4607 12216 4616
rect 12164 4573 12173 4607
rect 12173 4573 12207 4607
rect 12207 4573 12216 4607
rect 12164 4564 12216 4573
rect 12440 4564 12492 4616
rect 15660 4564 15712 4616
rect 17592 4607 17644 4616
rect 11612 4496 11664 4548
rect 15384 4496 15436 4548
rect 15568 4496 15620 4548
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 14924 4428 14976 4480
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 6644 4224 6696 4276
rect 8024 4224 8076 4276
rect 8576 4224 8628 4276
rect 9772 4224 9824 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 5816 4020 5868 4072
rect 388 3952 440 4004
rect 4620 3952 4672 4004
rect 6276 4088 6328 4140
rect 6644 4088 6696 4140
rect 7012 4020 7064 4072
rect 10324 4088 10376 4140
rect 13728 4224 13780 4276
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 14648 4224 14700 4276
rect 15660 4224 15712 4276
rect 8300 4020 8352 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 9220 4020 9272 4072
rect 6552 3952 6604 4004
rect 6644 3952 6696 4004
rect 3792 3884 3844 3936
rect 4436 3884 4488 3936
rect 5264 3884 5316 3936
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 5632 3884 5684 3893
rect 6184 3884 6236 3936
rect 7564 3884 7616 3936
rect 9312 3952 9364 4004
rect 10140 3952 10192 4004
rect 12716 3995 12768 4004
rect 10968 3884 11020 3936
rect 12716 3961 12750 3995
rect 12750 3961 12768 3995
rect 12716 3952 12768 3961
rect 12164 3884 12216 3936
rect 14372 3884 14424 3936
rect 16396 4020 16448 4072
rect 16948 4088 17000 4140
rect 17776 4156 17828 4208
rect 17040 4020 17092 4072
rect 17500 4020 17552 4072
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 16764 3952 16816 4004
rect 17592 3952 17644 4004
rect 15568 3884 15620 3936
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 1400 3680 1452 3732
rect 2320 3680 2372 3732
rect 2412 3680 2464 3732
rect 3056 3612 3108 3664
rect 2412 3544 2464 3596
rect 3240 3680 3292 3732
rect 4528 3680 4580 3732
rect 5632 3680 5684 3732
rect 6736 3680 6788 3732
rect 3700 3612 3752 3664
rect 5080 3655 5132 3664
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 5080 3621 5089 3655
rect 5089 3621 5123 3655
rect 5123 3621 5132 3655
rect 5080 3612 5132 3621
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 2504 3408 2556 3460
rect 4896 3476 4948 3528
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 5540 3476 5592 3528
rect 7472 3544 7524 3596
rect 8392 3680 8444 3732
rect 9680 3680 9732 3732
rect 11520 3680 11572 3732
rect 11980 3723 12032 3732
rect 11980 3689 11989 3723
rect 11989 3689 12023 3723
rect 12023 3689 12032 3723
rect 11980 3680 12032 3689
rect 12256 3680 12308 3732
rect 12532 3680 12584 3732
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 14464 3680 14516 3732
rect 17224 3680 17276 3732
rect 17408 3680 17460 3732
rect 9128 3612 9180 3664
rect 10600 3612 10652 3664
rect 15016 3612 15068 3664
rect 9588 3544 9640 3596
rect 10140 3544 10192 3596
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 12624 3544 12676 3596
rect 14372 3544 14424 3596
rect 16488 3612 16540 3664
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 17040 3587 17092 3596
rect 17040 3553 17049 3587
rect 17049 3553 17083 3587
rect 17083 3553 17092 3587
rect 17040 3544 17092 3553
rect 10416 3476 10468 3528
rect 11244 3476 11296 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 15660 3476 15712 3528
rect 18052 3519 18104 3528
rect 3516 3408 3568 3460
rect 4344 3340 4396 3392
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 5540 3340 5592 3392
rect 6460 3340 6512 3392
rect 7196 3340 7248 3392
rect 11704 3408 11756 3460
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 18512 3408 18564 3460
rect 9312 3340 9364 3392
rect 11060 3340 11112 3392
rect 11612 3340 11664 3392
rect 17316 3340 17368 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 2688 3136 2740 3188
rect 6092 3136 6144 3188
rect 7196 3136 7248 3188
rect 8944 3136 8996 3188
rect 9588 3179 9640 3188
rect 9588 3145 9597 3179
rect 9597 3145 9631 3179
rect 9631 3145 9640 3179
rect 9588 3136 9640 3145
rect 9772 3136 9824 3188
rect 10508 3136 10560 3188
rect 4988 3068 5040 3120
rect 5448 3068 5500 3120
rect 7380 3068 7432 3120
rect 8760 3068 8812 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2780 3000 2832 3052
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 3332 2932 3384 2984
rect 6184 3000 6236 3052
rect 6276 3043 6328 3052
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 6276 3000 6328 3009
rect 6552 3000 6604 3052
rect 7748 3000 7800 3052
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 8300 3000 8352 3052
rect 10692 3068 10744 3120
rect 11428 3136 11480 3188
rect 13636 3136 13688 3188
rect 18420 3136 18472 3188
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 9312 3000 9364 3052
rect 10876 3000 10928 3052
rect 11244 3043 11296 3052
rect 11244 3009 11253 3043
rect 11253 3009 11287 3043
rect 11287 3009 11296 3043
rect 11244 3000 11296 3009
rect 6460 2932 6512 2984
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 2412 2864 2464 2916
rect 2780 2864 2832 2916
rect 4252 2864 4304 2916
rect 6092 2907 6144 2916
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 4712 2839 4764 2848
rect 3700 2796 3752 2805
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 6092 2873 6101 2907
rect 6101 2873 6135 2907
rect 6135 2873 6144 2907
rect 6092 2864 6144 2873
rect 6276 2864 6328 2916
rect 6736 2864 6788 2916
rect 9404 2932 9456 2984
rect 10968 2975 11020 2984
rect 9496 2864 9548 2916
rect 10968 2941 10977 2975
rect 10977 2941 11011 2975
rect 11011 2941 11020 2975
rect 10968 2932 11020 2941
rect 11336 2932 11388 2984
rect 12072 3068 12124 3120
rect 12716 3000 12768 3052
rect 13912 3068 13964 3120
rect 13820 2975 13872 2984
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 15476 3000 15528 3052
rect 15200 2975 15252 2984
rect 15200 2941 15209 2975
rect 15209 2941 15243 2975
rect 15243 2941 15252 2975
rect 15200 2932 15252 2941
rect 16120 2932 16172 2984
rect 16580 2932 16632 2984
rect 17408 3000 17460 3052
rect 19432 3000 19484 3052
rect 17316 2932 17368 2984
rect 6368 2796 6420 2848
rect 8024 2796 8076 2848
rect 9864 2796 9916 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 14096 2864 14148 2916
rect 14832 2864 14884 2916
rect 16764 2907 16816 2916
rect 16764 2873 16773 2907
rect 16773 2873 16807 2907
rect 16807 2873 16816 2907
rect 16764 2864 16816 2873
rect 10048 2796 10100 2805
rect 10784 2796 10836 2848
rect 17500 2796 17552 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1768 2592 1820 2644
rect 2044 2592 2096 2644
rect 2780 2592 2832 2644
rect 3700 2524 3752 2576
rect 4344 2592 4396 2644
rect 4712 2592 4764 2644
rect 5356 2592 5408 2644
rect 5724 2592 5776 2644
rect 5448 2524 5500 2576
rect 7840 2592 7892 2644
rect 8760 2592 8812 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 10508 2592 10560 2644
rect 12440 2592 12492 2644
rect 3424 2456 3476 2508
rect 4620 2456 4672 2508
rect 7288 2524 7340 2576
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 2780 2388 2832 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 5540 2388 5592 2440
rect 5908 2456 5960 2508
rect 7564 2388 7616 2440
rect 4068 2320 4120 2372
rect 4804 2252 4856 2304
rect 9864 2524 9916 2576
rect 10232 2456 10284 2508
rect 10600 2456 10652 2508
rect 8484 2388 8536 2440
rect 9496 2388 9548 2440
rect 11244 2524 11296 2576
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 11152 2456 11204 2508
rect 12348 2456 12400 2508
rect 16856 2592 16908 2644
rect 9036 2320 9088 2372
rect 10324 2320 10376 2372
rect 11336 2388 11388 2440
rect 12164 2388 12216 2440
rect 16396 2388 16448 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 1860 2048 1912 2100
rect 16396 2048 16448 2100
rect 1216 1980 1268 2032
rect 9220 1980 9272 2032
rect 3516 1300 3568 1352
rect 6644 1300 6696 1352
rect 3424 552 3476 604
rect 6000 552 6052 604
<< metal2 >>
rect 1674 16520 1730 17000
rect 4066 16824 4122 16833
rect 4066 16759 4122 16768
rect 3422 16552 3478 16561
rect 1688 14346 1716 16520
rect 3422 16487 3478 16496
rect 2962 16144 3018 16153
rect 2962 16079 3018 16088
rect 2870 15192 2926 15201
rect 2870 15127 2926 15136
rect 2778 14784 2834 14793
rect 2778 14719 2834 14728
rect 2792 14618 2820 14719
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2778 14512 2834 14521
rect 2044 14476 2096 14482
rect 2778 14447 2834 14456
rect 2044 14418 2096 14424
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1780 14113 1808 14350
rect 1766 14104 1822 14113
rect 1766 14039 1822 14048
rect 1860 13864 1912 13870
rect 1858 13832 1860 13841
rect 1912 13832 1914 13841
rect 1676 13796 1728 13802
rect 1858 13767 1914 13776
rect 1676 13738 1728 13744
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1306 11520 1362 11529
rect 1306 11455 1362 11464
rect 570 9072 626 9081
rect 570 9007 626 9016
rect 584 8537 612 9007
rect 570 8528 626 8537
rect 570 8463 626 8472
rect 1320 8430 1348 11455
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1504 10606 1532 10911
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9518 1440 9998
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9042 1440 9454
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1308 8424 1360 8430
rect 1308 8366 1360 8372
rect 1214 8120 1270 8129
rect 1214 8055 1270 8064
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1228 4622 1256 8055
rect 1412 7954 1440 8055
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1306 7440 1362 7449
rect 1306 7375 1362 7384
rect 1320 5001 1348 7375
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6390 1440 6734
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1412 5234 1440 6326
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1306 4992 1362 5001
rect 1306 4927 1362 4936
rect 1216 4616 1268 4622
rect 1216 4558 1268 4564
rect 388 4004 440 4010
rect 388 3946 440 3952
rect 400 480 428 3946
rect 1320 3754 1348 4927
rect 1412 4146 1440 5170
rect 1504 4690 1532 8434
rect 1596 5250 1624 13330
rect 1688 12782 1716 13738
rect 1858 13560 1914 13569
rect 1858 13495 1914 13504
rect 1872 13462 1900 13495
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 2056 13394 2084 14418
rect 2792 13938 2820 14447
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2240 13394 2268 13670
rect 2884 13530 2912 15127
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 1950 13152 2006 13161
rect 1950 13087 2006 13096
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1688 5409 1716 12718
rect 1780 6866 1808 12718
rect 1964 11286 1992 13087
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11354 2084 12174
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1858 9616 1914 9625
rect 1858 9551 1914 9560
rect 1872 8498 1900 9551
rect 1964 9042 1992 11086
rect 2148 10810 2176 12242
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2240 10690 2268 13330
rect 2976 12986 3004 16079
rect 3238 15872 3294 15881
rect 3238 15807 3294 15816
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3068 13870 3096 14350
rect 3252 14074 3280 15807
rect 3436 14074 3464 16487
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3804 13954 3832 15399
rect 4080 14414 4108 16759
rect 4986 16520 5042 17000
rect 8298 16520 8354 17000
rect 11610 16520 11666 17000
rect 14922 16520 14978 17000
rect 15290 16824 15346 16833
rect 15290 16759 15346 16768
rect 5000 14618 5028 16520
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 5184 14278 5212 14418
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3804 13926 4016 13954
rect 3988 13870 4016 13926
rect 3056 13864 3108 13870
rect 3054 13832 3056 13841
rect 3976 13864 4028 13870
rect 3108 13832 3110 13841
rect 3976 13806 4028 13812
rect 3054 13767 3110 13776
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 4528 12912 4580 12918
rect 3330 12880 3386 12889
rect 2688 12844 2740 12850
rect 4528 12854 4580 12860
rect 3330 12815 3386 12824
rect 4068 12844 4120 12850
rect 2688 12786 2740 12792
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2056 10662 2268 10690
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7546 1900 8230
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6458 1808 6802
rect 2056 6610 2084 10662
rect 2134 9480 2190 9489
rect 2134 9415 2190 9424
rect 2148 7342 2176 9415
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2240 8362 2268 8434
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2240 7818 2268 8298
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2240 7410 2268 7754
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 1872 6582 2084 6610
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1780 5953 1808 6190
rect 1766 5944 1822 5953
rect 1766 5879 1822 5888
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1674 5400 1730 5409
rect 1674 5335 1730 5344
rect 1596 5222 1716 5250
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1320 3738 1440 3754
rect 1320 3732 1452 3738
rect 1320 3726 1400 3732
rect 1400 3674 1452 3680
rect 1596 2825 1624 4422
rect 1688 3641 1716 5222
rect 1674 3632 1730 3641
rect 1674 3567 1730 3576
rect 1582 2816 1638 2825
rect 1582 2751 1638 2760
rect 1780 2650 1808 5714
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1872 2106 1900 6582
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1964 5030 1992 6394
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5166 2084 6054
rect 2148 5250 2176 6258
rect 2240 6202 2268 7346
rect 2332 6322 2360 12582
rect 2608 12442 2636 12582
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2424 11626 2452 12174
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 10198 2452 11562
rect 2516 10554 2544 12310
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 11150 2636 11630
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2608 10674 2636 11086
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2516 10526 2636 10554
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2424 8498 2452 9454
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2608 7936 2636 10526
rect 2700 9994 2728 12786
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2962 12336 3018 12345
rect 2962 12271 3018 12280
rect 2778 11656 2834 11665
rect 2778 11591 2834 11600
rect 2792 11354 2820 11591
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2700 9450 2728 9930
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8362 2728 8774
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2516 7908 2636 7936
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 7313 2452 7822
rect 2410 7304 2466 7313
rect 2410 7239 2466 7248
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2516 6254 2544 7908
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2504 6248 2556 6254
rect 2240 6174 2360 6202
rect 2504 6190 2556 6196
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2332 6066 2360 6174
rect 2240 5914 2268 6054
rect 2332 6038 2544 6066
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2148 5222 2452 5250
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2136 5092 2188 5098
rect 2136 5034 2188 5040
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2650 2084 2790
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1860 2100 1912 2106
rect 1860 2042 1912 2048
rect 1216 2032 1268 2038
rect 1216 1974 1268 1980
rect 1228 480 1256 1974
rect 2148 480 2176 5034
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 3040 2268 4966
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2332 3738 2360 4626
rect 2424 3738 2452 5222
rect 2516 4622 2544 6038
rect 2608 4826 2636 7142
rect 2792 5817 2820 10678
rect 2884 10606 2912 11086
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2884 7041 2912 10095
rect 2870 7032 2926 7041
rect 2870 6967 2926 6976
rect 2870 6896 2926 6905
rect 2976 6882 3004 12271
rect 3068 10810 3096 12582
rect 3252 12345 3280 12650
rect 3238 12336 3294 12345
rect 3238 12271 3240 12280
rect 3292 12271 3294 12280
rect 3240 12242 3292 12248
rect 3344 12186 3372 12815
rect 4068 12786 4120 12792
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3620 12209 3648 12582
rect 3712 12345 3740 12582
rect 4080 12481 4108 12786
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4066 12472 4122 12481
rect 4066 12407 4122 12416
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3252 12158 3372 12186
rect 3606 12200 3662 12209
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3054 10160 3110 10169
rect 3054 10095 3056 10104
rect 3108 10095 3110 10104
rect 3056 10066 3108 10072
rect 3054 10024 3110 10033
rect 3054 9959 3110 9968
rect 3068 9450 3096 9959
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3160 9382 3188 12106
rect 3252 10062 3280 12158
rect 3606 12135 3662 12144
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2926 6854 3004 6882
rect 2870 6831 2926 6840
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2688 5704 2740 5710
rect 2884 5681 2912 6831
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2688 5646 2740 5652
rect 2870 5672 2926 5681
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2320 3052 2372 3058
rect 2240 3012 2320 3040
rect 2320 2994 2372 3000
rect 2332 2446 2360 2994
rect 2424 2922 2452 3538
rect 2516 3466 2544 4422
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2608 2394 2636 3470
rect 2700 3194 2728 5646
rect 2870 5607 2926 5616
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2792 4282 2820 5034
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3058 2820 4218
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2792 2650 2820 2858
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2780 2440 2832 2446
rect 2608 2388 2780 2394
rect 2608 2382 2832 2388
rect 2608 2366 2820 2382
rect 2884 2145 2912 5510
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 2976 1873 3004 6122
rect 3068 4185 3096 8774
rect 3160 8362 3188 8910
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2962 1864 3018 1873
rect 2962 1799 3018 1808
rect 3068 480 3096 3606
rect 3160 513 3188 8026
rect 3252 5273 3280 9862
rect 3238 5264 3294 5273
rect 3238 5199 3294 5208
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3252 4690 3280 5034
rect 3344 4826 3372 12038
rect 3620 11830 3648 12135
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3608 11824 3660 11830
rect 3712 11801 3740 12038
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3608 11766 3660 11772
rect 3698 11792 3754 11801
rect 3424 11756 3476 11762
rect 3698 11727 3754 11736
rect 4344 11756 4396 11762
rect 3424 11698 3476 11704
rect 4344 11698 4396 11704
rect 3436 11558 3464 11698
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3436 10742 3464 11494
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3528 10674 3556 11494
rect 4080 11218 4108 11562
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 9722 3464 10406
rect 3620 10266 3648 11086
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10441 3832 10950
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4264 10810 4292 11630
rect 4356 11354 4384 11698
rect 4448 11370 4476 12582
rect 4540 12442 4568 12854
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12442 4752 12582
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4344 11348 4396 11354
rect 4448 11342 4568 11370
rect 4344 11290 4396 11296
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4356 10606 4384 11290
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 3976 10464 4028 10470
rect 3790 10432 3846 10441
rect 3976 10406 4028 10412
rect 3790 10367 3846 10376
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3436 8090 3464 9046
rect 3528 8401 3556 9998
rect 3620 9518 3648 10202
rect 3712 9897 3740 10202
rect 3884 10056 3936 10062
rect 3804 10004 3884 10010
rect 3988 10033 4016 10406
rect 4356 10112 4384 10542
rect 4347 10084 4384 10112
rect 4347 10033 4375 10084
rect 3804 9998 3936 10004
rect 3974 10024 4030 10033
rect 3804 9982 3924 9998
rect 3698 9888 3754 9897
rect 3698 9823 3754 9832
rect 3804 9586 3832 9982
rect 3974 9959 4030 9968
rect 4342 10024 4398 10033
rect 4342 9959 4398 9968
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4342 9752 4398 9761
rect 4342 9687 4398 9696
rect 4436 9716 4488 9722
rect 4356 9586 4384 9687
rect 4436 9658 4488 9664
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 3608 9512 3660 9518
rect 4448 9466 4476 9658
rect 3608 9454 3660 9460
rect 3620 9042 3648 9454
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 4356 9438 4476 9466
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8634 3648 8774
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3528 7954 3556 8327
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 7410 3464 7822
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 6186 3464 6666
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3436 5710 3464 6122
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3240 4684 3292 4690
rect 3292 4644 3372 4672
rect 3240 4626 3292 4632
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3252 3738 3280 4014
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3252 2446 3280 2994
rect 3344 2990 3372 4644
rect 3436 3233 3464 5510
rect 3528 5370 3556 6870
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3528 4593 3556 5170
rect 3514 4584 3570 4593
rect 3514 4519 3570 4528
rect 3514 3496 3570 3505
rect 3514 3431 3516 3440
rect 3568 3431 3570 3440
rect 3516 3402 3568 3408
rect 3422 3224 3478 3233
rect 3422 3159 3478 3168
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3436 2514 3464 3023
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3620 1465 3648 6598
rect 3712 5692 3740 9318
rect 3988 8945 4016 9386
rect 4356 9042 4384 9438
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 3974 8936 4030 8945
rect 3974 8871 4030 8880
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 4356 8634 4384 8978
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 7857 4108 8366
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7410 3832 7686
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 6905 3924 7278
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4068 6248 4120 6254
rect 4066 6216 4068 6225
rect 4120 6216 4122 6225
rect 4066 6151 4122 6160
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5710 4108 6054
rect 4160 5840 4212 5846
rect 4158 5808 4160 5817
rect 4212 5808 4214 5817
rect 4158 5743 4214 5752
rect 4068 5704 4120 5710
rect 3712 5664 3832 5692
rect 3698 5536 3754 5545
rect 3698 5471 3754 5480
rect 3712 5370 3740 5471
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 3712 3670 3740 5199
rect 3804 4622 3832 5664
rect 4068 5646 4120 5652
rect 4264 5658 4292 8230
rect 4448 7886 4476 8298
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 7410 4384 7754
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4448 6798 4476 7346
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4356 5846 4384 6394
rect 4448 6118 4476 6734
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4264 5630 4384 5658
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4158 5128 4214 5137
rect 4158 5063 4214 5072
rect 4172 4622 4200 5063
rect 4264 4865 4292 5510
rect 4356 5234 4384 5630
rect 4448 5234 4476 6054
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4250 4856 4306 4865
rect 4250 4791 4306 4800
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4160 4616 4212 4622
rect 4264 4593 4292 4694
rect 4356 4690 4384 4966
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4160 4558 4212 4564
rect 4250 4584 4306 4593
rect 4250 4519 4306 4528
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2582 3740 2790
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 3606 1456 3662 1465
rect 3804 1442 3832 3878
rect 4080 3602 4108 4111
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4264 2922 4292 4519
rect 4448 3942 4476 5034
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4540 3738 4568 11342
rect 4632 6866 4660 12174
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10674 4752 11154
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4724 10441 4752 10610
rect 4710 10432 4766 10441
rect 4710 10367 4766 10376
rect 4724 10062 4752 10367
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9217 4752 9862
rect 4710 9208 4766 9217
rect 4710 9143 4766 9152
rect 4816 8838 4844 12174
rect 4908 9518 4936 12786
rect 5184 11801 5212 14214
rect 8312 13938 8340 16520
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 13530 5764 13670
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5724 13320 5776 13326
rect 6380 13274 6408 13874
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7300 13530 7328 13806
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 5724 13262 5776 13268
rect 5736 12986 5764 13262
rect 6288 13258 6408 13274
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6276 13252 6408 13258
rect 6328 13246 6408 13252
rect 6276 13194 6328 13200
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5170 11792 5226 11801
rect 5170 11727 5226 11736
rect 5276 11642 5304 12378
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5092 11614 5304 11642
rect 4986 11248 5042 11257
rect 4986 11183 5042 11192
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 9178 4936 9454
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4894 8800 4950 8809
rect 4894 8735 4950 8744
rect 4908 8498 4936 8735
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4724 8072 4752 8434
rect 4804 8424 4856 8430
rect 4802 8392 4804 8401
rect 4856 8392 4858 8401
rect 4802 8327 4858 8336
rect 4724 8044 4844 8072
rect 4710 7984 4766 7993
rect 4710 7919 4766 7928
rect 4724 7886 4752 7919
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4816 6361 4844 8044
rect 4802 6352 4858 6361
rect 4802 6287 4858 6296
rect 4908 6236 4936 8434
rect 5000 8294 5028 11183
rect 5092 10146 5120 11614
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 10810 5212 11494
rect 5262 11248 5318 11257
rect 5262 11183 5264 11192
rect 5316 11183 5318 11192
rect 5264 11154 5316 11160
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5170 10704 5226 10713
rect 5170 10639 5226 10648
rect 5184 10470 5212 10639
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5092 10118 5212 10146
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5092 8022 5120 9998
rect 5184 8090 5212 10118
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5276 7954 5304 11018
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4724 6208 4936 6236
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4632 4010 4660 4558
rect 4724 4185 4752 6208
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4816 5846 4844 6054
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4804 5160 4856 5166
rect 4908 5148 4936 6054
rect 4986 5536 5042 5545
rect 5092 5522 5120 7754
rect 5092 5494 5212 5522
rect 4986 5471 5042 5480
rect 4856 5120 4936 5148
rect 4804 5102 4856 5108
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4710 4176 4766 4185
rect 4710 4111 4766 4120
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4356 2650 4384 3334
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4066 2544 4122 2553
rect 4632 2514 4660 3334
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4724 2650 4752 2790
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4066 2479 4122 2488
rect 4620 2508 4672 2514
rect 4080 2378 4108 2479
rect 4620 2450 4672 2456
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4816 2310 4844 4490
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3804 1414 4016 1442
rect 3606 1391 3662 1400
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3528 1193 3556 1294
rect 3514 1184 3570 1193
rect 3514 1119 3570 1128
rect 3424 604 3476 610
rect 3424 546 3476 552
rect 3146 504 3202 513
rect 386 0 442 480
rect 1214 0 1270 480
rect 2134 0 2190 480
rect 3054 0 3110 480
rect 3146 439 3202 448
rect 3436 241 3464 546
rect 3988 480 4016 1414
rect 4908 480 4936 3470
rect 5000 3126 5028 5471
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5092 3670 5120 4422
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5184 2961 5212 5494
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5276 4826 5304 5034
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3534 5304 3878
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 3058 5304 3470
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5170 2952 5226 2961
rect 5170 2887 5226 2896
rect 5368 2650 5396 12242
rect 5538 11792 5594 11801
rect 5538 11727 5594 11736
rect 5552 11098 5580 11727
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5460 11070 5580 11098
rect 5460 7818 5488 11070
rect 5644 10810 5672 11630
rect 5736 11354 5764 12718
rect 5906 12336 5962 12345
rect 5906 12271 5962 12280
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5736 10606 5764 10746
rect 5724 10600 5776 10606
rect 5552 10560 5724 10588
rect 5552 9081 5580 10560
rect 5724 10542 5776 10548
rect 5828 10282 5856 11290
rect 5920 10713 5948 12271
rect 5998 12200 6054 12209
rect 5998 12135 6054 12144
rect 5906 10704 5962 10713
rect 5906 10639 5962 10648
rect 6012 10470 6040 12135
rect 6104 11393 6132 13126
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12442 6224 12582
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6090 11384 6146 11393
rect 6090 11319 6146 11328
rect 6196 11150 6224 12174
rect 6288 11898 6316 13194
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6380 11694 6408 12582
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6472 12209 6500 12378
rect 6656 12374 6684 13262
rect 6840 12986 6868 13330
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 7208 12918 7236 13330
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 12368 6696 12374
rect 6748 12345 6776 12650
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6644 12310 6696 12316
rect 6734 12336 6790 12345
rect 6552 12300 6604 12306
rect 6734 12271 6790 12280
rect 6552 12242 6604 12248
rect 6458 12200 6514 12209
rect 6458 12135 6514 12144
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6380 11286 6408 11630
rect 6458 11384 6514 11393
rect 6458 11319 6514 11328
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6000 10464 6052 10470
rect 6104 10441 6132 10610
rect 6000 10406 6052 10412
rect 6090 10432 6146 10441
rect 5644 10254 5856 10282
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8498 5580 8910
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 7954 5580 8434
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 6322 5488 7210
rect 5552 7002 5580 7686
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6882 5672 10254
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5722 10024 5778 10033
rect 5722 9959 5724 9968
rect 5776 9959 5778 9968
rect 5724 9930 5776 9936
rect 5736 9500 5764 9930
rect 5828 9654 5856 10134
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5736 9472 5856 9500
rect 5828 8820 5856 9472
rect 6012 9081 6040 10406
rect 6090 10367 6146 10376
rect 5998 9072 6054 9081
rect 5998 9007 6054 9016
rect 6000 8832 6052 8838
rect 5828 8792 5948 8820
rect 5920 8276 5948 8792
rect 6000 8774 6052 8780
rect 6012 8430 6040 8774
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5920 8248 6040 8276
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5736 7478 5764 7822
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5736 7206 5764 7414
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5552 6854 5672 6882
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5166 5488 5510
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5460 4554 5488 5102
rect 5552 5030 5580 6854
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5538 4720 5594 4729
rect 5538 4655 5594 4664
rect 5552 4622 5580 4655
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 3534 5580 4422
rect 5644 4026 5672 6598
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5914 5764 6054
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5828 5098 5856 7482
rect 6012 7426 6040 8248
rect 6104 7546 6132 10367
rect 6196 9722 6224 11086
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6288 9654 6316 10474
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6012 7398 6132 7426
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6322 5948 6598
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 6104 6100 6132 7398
rect 6196 7206 6224 9454
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6274 8528 6330 8537
rect 6380 8498 6408 9386
rect 6274 8463 6330 8472
rect 6368 8492 6420 8498
rect 6288 7274 6316 8463
rect 6368 8434 6420 8440
rect 6472 7834 6500 11319
rect 6564 10810 6592 12242
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6656 10198 6684 12174
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6840 11694 6868 11834
rect 6828 11688 6880 11694
rect 6748 11648 6828 11676
rect 6748 10810 6776 11648
rect 6828 11630 6880 11636
rect 7300 11626 7328 12786
rect 7392 12442 7420 13670
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6748 10674 6776 10746
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6656 9586 6684 10134
rect 6748 10130 6776 10610
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7300 10266 7328 11562
rect 7484 11121 7512 13670
rect 7576 13326 7604 13874
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12850 7604 13262
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7470 11112 7526 11121
rect 7470 11047 7526 11056
rect 7576 10996 7604 12650
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7484 10968 7604 10996
rect 7484 10305 7512 10968
rect 7668 10849 7696 11154
rect 7654 10840 7710 10849
rect 7654 10775 7710 10784
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7470 10296 7526 10305
rect 7288 10260 7340 10266
rect 7470 10231 7526 10240
rect 7288 10202 7340 10208
rect 7484 10198 7512 10231
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9586 6776 10066
rect 7472 10056 7524 10062
rect 6826 10024 6882 10033
rect 7472 9998 7524 10004
rect 6826 9959 6828 9968
rect 6880 9959 6882 9968
rect 6828 9930 6880 9936
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6564 9042 6592 9454
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6550 8800 6606 8809
rect 6550 8735 6606 8744
rect 6564 8537 6592 8735
rect 6550 8528 6606 8537
rect 6550 8463 6606 8472
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6564 7886 6592 8327
rect 6656 7886 6684 9386
rect 6748 9042 6776 9522
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7392 9178 7420 9386
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7378 8936 7434 8945
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 8090 6776 8570
rect 7024 8498 7052 8910
rect 7378 8871 7434 8880
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6826 8392 6882 8401
rect 6826 8327 6828 8336
rect 6880 8327 6882 8336
rect 6828 8298 6880 8304
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6380 7806 6500 7834
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 6254 6224 7142
rect 6276 6792 6328 6798
rect 6274 6760 6276 6769
rect 6328 6760 6330 6769
rect 6274 6695 6330 6704
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6104 6072 6316 6100
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5736 4457 5764 4626
rect 5722 4448 5778 4457
rect 5722 4383 5778 4392
rect 5828 4162 5856 4694
rect 5920 4690 5948 5782
rect 6184 5704 6236 5710
rect 6090 5672 6146 5681
rect 6184 5646 6236 5652
rect 6090 5607 6146 5616
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5920 4321 5948 4626
rect 5906 4312 5962 4321
rect 5906 4247 5962 4256
rect 5828 4134 5948 4162
rect 5816 4072 5868 4078
rect 5644 3998 5764 4026
rect 5816 4014 5868 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3738 5672 3878
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5460 2582 5488 3062
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5552 2446 5580 3334
rect 5736 2650 5764 3998
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5828 480 5856 4014
rect 5920 3777 5948 4134
rect 5906 3768 5962 3777
rect 5906 3703 5962 3712
rect 5906 3496 5962 3505
rect 5906 3431 5962 3440
rect 5920 2514 5948 3431
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6012 610 6040 5510
rect 6104 5166 6132 5607
rect 6196 5370 6224 5646
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6288 5250 6316 6072
rect 6196 5222 6316 5250
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6104 3194 6132 5102
rect 6196 4049 6224 5222
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4146 6316 4966
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6182 4040 6238 4049
rect 6182 3975 6238 3984
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6196 3058 6224 3878
rect 6288 3058 6316 4082
rect 6380 3210 6408 7806
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6322 6500 6598
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6472 5710 6500 6258
rect 6564 5914 6592 7142
rect 6656 6497 6684 7686
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 6642 6488 6698 6497
rect 6748 6458 6776 6695
rect 6642 6423 6698 6432
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6642 5944 6698 5953
rect 6552 5908 6604 5914
rect 6642 5879 6698 5888
rect 6552 5850 6604 5856
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6564 5545 6592 5714
rect 6550 5536 6606 5545
rect 6550 5471 6606 5480
rect 6460 5024 6512 5030
rect 6458 4992 6460 5001
rect 6512 4992 6514 5001
rect 6458 4927 6514 4936
rect 6472 4826 6500 4927
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 3398 6500 4626
rect 6656 4282 6684 5879
rect 6748 5710 6776 6394
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 4486 6776 5646
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6550 4176 6606 4185
rect 6656 4146 6684 4218
rect 6550 4111 6606 4120
rect 6644 4140 6696 4146
rect 6564 4010 6592 4111
rect 6644 4082 6696 4088
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6380 3182 6500 3210
rect 6366 3088 6422 3097
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6276 3052 6328 3058
rect 6366 3023 6422 3032
rect 6276 2994 6328 3000
rect 6104 2922 6316 2938
rect 6092 2916 6328 2922
rect 6144 2910 6276 2916
rect 6092 2858 6144 2864
rect 6276 2858 6328 2864
rect 6380 2854 6408 3023
rect 6472 2990 6500 3182
rect 6564 3058 6592 3946
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6656 1358 6684 3946
rect 6748 3738 6776 4422
rect 7010 4176 7066 4185
rect 7010 4111 7066 4120
rect 7024 4078 7052 4111
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 3194 7236 3334
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6000 604 6052 610
rect 6000 546 6052 552
rect 6748 480 6776 2858
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7300 2582 7328 8570
rect 7392 7886 7420 8871
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 6866 7420 7346
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6322 7420 6802
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 5234 7420 6258
rect 7484 6254 7512 9998
rect 7576 8090 7604 10406
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7668 9382 7696 10134
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 8498 7696 9318
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7760 8242 7788 13806
rect 11624 13802 11652 16520
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 14278 14512 14334 14521
rect 14278 14447 14334 14456
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11801 7880 12038
rect 7838 11792 7894 11801
rect 7838 11727 7894 11736
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10538 7880 10950
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7668 8214 7788 8242
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7576 7954 7604 8026
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7562 7304 7618 7313
rect 7562 7239 7618 7248
rect 7576 6254 7604 7239
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 3126 7420 4626
rect 7470 4312 7526 4321
rect 7470 4247 7526 4256
rect 7484 3602 7512 4247
rect 7576 3942 7604 5850
rect 7668 4049 7696 8214
rect 7852 7954 7880 8978
rect 7944 8838 7972 12582
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 8036 8430 8064 12038
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8128 11082 8156 11562
rect 8220 11558 8248 13398
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8128 8294 8156 11018
rect 8220 10606 8248 11494
rect 8208 10600 8260 10606
rect 8312 10577 8340 12582
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8208 10542 8260 10548
rect 8298 10568 8354 10577
rect 8298 10503 8354 10512
rect 8312 10266 8340 10503
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8206 9072 8262 9081
rect 8206 9007 8262 9016
rect 8220 8401 8248 9007
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 8206 8392 8262 8401
rect 8206 8327 8262 8336
rect 8312 8294 8340 8871
rect 8404 8430 8432 12174
rect 8496 11354 8524 13126
rect 8588 12374 8616 13194
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11665 8616 12038
rect 8574 11656 8630 11665
rect 8574 11591 8630 11600
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8496 11121 8524 11154
rect 8668 11144 8720 11150
rect 8482 11112 8538 11121
rect 8668 11086 8720 11092
rect 8482 11047 8538 11056
rect 8482 10296 8538 10305
rect 8482 10231 8538 10240
rect 8496 10198 8524 10231
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8680 9654 8708 11086
rect 8772 10810 8800 13194
rect 8864 12782 8892 13262
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 9048 12714 9076 13330
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8772 9110 8800 10746
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8864 8945 8892 12582
rect 8944 12368 8996 12374
rect 8942 12336 8944 12345
rect 8996 12336 8998 12345
rect 8942 12271 8998 12280
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 12209 9076 12242
rect 9140 12238 9168 12786
rect 9784 12730 9812 13330
rect 10968 13320 11020 13326
rect 10966 13288 10968 13297
rect 11020 13288 11022 13297
rect 10966 13223 11022 13232
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 9692 12702 9812 12730
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10140 12708 10192 12714
rect 9128 12232 9180 12238
rect 9034 12200 9090 12209
rect 9128 12174 9180 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9034 12135 9090 12144
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8956 10810 8984 11290
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9048 9926 9076 10202
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9036 9512 9088 9518
rect 9140 9500 9168 12174
rect 9232 11626 9260 12174
rect 9692 11778 9720 12702
rect 10140 12650 10192 12656
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9508 11750 9720 11778
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11150 9260 11562
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 9586 9352 10610
rect 9508 9625 9536 11750
rect 9680 11620 9732 11626
rect 9600 11580 9680 11608
rect 9600 10674 9628 11580
rect 9680 11562 9732 11568
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9494 9616 9550 9625
rect 9312 9580 9364 9586
rect 9494 9551 9550 9560
rect 9312 9522 9364 9528
rect 9088 9472 9168 9500
rect 9036 9454 9088 9460
rect 9140 9178 9168 9472
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8850 8936 8906 8945
rect 8850 8871 8906 8880
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8634 8984 8842
rect 9692 8650 9720 11290
rect 9784 9450 9812 12582
rect 9968 12306 9996 12582
rect 10152 12345 10180 12650
rect 10138 12336 10194 12345
rect 9956 12300 10008 12306
rect 10138 12271 10194 12280
rect 9956 12242 10008 12248
rect 9968 12209 9996 12242
rect 9954 12200 10010 12209
rect 9954 12135 10010 12144
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10140 11688 10192 11694
rect 10138 11656 10140 11665
rect 10192 11656 10194 11665
rect 10138 11591 10194 11600
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9864 11280 9916 11286
rect 9862 11248 9864 11257
rect 9916 11248 9918 11257
rect 9862 11183 9918 11192
rect 10152 11132 10180 11494
rect 10244 11234 10272 12718
rect 10336 12442 10364 12786
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11354 10364 12038
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10244 11206 10364 11234
rect 10232 11144 10284 11150
rect 10152 11104 10232 11132
rect 10232 11086 10284 11092
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10060 10198 10088 10639
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9956 9512 10008 9518
rect 10244 9500 10272 11086
rect 10336 10033 10364 11206
rect 10322 10024 10378 10033
rect 10322 9959 10378 9968
rect 10008 9472 10272 9500
rect 9956 9454 10008 9460
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9876 9042 9904 9386
rect 10046 9208 10102 9217
rect 10046 9143 10102 9152
rect 10060 9042 10088 9143
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9508 8622 9720 8650
rect 9784 8634 9812 8842
rect 10060 8820 10088 8978
rect 10232 8968 10284 8974
rect 10336 8956 10364 9959
rect 10428 9178 10456 12650
rect 10520 11121 10548 12786
rect 10796 12306 10824 12922
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10506 11112 10562 11121
rect 10506 11047 10562 11056
rect 10520 10606 10548 11047
rect 10612 10810 10640 11591
rect 10704 11354 10732 12242
rect 10782 11928 10838 11937
rect 10782 11863 10784 11872
rect 10836 11863 10838 11872
rect 10784 11834 10836 11840
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10600 10804 10652 10810
rect 10652 10764 10732 10792
rect 10600 10746 10652 10752
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 10062 10548 10542
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 10130 10640 10474
rect 10704 10266 10732 10764
rect 10692 10260 10744 10266
rect 10744 10220 10824 10248
rect 10692 10202 10744 10208
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10506 9888 10562 9897
rect 10506 9823 10562 9832
rect 10520 9217 10548 9823
rect 10598 9752 10654 9761
rect 10704 9738 10732 9787
rect 10796 9738 10824 10220
rect 10704 9722 10824 9738
rect 10598 9687 10654 9696
rect 10692 9716 10824 9722
rect 10612 9489 10640 9687
rect 10744 9710 10824 9716
rect 10692 9658 10744 9664
rect 10598 9480 10654 9489
rect 10598 9415 10654 9424
rect 10506 9208 10562 9217
rect 10416 9172 10468 9178
rect 10506 9143 10562 9152
rect 10416 9114 10468 9120
rect 10284 8928 10364 8956
rect 10232 8910 10284 8916
rect 10060 8792 10272 8820
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 9772 8628 9824 8634
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8760 8424 8812 8430
rect 9508 8412 9536 8622
rect 9772 8570 9824 8576
rect 9588 8560 9640 8566
rect 9640 8508 9812 8514
rect 9588 8502 9812 8508
rect 9600 8486 9812 8502
rect 9508 8384 9720 8412
rect 8760 8366 8812 8372
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8128 7954 8156 8230
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7177 7788 7822
rect 7840 7336 7892 7342
rect 8208 7336 8260 7342
rect 7840 7278 7892 7284
rect 7746 7168 7802 7177
rect 7746 7103 7802 7112
rect 7760 5914 7788 7103
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7746 4720 7802 4729
rect 7746 4655 7802 4664
rect 7654 4040 7710 4049
rect 7654 3975 7710 3984
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7576 2825 7604 3878
rect 7760 3058 7788 4655
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7852 2650 7880 7278
rect 7944 7262 8156 7290
rect 8208 7278 8260 7284
rect 7944 7206 7972 7262
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7944 5166 7972 6938
rect 8036 5302 8064 7142
rect 8128 7018 8156 7262
rect 8220 7206 8248 7278
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8312 7018 8340 8230
rect 8128 6990 8340 7018
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 6458 8156 6734
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5778 8156 6190
rect 8220 5914 8248 6258
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7932 5160 7984 5166
rect 8128 5114 8156 5578
rect 7932 5102 7984 5108
rect 8036 5086 8156 5114
rect 7932 4616 7984 4622
rect 8036 4604 8064 5086
rect 7984 4576 8064 4604
rect 7932 4558 7984 4564
rect 8024 4480 8076 4486
rect 7930 4448 7986 4457
rect 8076 4428 8156 4434
rect 8024 4422 8156 4428
rect 8036 4406 8156 4422
rect 7930 4383 7986 4392
rect 7944 2990 7972 4383
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 8036 2854 8064 4218
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7576 480 7604 2382
rect 8128 785 8156 4406
rect 8220 3058 8248 5646
rect 8312 4554 8340 6990
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8588 6361 8616 6938
rect 8574 6352 8630 6361
rect 8574 6287 8630 6296
rect 8588 6254 8616 6287
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5817 8432 6054
rect 8496 5914 8524 6122
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8390 5808 8446 5817
rect 8390 5743 8446 5752
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8404 5234 8432 5578
rect 8482 5536 8538 5545
rect 8482 5471 8538 5480
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8496 5030 8524 5471
rect 8772 5030 8800 8366
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 7274 8892 8230
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8956 7342 8984 7414
rect 9048 7342 9076 7482
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 9048 5778 9076 7278
rect 9232 6934 9260 7686
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9586 6896 9642 6905
rect 9692 6882 9720 8384
rect 9784 7426 9812 8486
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9968 8129 9996 8434
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10152 8265 10180 8366
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 9954 8120 10010 8129
rect 9954 8055 10010 8064
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10244 7546 10272 8792
rect 10336 7886 10364 8928
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9784 7398 9904 7426
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9784 7002 9812 7210
rect 9876 7002 9904 7398
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9692 6854 10272 6882
rect 10428 6866 10456 8871
rect 10506 8664 10562 8673
rect 10506 8599 10562 8608
rect 10520 8566 10548 8599
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10612 8106 10640 9415
rect 10704 8974 10732 9658
rect 10692 8968 10744 8974
rect 10744 8928 10824 8956
rect 10692 8910 10744 8916
rect 10612 8078 10732 8106
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10520 7546 10548 7890
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 9586 6831 9642 6840
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6254 9536 6598
rect 9600 6254 9628 6831
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8496 4264 8524 4966
rect 8772 4826 8800 4966
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8576 4276 8628 4282
rect 8496 4236 8576 4264
rect 8576 4218 8628 4224
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 8312 4078 8340 4111
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8312 3058 8340 4014
rect 8404 3738 8432 4014
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8956 3194 8984 4626
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8772 2650 8800 3062
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8114 776 8170 785
rect 8114 711 8170 720
rect 8496 480 8524 2382
rect 9048 2378 9076 4762
rect 9232 4706 9260 5850
rect 9508 5234 9536 6190
rect 9680 5704 9732 5710
rect 9784 5692 9812 6666
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5778 9996 6054
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9732 5664 9812 5692
rect 9680 5646 9732 5652
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9600 5522 9628 5578
rect 9600 5494 9720 5522
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9692 5098 9720 5494
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9140 4678 9260 4706
rect 9140 3670 9168 4678
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9586 4584 9642 4593
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9140 3058 9168 3606
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9232 2038 9260 4014
rect 9324 4010 9352 4558
rect 9586 4519 9588 4528
rect 9640 4519 9642 4528
rect 9588 4490 9640 4496
rect 9784 4486 9812 5664
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 10046 4720 10102 4729
rect 10046 4655 10102 4664
rect 10060 4554 10088 4655
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9324 3398 9352 3946
rect 9692 3738 9720 4422
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3058 9352 3334
rect 9600 3194 9628 3538
rect 9784 3194 9812 4218
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3602 10180 3946
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9416 480 9444 2926
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9508 2446 9536 2858
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 9876 2582 9904 2790
rect 10060 2650 10088 2790
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 10244 2514 10272 6854
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6390 10364 6734
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10336 4758 10364 6122
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4146 10364 4422
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10428 3534 10456 5238
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10520 3194 10548 7482
rect 10704 5778 10732 8078
rect 10796 8022 10824 8928
rect 10784 8016 10836 8022
rect 10888 7993 10916 12582
rect 10980 9654 11008 13126
rect 11150 12880 11206 12889
rect 11150 12815 11206 12824
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 9110 11008 9590
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11072 8838 11100 12582
rect 11164 9994 11192 12815
rect 11612 12368 11664 12374
rect 11426 12336 11482 12345
rect 11664 12328 11744 12356
rect 11612 12310 11664 12316
rect 11426 12271 11482 12280
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11256 11898 11284 12135
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11242 11792 11298 11801
rect 11242 11727 11298 11736
rect 11256 11694 11284 11727
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11354 11284 11494
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9625 11284 9862
rect 11242 9616 11298 9625
rect 11242 9551 11298 9560
rect 11150 9072 11206 9081
rect 11150 9007 11206 9016
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10784 7958 10836 7964
rect 10874 7984 10930 7993
rect 10874 7919 10930 7928
rect 10980 7886 11008 8434
rect 11164 8430 11192 9007
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10612 3505 10640 3606
rect 10598 3496 10654 3505
rect 10598 3431 10654 3440
rect 10598 3224 10654 3233
rect 10508 3188 10560 3194
rect 10598 3159 10654 3168
rect 10508 3130 10560 3136
rect 10506 2816 10562 2825
rect 10506 2751 10562 2760
rect 10520 2650 10548 2751
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10612 2514 10640 3159
rect 10704 3126 10732 5578
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10796 2854 10824 7822
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10888 4690 10916 7754
rect 11072 7546 11100 8298
rect 11256 8294 11284 8366
rect 11244 8288 11296 8294
rect 11150 8256 11206 8265
rect 11244 8230 11296 8236
rect 11336 8288 11388 8294
rect 11440 8265 11468 12271
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11532 11898 11560 12174
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11150 11560 11562
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10810 11560 11086
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11336 8230 11388 8236
rect 11426 8256 11482 8265
rect 11150 8191 11206 8200
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10966 6488 11022 6497
rect 11164 6458 11192 8191
rect 11256 7886 11284 8230
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11348 7732 11376 8230
rect 11426 8191 11482 8200
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11256 7704 11376 7732
rect 11256 7274 11284 7704
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11256 6458 11284 7210
rect 11336 7200 11388 7206
rect 11440 7188 11468 7958
rect 11532 7410 11560 10066
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11388 7160 11468 7188
rect 11336 7142 11388 7148
rect 10966 6423 10968 6432
rect 11020 6423 11022 6432
rect 11152 6452 11204 6458
rect 10968 6394 11020 6400
rect 11152 6394 11204 6400
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5166 11008 6190
rect 11624 6186 11652 12174
rect 11716 11665 11744 12328
rect 11808 12238 11836 14010
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11702 11656 11758 11665
rect 11900 11626 11928 12174
rect 12084 11762 12112 12786
rect 12360 12782 12388 13738
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 12532 12844 12584 12850
rect 12452 12804 12532 12832
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11702 11591 11758 11600
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11980 11076 12032 11082
rect 11900 11036 11980 11064
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10810 11744 10950
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 10130 11744 10542
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 8634 11744 9318
rect 11808 9058 11836 10406
rect 11900 9450 11928 11036
rect 11980 11018 12032 11024
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11808 9030 11928 9058
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11704 8288 11756 8294
rect 11702 8256 11704 8265
rect 11756 8256 11758 8265
rect 11702 8191 11758 8200
rect 11808 8090 11836 8910
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11900 7585 11928 9030
rect 11886 7576 11942 7585
rect 11886 7511 11942 7520
rect 11794 7440 11850 7449
rect 11704 7404 11756 7410
rect 11794 7375 11796 7384
rect 11704 7346 11756 7352
rect 11848 7375 11850 7384
rect 11796 7346 11848 7352
rect 11716 7002 11744 7346
rect 11900 7342 11928 7511
rect 11888 7336 11940 7342
rect 11794 7304 11850 7313
rect 11888 7278 11940 7284
rect 11794 7239 11850 7248
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11716 6322 11744 6938
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11808 6118 11836 7239
rect 11992 7206 12020 10095
rect 12084 9178 12112 11698
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 9466 12204 11630
rect 12254 11248 12310 11257
rect 12254 11183 12256 11192
rect 12308 11183 12310 11192
rect 12256 11154 12308 11160
rect 12268 10577 12296 11154
rect 12254 10568 12310 10577
rect 12254 10503 12310 10512
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12268 9625 12296 9658
rect 12254 9616 12310 9625
rect 12254 9551 12310 9560
rect 12176 9438 12296 9466
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 9178 12204 9318
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12070 8120 12126 8129
rect 12070 8055 12126 8064
rect 12084 7954 12112 8055
rect 12176 8022 12204 8230
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 12084 6730 12112 7890
rect 12268 7834 12296 9438
rect 12360 7993 12388 12038
rect 12346 7984 12402 7993
rect 12346 7919 12402 7928
rect 12176 7806 12296 7834
rect 12348 7812 12400 7818
rect 12176 7313 12204 7806
rect 12348 7754 12400 7760
rect 12256 7744 12308 7750
rect 12254 7712 12256 7721
rect 12308 7712 12310 7721
rect 12254 7647 12310 7656
rect 12162 7304 12218 7313
rect 12162 7239 12218 7248
rect 12164 7200 12216 7206
rect 12162 7168 12164 7177
rect 12216 7168 12218 7177
rect 12162 7103 12218 7112
rect 12360 6866 12388 7754
rect 12452 7478 12480 12804
rect 12532 12786 12584 12792
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 12714 11656 12770 11665
rect 12714 11591 12770 11600
rect 13358 11656 13414 11665
rect 13358 11591 13414 11600
rect 12532 11144 12584 11150
rect 12530 11112 12532 11121
rect 12584 11112 12586 11121
rect 12728 11082 12756 11591
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12530 11047 12586 11056
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12530 9752 12586 9761
rect 12530 9687 12532 9696
rect 12584 9687 12586 9696
rect 12532 9658 12584 9664
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 8838 12572 9454
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12636 8430 12664 10746
rect 13266 10704 13322 10713
rect 13266 10639 13322 10648
rect 13174 10568 13230 10577
rect 12716 10532 12768 10538
rect 13280 10538 13308 10639
rect 13174 10503 13230 10512
rect 13268 10532 13320 10538
rect 12716 10474 12768 10480
rect 12728 9926 12756 10474
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12820 10033 12848 10134
rect 12806 10024 12862 10033
rect 12806 9959 12862 9968
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9654 13032 9862
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12530 8256 12586 8265
rect 12530 8191 12586 8200
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10874 3088 10930 3097
rect 10874 3023 10876 3032
rect 10928 3023 10930 3032
rect 10876 2994 10928 3000
rect 10980 2990 11008 3878
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 11072 2514 11100 3334
rect 11164 2514 11192 4966
rect 11256 4570 11284 5034
rect 11348 4690 11376 5170
rect 11532 5166 11560 5510
rect 11900 5370 11928 5850
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11532 4826 11560 4966
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11336 4684 11388 4690
rect 11388 4644 11468 4672
rect 11336 4626 11388 4632
rect 11334 4584 11390 4593
rect 11256 4542 11334 4570
rect 11334 4519 11390 4528
rect 11348 3602 11376 4519
rect 11440 3618 11468 4644
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11532 3738 11560 4558
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11336 3596 11388 3602
rect 11440 3590 11560 3618
rect 11336 3538 11388 3544
rect 11532 3534 11560 3590
rect 11244 3528 11296 3534
rect 11428 3528 11480 3534
rect 11296 3476 11376 3482
rect 11244 3470 11376 3476
rect 11428 3470 11480 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11256 3454 11376 3470
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11256 2582 11284 2994
rect 11348 2990 11376 3454
rect 11440 3194 11468 3470
rect 11624 3398 11652 4490
rect 11716 3466 11744 4966
rect 11992 3738 12020 5646
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 12084 3126 12112 6666
rect 12164 6656 12216 6662
rect 12216 6616 12388 6644
rect 12164 6598 12216 6604
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 5098 12204 5646
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12176 4622 12204 5034
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12162 4040 12218 4049
rect 12162 3975 12218 3984
rect 12176 3942 12204 3975
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12268 3738 12296 6394
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 12360 2514 12388 6616
rect 12452 5642 12480 7278
rect 12544 7154 12572 8191
rect 12636 7750 12664 8366
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12636 7274 12664 7414
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12544 7126 12664 7154
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6254 12572 6598
rect 12636 6497 12664 7126
rect 12622 6488 12678 6497
rect 12622 6423 12678 6432
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12452 4622 12480 5102
rect 12544 5030 12572 5238
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12636 4842 12664 6423
rect 12544 4814 12664 4842
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12452 4146 12480 4558
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12438 3904 12494 3913
rect 12438 3839 12494 3848
rect 12452 2650 12480 3839
rect 12544 3738 12572 4814
rect 12728 4162 12756 9454
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8673 12940 8978
rect 12898 8664 12954 8673
rect 12898 8599 12954 8608
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12992 7880 13044 7886
rect 12990 7848 12992 7857
rect 13044 7848 13046 7857
rect 12990 7783 13046 7792
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12820 7342 12848 7686
rect 13004 7342 13032 7686
rect 13188 7410 13216 10503
rect 13268 10474 13320 10480
rect 13280 9926 13308 10474
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8498 13308 8910
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13372 7936 13400 11591
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 9110 13492 11494
rect 13648 10062 13676 11698
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 10470 13768 11154
rect 13832 10674 13860 12854
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14002 11928 14058 11937
rect 14002 11863 14058 11872
rect 14016 11694 14044 11863
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13280 7908 13400 7936
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12992 7336 13044 7342
rect 13280 7290 13308 7908
rect 13358 7848 13414 7857
rect 13358 7783 13414 7792
rect 12992 7278 13044 7284
rect 13188 7262 13308 7290
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 6458 12940 6802
rect 13188 6633 13216 7262
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13280 7002 13308 7142
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13372 6798 13400 7783
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13174 6624 13230 6633
rect 13174 6559 13230 6568
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13188 6322 13216 6559
rect 13372 6458 13400 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13188 5642 13216 6054
rect 13372 5778 13400 6394
rect 13464 6322 13492 6802
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 13188 4758 13216 5578
rect 13556 5574 13584 9930
rect 13648 9518 13676 9998
rect 13740 9586 13768 10406
rect 13818 9752 13874 9761
rect 13818 9687 13820 9696
rect 13872 9687 13874 9696
rect 13820 9658 13872 9664
rect 13924 9586 13952 11562
rect 14108 11286 14136 11630
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14108 11150 14136 11222
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10810 14136 11086
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 10266 14044 10542
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9042 13676 9454
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13634 7576 13690 7585
rect 13634 7511 13690 7520
rect 13648 7342 13676 7511
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13832 7274 13860 8230
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 12636 4134 12756 4162
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12636 3602 12664 4134
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12728 3058 12756 3946
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 9496 2440 9548 2446
rect 11336 2440 11388 2446
rect 9496 2382 9548 2388
rect 11256 2400 11336 2428
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10336 480 10364 2314
rect 11256 480 11284 2400
rect 11336 2382 11388 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12176 480 12204 2382
rect 13188 1442 13216 3470
rect 13648 3194 13676 6326
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13740 5370 13768 5782
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13740 4282 13768 4626
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13832 2990 13860 6938
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 14016 6610 14044 9862
rect 14108 7970 14136 10610
rect 14200 10266 14228 12174
rect 14292 11558 14320 14447
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14660 13870 14688 14282
rect 14936 13938 14964 16520
rect 15198 14784 15254 14793
rect 15198 14719 15254 14728
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14660 12646 14688 13466
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14384 10130 14412 11766
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14476 10266 14504 10610
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14476 9518 14504 9998
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14568 9194 14596 9386
rect 14200 9166 14596 9194
rect 14200 8090 14228 9166
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14280 8424 14332 8430
rect 14278 8392 14280 8401
rect 14332 8392 14334 8401
rect 14384 8362 14412 8978
rect 14660 8616 14688 12582
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14752 11014 14780 11562
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10062 14780 10950
rect 14844 10810 14872 11562
rect 15028 11558 15056 12106
rect 15212 12102 15240 14719
rect 15304 12782 15332 16759
rect 15566 16552 15622 16561
rect 18234 16520 18290 17000
rect 15566 16487 15622 16496
rect 15474 13832 15530 13841
rect 15474 13767 15530 13776
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15304 11914 15332 12242
rect 15212 11886 15332 11914
rect 15016 11552 15068 11558
rect 14922 11520 14978 11529
rect 15016 11494 15068 11500
rect 14922 11455 14978 11464
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14830 10704 14886 10713
rect 14830 10639 14886 10648
rect 14844 10130 14872 10639
rect 14936 10606 14964 11455
rect 15028 11218 15056 11494
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15028 10674 15056 11154
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 10600 14976 10606
rect 14922 10568 14924 10577
rect 14976 10568 14978 10577
rect 14922 10503 14978 10512
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14844 9738 14872 10066
rect 15028 9897 15056 10202
rect 15120 10130 15148 11086
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15014 9888 15070 9897
rect 15014 9823 15070 9832
rect 14844 9710 15056 9738
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14476 8588 14688 8616
rect 14278 8327 14334 8336
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14384 8090 14412 8298
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14108 7942 14412 7970
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14108 7449 14136 7822
rect 14094 7440 14150 7449
rect 14094 7375 14150 7384
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14108 7002 14136 7278
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14280 6656 14332 6662
rect 14278 6624 14280 6633
rect 14332 6624 14334 6633
rect 13924 3738 13952 6598
rect 14016 6582 14228 6610
rect 14200 6304 14228 6582
rect 14278 6559 14334 6568
rect 14280 6316 14332 6322
rect 14200 6276 14280 6304
rect 14280 6258 14332 6264
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5778 14044 6054
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14016 4826 14044 5034
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13096 1414 13216 1442
rect 13096 480 13124 1414
rect 13924 480 13952 3062
rect 14108 2922 14136 6190
rect 14292 4690 14320 6258
rect 14384 5114 14412 7942
rect 14476 6118 14504 8588
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14568 6254 14596 8434
rect 14752 8294 14780 9590
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14936 9178 14964 9522
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14844 8498 14872 9046
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14568 5574 14596 6190
rect 14660 5710 14688 6394
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14752 5658 14780 8230
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14844 6934 14872 7278
rect 14832 6928 14884 6934
rect 14832 6870 14884 6876
rect 14844 6458 14872 6870
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 5914 14872 6054
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14936 5710 14964 6258
rect 14924 5704 14976 5710
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14384 5086 14504 5114
rect 14372 5024 14424 5030
rect 14476 5001 14504 5086
rect 14372 4966 14424 4972
rect 14462 4992 14518 5001
rect 14384 4826 14412 4966
rect 14462 4927 14518 4936
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3602 14412 3878
rect 14476 3738 14504 4927
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14568 3534 14596 5510
rect 14660 5370 14688 5646
rect 14752 5630 14872 5658
rect 14924 5646 14976 5652
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14660 4282 14688 5306
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14844 3233 14872 5630
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 5166 14964 5510
rect 15028 5370 15056 9710
rect 15120 9586 15148 10066
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 9110 15148 9522
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15212 8650 15240 11886
rect 15382 11792 15438 11801
rect 15382 11727 15438 11736
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15120 8622 15240 8650
rect 15120 7970 15148 8622
rect 15198 8528 15254 8537
rect 15198 8463 15254 8472
rect 15212 8090 15240 8463
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15120 7942 15240 7970
rect 15212 7886 15240 7942
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15200 7744 15252 7750
rect 15304 7721 15332 10542
rect 15396 9654 15424 11727
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15488 9330 15516 13767
rect 15580 12918 15608 16487
rect 18050 16144 18106 16153
rect 18050 16079 18106 16088
rect 15658 15872 15714 15881
rect 15658 15807 15714 15816
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 10606 15608 12718
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15396 9302 15516 9330
rect 15396 8401 15424 9302
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15382 8392 15438 8401
rect 15382 8327 15438 8336
rect 15382 8120 15438 8129
rect 15488 8090 15516 8774
rect 15382 8055 15438 8064
rect 15476 8084 15528 8090
rect 15200 7686 15252 7692
rect 15290 7712 15346 7721
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14936 4486 14964 5102
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15028 3670 15056 5306
rect 15120 4826 15148 6734
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 14830 3224 14886 3233
rect 14830 3159 14886 3168
rect 15212 2990 15240 7686
rect 15290 7647 15346 7656
rect 15304 6322 15332 7647
rect 15396 7206 15424 8055
rect 15476 8026 15528 8032
rect 15474 7848 15530 7857
rect 15474 7783 15476 7792
rect 15528 7783 15530 7792
rect 15476 7754 15528 7760
rect 15580 7698 15608 10406
rect 15672 9450 15700 15807
rect 17406 15464 17462 15473
rect 17406 15399 17462 15408
rect 16302 15192 16358 15201
rect 16302 15127 16358 15136
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 16210 14104 16266 14113
rect 16210 14039 16212 14048
rect 16264 14039 16266 14048
rect 16212 14010 16264 14016
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16224 13161 16252 13330
rect 16210 13152 16266 13161
rect 15782 13084 16078 13104
rect 16210 13087 16266 13096
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15764 12306 15792 12854
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16132 11665 16160 12378
rect 16118 11656 16174 11665
rect 16118 11591 16174 11600
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16132 10606 16160 11494
rect 16316 10792 16344 15127
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11762 16528 12038
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16394 11112 16450 11121
rect 16394 11047 16450 11056
rect 16224 10764 16344 10792
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 16132 9081 16160 10406
rect 16118 9072 16174 9081
rect 15660 9036 15712 9042
rect 16118 9007 16174 9016
rect 15660 8978 15712 8984
rect 15488 7670 15608 7698
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15382 6896 15438 6905
rect 15382 6831 15438 6840
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15304 4826 15332 5510
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15396 4554 15424 6831
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 3602 15332 4422
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15488 3058 15516 7670
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15580 7449 15608 7482
rect 15566 7440 15622 7449
rect 15566 7375 15622 7384
rect 15672 6458 15700 8978
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16132 8294 16160 8910
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7818 16160 8230
rect 16224 7970 16252 10764
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16316 9926 16344 10610
rect 16408 10470 16436 11047
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9518 16344 9862
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 8634 16344 8978
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16224 7942 16344 7970
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 16132 7274 16160 7754
rect 16224 7546 16252 7822
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16224 6934 16252 7482
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16316 6746 16344 7942
rect 16132 6718 16344 6746
rect 16408 6746 16436 9998
rect 16500 7177 16528 11494
rect 16592 9518 16620 11630
rect 16776 10062 16804 11630
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9874 16804 9998
rect 16684 9846 16804 9874
rect 16684 9722 16712 9846
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16776 9110 16804 9658
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16578 8392 16634 8401
rect 16578 8327 16634 8336
rect 16592 7410 16620 8327
rect 16868 7970 16896 13942
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16946 11792 17002 11801
rect 16946 11727 17002 11736
rect 16960 10010 16988 11727
rect 17052 10674 17080 12038
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17144 11014 17172 11698
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10674 17172 10950
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 10130 17172 10610
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 16960 9982 17080 10010
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16960 8498 16988 9862
rect 17052 8945 17080 9982
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 16776 7942 16896 7970
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16578 7304 16634 7313
rect 16578 7239 16634 7248
rect 16486 7168 16542 7177
rect 16486 7103 16542 7112
rect 16592 7002 16620 7239
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16408 6718 16528 6746
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 16132 6118 16160 6718
rect 16396 6656 16448 6662
rect 16316 6616 16396 6644
rect 16210 6488 16266 6497
rect 16210 6423 16266 6432
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16224 5846 16252 6423
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15580 3942 15608 4490
rect 15672 4282 15700 4558
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 16316 4010 16344 6616
rect 16396 6598 16448 6604
rect 16394 6352 16450 6361
rect 16394 6287 16396 6296
rect 16448 6287 16450 6296
rect 16396 6258 16448 6264
rect 16500 6118 16528 6718
rect 16684 6322 16712 7346
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5030 16436 5646
rect 16486 5128 16542 5137
rect 16486 5063 16542 5072
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4078 16436 4966
rect 16500 4826 16528 5063
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16486 4720 16542 4729
rect 16486 4655 16488 4664
rect 16540 4655 16542 4664
rect 16488 4626 16540 4632
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16776 4010 16804 7942
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16868 7546 16896 7822
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17052 5098 17080 8230
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17144 5778 17172 6598
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5234 17172 5714
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17040 5092 17092 5098
rect 17040 5034 17092 5040
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4146 16988 4966
rect 17052 4593 17080 5034
rect 17038 4584 17094 4593
rect 17038 4519 17094 4528
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17052 4078 17080 4422
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 17236 3738 17264 13806
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10606 17356 10950
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17314 10432 17370 10441
rect 17314 10367 17370 10376
rect 17328 10266 17356 10367
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17420 10169 17448 15399
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 14074 17724 14350
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17590 13560 17646 13569
rect 17590 13495 17646 13504
rect 17604 12646 17632 13495
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12442 17632 12582
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17592 10124 17644 10130
rect 17420 6322 17448 10095
rect 17592 10066 17644 10072
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9722 17540 9998
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17604 9466 17632 10066
rect 17512 9438 17632 9466
rect 17512 8378 17540 9438
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 9217 17632 9318
rect 17590 9208 17646 9217
rect 17590 9143 17646 9152
rect 17696 8838 17724 10542
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17512 8350 17632 8378
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17512 8090 17540 8230
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17604 6118 17632 8350
rect 17696 7342 17724 8774
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17788 7002 17816 11630
rect 17880 9518 17908 12310
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 10130 18000 12242
rect 18064 11286 18092 16079
rect 18248 13870 18276 16520
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18156 11354 18184 12174
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8498 17908 8774
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 8022 17908 8434
rect 18064 8430 18092 10678
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18156 10169 18184 10202
rect 18142 10160 18198 10169
rect 18142 10095 18198 10104
rect 18248 9897 18276 10406
rect 18234 9888 18290 9897
rect 18234 9823 18290 9832
rect 18234 9480 18290 9489
rect 18234 9415 18290 9424
rect 18248 9382 18276 9415
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18340 8809 18368 11494
rect 18326 8800 18382 8809
rect 18326 8735 18382 8744
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7410 17908 7958
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17972 7342 18000 8298
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17696 6254 17724 6802
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17788 6322 17816 6666
rect 17880 6390 17908 6734
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17328 5030 17356 5306
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17316 5024 17368 5030
rect 17408 5024 17460 5030
rect 17316 4966 17368 4972
rect 17406 4992 17408 5001
rect 17460 4992 17462 5001
rect 17406 4927 17462 4936
rect 17420 4672 17448 4927
rect 17500 4684 17552 4690
rect 17420 4644 17500 4672
rect 17500 4626 17552 4632
rect 17604 4622 17632 5170
rect 17696 4826 17724 6190
rect 17788 5574 17816 6258
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5166 17816 5510
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17788 4214 17816 5102
rect 17880 4865 17908 6054
rect 18156 5914 18184 6122
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18248 5545 18276 7142
rect 18340 6225 18368 8502
rect 18326 6216 18382 6225
rect 18326 6151 18382 6160
rect 18418 5808 18474 5817
rect 18418 5743 18474 5752
rect 18234 5536 18290 5545
rect 18234 5471 18290 5480
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 17866 4856 17922 4865
rect 17866 4791 17922 4800
rect 18236 4480 18288 4486
rect 18340 4457 18368 4966
rect 18236 4422 18288 4428
rect 18326 4448 18382 4457
rect 17776 4208 17828 4214
rect 18248 4185 18276 4422
rect 18326 4383 18382 4392
rect 17776 4150 17828 4156
rect 18234 4176 18290 4185
rect 18234 4111 18290 4120
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 17038 3632 17094 3641
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 15660 3528 15712 3534
rect 16316 3505 16344 3538
rect 15660 3470 15712 3476
rect 16118 3496 16174 3505
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14844 480 14872 2858
rect 15672 1442 15700 3470
rect 16118 3431 16174 3440
rect 16302 3496 16358 3505
rect 16302 3431 16358 3440
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16132 2990 16160 3431
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16500 2666 16528 3606
rect 17094 3576 17172 3584
rect 17038 3567 17040 3576
rect 17092 3556 17172 3576
rect 17040 3538 17092 3544
rect 16578 3224 16634 3233
rect 16578 3159 16634 3168
rect 16592 2990 16620 3159
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16670 2952 16726 2961
rect 16670 2887 16726 2896
rect 16764 2916 16816 2922
rect 16500 2638 16620 2666
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16408 2145 16436 2382
rect 16394 2136 16450 2145
rect 16394 2071 16396 2080
rect 16448 2071 16450 2080
rect 16396 2042 16448 2048
rect 16408 2011 16436 2042
rect 16592 1714 16620 2638
rect 16500 1686 16620 1714
rect 15672 1414 15792 1442
rect 15764 480 15792 1414
rect 3422 232 3478 241
rect 3422 167 3478 176
rect 3974 0 4030 480
rect 4894 0 4950 480
rect 5814 0 5870 480
rect 6734 0 6790 480
rect 7562 0 7618 480
rect 8482 0 8538 480
rect 9402 0 9458 480
rect 10322 0 10378 480
rect 11242 0 11298 480
rect 12162 0 12218 480
rect 13082 0 13138 480
rect 13910 0 13966 480
rect 14830 0 14886 480
rect 15750 0 15806 480
rect 16500 241 16528 1686
rect 16684 480 16712 2887
rect 16764 2858 16816 2864
rect 16776 1465 16804 2858
rect 16854 2816 16910 2825
rect 16854 2751 16910 2760
rect 16868 2650 16896 2751
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 16762 1456 16818 1465
rect 16762 1391 16818 1400
rect 17052 1193 17080 2382
rect 17144 1873 17172 3556
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 2990 17356 3334
rect 17420 3058 17448 3674
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17420 2553 17448 2994
rect 17512 2854 17540 4014
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17406 2544 17462 2553
rect 17406 2479 17462 2488
rect 17130 1864 17186 1873
rect 17130 1799 17186 1808
rect 17038 1184 17094 1193
rect 17038 1119 17094 1128
rect 17604 480 17632 3946
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3777 18276 3878
rect 18234 3768 18290 3777
rect 18234 3703 18290 3712
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17788 513 17816 2382
rect 18064 785 18092 3470
rect 18432 3194 18460 5743
rect 18512 3460 18564 3466
rect 18512 3402 18564 3408
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18050 776 18106 785
rect 18050 711 18106 720
rect 17774 504 17830 513
rect 16486 232 16542 241
rect 16486 167 16542 176
rect 16670 0 16726 480
rect 17590 0 17646 480
rect 18524 480 18552 3402
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 17774 439 17830 448
rect 18510 0 18566 480
rect 19430 0 19486 480
<< via2 >>
rect 4066 16768 4122 16824
rect 3422 16496 3478 16552
rect 2962 16088 3018 16144
rect 2870 15136 2926 15192
rect 2778 14728 2834 14784
rect 2778 14456 2834 14512
rect 1766 14048 1822 14104
rect 1858 13812 1860 13832
rect 1860 13812 1912 13832
rect 1912 13812 1914 13832
rect 1858 13776 1914 13812
rect 1306 11464 1362 11520
rect 570 9016 626 9072
rect 570 8472 626 8528
rect 1490 10920 1546 10976
rect 1214 8064 1270 8120
rect 1398 8064 1454 8120
rect 1306 7384 1362 7440
rect 1306 4936 1362 4992
rect 1858 13504 1914 13560
rect 1950 13096 2006 13152
rect 1858 9560 1914 9616
rect 3238 15816 3294 15872
rect 3790 15408 3846 15464
rect 15290 16768 15346 16824
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3054 13812 3056 13832
rect 3056 13812 3108 13832
rect 3108 13812 3110 13832
rect 3054 13776 3110 13812
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3330 12824 3386 12880
rect 2134 9424 2190 9480
rect 1766 5888 1822 5944
rect 1674 5344 1730 5400
rect 1674 3576 1730 3632
rect 1582 2760 1638 2816
rect 2962 12280 3018 12336
rect 2778 11600 2834 11656
rect 2410 7248 2466 7304
rect 2870 10104 2926 10160
rect 2870 6976 2926 7032
rect 2870 6840 2926 6896
rect 3238 12300 3294 12336
rect 3238 12280 3240 12300
rect 3240 12280 3292 12300
rect 3292 12280 3294 12300
rect 4066 12416 4122 12472
rect 3698 12280 3754 12336
rect 3054 10124 3110 10160
rect 3054 10104 3056 10124
rect 3056 10104 3108 10124
rect 3108 10104 3110 10124
rect 3054 9968 3110 10024
rect 3606 12144 3662 12200
rect 2778 5752 2834 5808
rect 2870 5616 2926 5672
rect 2870 2080 2926 2136
rect 3054 4120 3110 4176
rect 2962 1808 3018 1864
rect 3238 5208 3294 5264
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3698 11736 3754 11792
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3790 10376 3846 10432
rect 3698 9832 3754 9888
rect 3974 9968 4030 10024
rect 4342 9968 4398 10024
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4342 9696 4398 9752
rect 3514 8336 3570 8392
rect 3514 4528 3570 4584
rect 3514 3460 3570 3496
rect 3514 3440 3516 3460
rect 3516 3440 3568 3460
rect 3568 3440 3570 3460
rect 3422 3168 3478 3224
rect 3422 3032 3478 3088
rect 3974 8880 4030 8936
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 4066 7792 4122 7848
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3882 6840 3938 6896
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 4066 6196 4068 6216
rect 4068 6196 4120 6216
rect 4120 6196 4122 6216
rect 4066 6160 4122 6196
rect 4158 5788 4160 5808
rect 4160 5788 4212 5808
rect 4212 5788 4214 5808
rect 4158 5752 4214 5788
rect 3698 5480 3754 5536
rect 3698 5208 3754 5264
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 4158 5072 4214 5128
rect 4250 4800 4306 4856
rect 4250 4528 4306 4584
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 4066 4120 4122 4176
rect 3606 1400 3662 1456
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 4710 10376 4766 10432
rect 4710 9152 4766 9208
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 5170 11736 5226 11792
rect 4986 11192 5042 11248
rect 4894 8744 4950 8800
rect 4802 8372 4804 8392
rect 4804 8372 4856 8392
rect 4856 8372 4858 8392
rect 4802 8336 4858 8372
rect 4710 7928 4766 7984
rect 4802 6296 4858 6352
rect 5262 11212 5318 11248
rect 5262 11192 5264 11212
rect 5264 11192 5316 11212
rect 5316 11192 5318 11212
rect 5170 10648 5226 10704
rect 4986 5480 5042 5536
rect 4710 4120 4766 4176
rect 4066 2488 4122 2544
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 3514 1128 3570 1184
rect 3146 448 3202 504
rect 5170 2896 5226 2952
rect 5538 11736 5594 11792
rect 5906 12280 5962 12336
rect 5998 12144 6054 12200
rect 5906 10648 5962 10704
rect 6090 11328 6146 11384
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6734 12280 6790 12336
rect 6458 12144 6514 12200
rect 6458 11328 6514 11384
rect 5538 9016 5594 9072
rect 5722 9988 5778 10024
rect 5722 9968 5724 9988
rect 5724 9968 5776 9988
rect 5776 9968 5778 9988
rect 6090 10376 6146 10432
rect 5998 9016 6054 9072
rect 5538 4664 5594 4720
rect 6274 8472 6330 8528
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 7470 11056 7526 11112
rect 7654 10784 7710 10840
rect 7470 10240 7526 10296
rect 6826 9988 6882 10024
rect 6826 9968 6828 9988
rect 6828 9968 6880 9988
rect 6880 9968 6882 9988
rect 6550 8744 6606 8800
rect 6550 8472 6606 8528
rect 6550 8336 6606 8392
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7378 8880 7434 8936
rect 6826 8356 6882 8392
rect 6826 8336 6828 8356
rect 6828 8336 6880 8356
rect 6880 8336 6882 8356
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6274 6740 6276 6760
rect 6276 6740 6328 6760
rect 6328 6740 6330 6760
rect 6274 6704 6330 6740
rect 5722 4392 5778 4448
rect 6090 5616 6146 5672
rect 5906 4256 5962 4312
rect 5906 3712 5962 3768
rect 5906 3440 5962 3496
rect 6182 3984 6238 4040
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6734 6704 6790 6760
rect 6642 6432 6698 6488
rect 6642 5888 6698 5944
rect 6550 5480 6606 5536
rect 6458 4972 6460 4992
rect 6460 4972 6512 4992
rect 6512 4972 6514 4992
rect 6458 4936 6514 4972
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6550 4120 6606 4176
rect 6366 3032 6422 3088
rect 7010 4120 7066 4176
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 14278 14456 14334 14512
rect 7838 11736 7894 11792
rect 7562 7248 7618 7304
rect 7470 4256 7526 4312
rect 8298 10512 8354 10568
rect 8206 9016 8262 9072
rect 8298 8880 8354 8936
rect 8206 8336 8262 8392
rect 8574 11600 8630 11656
rect 8482 11056 8538 11112
rect 8482 10240 8538 10296
rect 8942 12316 8944 12336
rect 8944 12316 8996 12336
rect 8996 12316 8998 12336
rect 8942 12280 8998 12316
rect 10966 13268 10968 13288
rect 10968 13268 11020 13288
rect 11020 13268 11022 13288
rect 10966 13232 11022 13268
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9034 12144 9090 12200
rect 9494 9560 9550 9616
rect 8850 8880 8906 8936
rect 10138 12280 10194 12336
rect 9954 12144 10010 12200
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10138 11636 10140 11656
rect 10140 11636 10192 11656
rect 10192 11636 10194 11656
rect 10138 11600 10194 11636
rect 9862 11228 9864 11248
rect 9864 11228 9916 11248
rect 9916 11228 9918 11248
rect 9862 11192 9918 11228
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10046 10648 10102 10704
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10322 9968 10378 10024
rect 10046 9152 10102 9208
rect 10598 11600 10654 11656
rect 10506 11056 10562 11112
rect 10782 11892 10838 11928
rect 10782 11872 10784 11892
rect 10784 11872 10836 11892
rect 10836 11872 10838 11892
rect 10506 9832 10562 9888
rect 10598 9696 10654 9752
rect 10598 9424 10654 9480
rect 10506 9152 10562 9208
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 7746 7112 7802 7168
rect 7746 4664 7802 4720
rect 7654 3984 7710 4040
rect 7562 2760 7618 2816
rect 7930 4392 7986 4448
rect 8574 6296 8630 6352
rect 8390 5752 8446 5808
rect 8482 5480 8538 5536
rect 9586 6840 9642 6896
rect 10138 8200 10194 8256
rect 9954 8064 10010 8120
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10414 8880 10470 8936
rect 10506 8608 10562 8664
rect 8298 4120 8354 4176
rect 8114 720 8170 776
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9586 4548 9642 4584
rect 9586 4528 9588 4548
rect 9588 4528 9640 4548
rect 9640 4528 9642 4548
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10046 4664 10102 4720
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 11150 12824 11206 12880
rect 11426 12280 11482 12336
rect 11242 12144 11298 12200
rect 11242 11736 11298 11792
rect 11242 9560 11298 9616
rect 11150 9016 11206 9072
rect 10874 7928 10930 7984
rect 10598 3440 10654 3496
rect 10598 3168 10654 3224
rect 10506 2760 10562 2816
rect 11150 8200 11206 8256
rect 10966 6452 11022 6488
rect 11426 8200 11482 8256
rect 10966 6432 10968 6452
rect 10968 6432 11020 6452
rect 11020 6432 11022 6452
rect 11702 11600 11758 11656
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 11978 10104 12034 10160
rect 11702 8236 11704 8256
rect 11704 8236 11756 8256
rect 11756 8236 11758 8256
rect 11702 8200 11758 8236
rect 11886 7520 11942 7576
rect 11794 7404 11850 7440
rect 11794 7384 11796 7404
rect 11796 7384 11848 7404
rect 11848 7384 11850 7404
rect 11794 7248 11850 7304
rect 12254 11212 12310 11248
rect 12254 11192 12256 11212
rect 12256 11192 12308 11212
rect 12308 11192 12310 11212
rect 12254 10512 12310 10568
rect 12254 9560 12310 9616
rect 12070 8064 12126 8120
rect 12346 7928 12402 7984
rect 12254 7692 12256 7712
rect 12256 7692 12308 7712
rect 12308 7692 12310 7712
rect 12254 7656 12310 7692
rect 12162 7248 12218 7304
rect 12162 7148 12164 7168
rect 12164 7148 12216 7168
rect 12216 7148 12218 7168
rect 12162 7112 12218 7148
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12714 11600 12770 11656
rect 13358 11600 13414 11656
rect 12530 11092 12532 11112
rect 12532 11092 12584 11112
rect 12584 11092 12586 11112
rect 12530 11056 12586 11092
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12530 9716 12586 9752
rect 12530 9696 12532 9716
rect 12532 9696 12584 9716
rect 12584 9696 12586 9716
rect 13266 10648 13322 10704
rect 13174 10512 13230 10568
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12806 9968 12862 10024
rect 12530 8200 12586 8256
rect 10874 3052 10930 3088
rect 10874 3032 10876 3052
rect 10876 3032 10928 3052
rect 10928 3032 10930 3052
rect 11334 4528 11390 4584
rect 12162 3984 12218 4040
rect 12622 6432 12678 6488
rect 12438 3848 12494 3904
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12898 8608 12954 8664
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12990 7828 12992 7848
rect 12992 7828 13044 7848
rect 13044 7828 13046 7848
rect 12990 7792 13046 7828
rect 14002 11872 14058 11928
rect 13358 7792 13414 7848
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 13174 6568 13230 6624
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13818 9716 13874 9752
rect 13818 9696 13820 9716
rect 13820 9696 13872 9716
rect 13872 9696 13874 9716
rect 13634 7520 13690 7576
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 15198 14728 15254 14784
rect 14278 8372 14280 8392
rect 14280 8372 14332 8392
rect 14332 8372 14334 8392
rect 14278 8336 14334 8372
rect 15566 16496 15622 16552
rect 15474 13776 15530 13832
rect 14922 11464 14978 11520
rect 14830 10648 14886 10704
rect 14922 10548 14924 10568
rect 14924 10548 14976 10568
rect 14976 10548 14978 10568
rect 14922 10512 14978 10548
rect 15014 9832 15070 9888
rect 14094 7384 14150 7440
rect 14278 6604 14280 6624
rect 14280 6604 14332 6624
rect 14332 6604 14334 6624
rect 14278 6568 14334 6604
rect 14462 4936 14518 4992
rect 15382 11736 15438 11792
rect 15198 8472 15254 8528
rect 18050 16088 18106 16144
rect 15658 15816 15714 15872
rect 15382 8336 15438 8392
rect 15382 8064 15438 8120
rect 14830 3168 14886 3224
rect 15290 7656 15346 7712
rect 15474 7812 15530 7848
rect 15474 7792 15476 7812
rect 15476 7792 15528 7812
rect 15528 7792 15530 7812
rect 17406 15408 17462 15464
rect 16302 15136 16358 15192
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 16210 14068 16266 14104
rect 16210 14048 16212 14068
rect 16212 14048 16264 14068
rect 16264 14048 16266 14068
rect 16210 13096 16266 13152
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16118 11600 16174 11656
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 16394 11056 16450 11112
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 16118 9016 16174 9072
rect 15382 6840 15438 6896
rect 15566 7384 15622 7440
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 16578 8336 16634 8392
rect 16946 11736 17002 11792
rect 17038 8880 17094 8936
rect 16578 7248 16634 7304
rect 16486 7112 16542 7168
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 16210 6432 16266 6488
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 16394 6316 16450 6352
rect 16394 6296 16396 6316
rect 16396 6296 16448 6316
rect 16448 6296 16450 6316
rect 16486 5072 16542 5128
rect 16486 4684 16542 4720
rect 16486 4664 16488 4684
rect 16488 4664 16540 4684
rect 16540 4664 16542 4684
rect 17038 4528 17094 4584
rect 17314 10376 17370 10432
rect 17590 13504 17646 13560
rect 17406 10104 17462 10160
rect 17590 9152 17646 9208
rect 18142 10104 18198 10160
rect 18234 9832 18290 9888
rect 18234 9424 18290 9480
rect 18326 8744 18382 8800
rect 17406 4972 17408 4992
rect 17408 4972 17460 4992
rect 17460 4972 17462 4992
rect 17406 4936 17462 4972
rect 18326 6160 18382 6216
rect 18418 5752 18474 5808
rect 18234 5480 18290 5536
rect 17866 4800 17922 4856
rect 18326 4392 18382 4448
rect 18234 4120 18290 4176
rect 16118 3440 16174 3496
rect 16302 3440 16358 3496
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 17038 3596 17094 3632
rect 17038 3576 17040 3596
rect 17040 3576 17092 3596
rect 17092 3576 17094 3596
rect 16578 3168 16634 3224
rect 16670 2896 16726 2952
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16394 2100 16450 2136
rect 16394 2080 16396 2100
rect 16396 2080 16448 2100
rect 16448 2080 16450 2100
rect 3422 176 3478 232
rect 16854 2760 16910 2816
rect 16762 1400 16818 1456
rect 17406 2488 17462 2544
rect 17130 1808 17186 1864
rect 17038 1128 17094 1184
rect 18234 3712 18290 3768
rect 18050 720 18106 776
rect 16486 176 16542 232
rect 17774 448 17830 504
<< metal3 >>
rect 0 16826 480 16856
rect 4061 16826 4127 16829
rect 0 16824 4127 16826
rect 0 16768 4066 16824
rect 4122 16768 4127 16824
rect 0 16766 4127 16768
rect 0 16736 480 16766
rect 4061 16763 4127 16766
rect 15285 16826 15351 16829
rect 19520 16826 20000 16856
rect 15285 16824 20000 16826
rect 15285 16768 15290 16824
rect 15346 16768 20000 16824
rect 15285 16766 20000 16768
rect 15285 16763 15351 16766
rect 19520 16736 20000 16766
rect 0 16554 480 16584
rect 3417 16554 3483 16557
rect 0 16552 3483 16554
rect 0 16496 3422 16552
rect 3478 16496 3483 16552
rect 0 16494 3483 16496
rect 0 16464 480 16494
rect 3417 16491 3483 16494
rect 15561 16554 15627 16557
rect 19520 16554 20000 16584
rect 15561 16552 20000 16554
rect 15561 16496 15566 16552
rect 15622 16496 20000 16552
rect 15561 16494 20000 16496
rect 15561 16491 15627 16494
rect 19520 16464 20000 16494
rect 0 16146 480 16176
rect 2957 16146 3023 16149
rect 0 16144 3023 16146
rect 0 16088 2962 16144
rect 3018 16088 3023 16144
rect 0 16086 3023 16088
rect 0 16056 480 16086
rect 2957 16083 3023 16086
rect 18045 16146 18111 16149
rect 19520 16146 20000 16176
rect 18045 16144 20000 16146
rect 18045 16088 18050 16144
rect 18106 16088 20000 16144
rect 18045 16086 20000 16088
rect 18045 16083 18111 16086
rect 19520 16056 20000 16086
rect 0 15874 480 15904
rect 3233 15874 3299 15877
rect 0 15872 3299 15874
rect 0 15816 3238 15872
rect 3294 15816 3299 15872
rect 0 15814 3299 15816
rect 0 15784 480 15814
rect 3233 15811 3299 15814
rect 15653 15874 15719 15877
rect 19520 15874 20000 15904
rect 15653 15872 20000 15874
rect 15653 15816 15658 15872
rect 15714 15816 20000 15872
rect 15653 15814 20000 15816
rect 15653 15811 15719 15814
rect 19520 15784 20000 15814
rect 0 15466 480 15496
rect 3785 15466 3851 15469
rect 0 15464 3851 15466
rect 0 15408 3790 15464
rect 3846 15408 3851 15464
rect 0 15406 3851 15408
rect 0 15376 480 15406
rect 3785 15403 3851 15406
rect 17401 15466 17467 15469
rect 19520 15466 20000 15496
rect 17401 15464 20000 15466
rect 17401 15408 17406 15464
rect 17462 15408 20000 15464
rect 17401 15406 20000 15408
rect 17401 15403 17467 15406
rect 19520 15376 20000 15406
rect 0 15194 480 15224
rect 2865 15194 2931 15197
rect 0 15192 2931 15194
rect 0 15136 2870 15192
rect 2926 15136 2931 15192
rect 0 15134 2931 15136
rect 0 15104 480 15134
rect 2865 15131 2931 15134
rect 16297 15194 16363 15197
rect 19520 15194 20000 15224
rect 16297 15192 20000 15194
rect 16297 15136 16302 15192
rect 16358 15136 20000 15192
rect 16297 15134 20000 15136
rect 16297 15131 16363 15134
rect 19520 15104 20000 15134
rect 0 14786 480 14816
rect 2773 14786 2839 14789
rect 0 14784 2839 14786
rect 0 14728 2778 14784
rect 2834 14728 2839 14784
rect 0 14726 2839 14728
rect 0 14696 480 14726
rect 2773 14723 2839 14726
rect 15193 14786 15259 14789
rect 19520 14786 20000 14816
rect 15193 14784 20000 14786
rect 15193 14728 15198 14784
rect 15254 14728 20000 14784
rect 15193 14726 20000 14728
rect 15193 14723 15259 14726
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 19520 14696 20000 14726
rect 12805 14655 13125 14656
rect 0 14514 480 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 480 14454
rect 2773 14451 2839 14454
rect 14273 14514 14339 14517
rect 19520 14514 20000 14544
rect 14273 14512 20000 14514
rect 14273 14456 14278 14512
rect 14334 14456 20000 14512
rect 14273 14454 20000 14456
rect 14273 14451 14339 14454
rect 19520 14424 20000 14454
rect 3909 14176 4229 14177
rect 0 14106 480 14136
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 14111 16090 14112
rect 1761 14106 1827 14109
rect 0 14104 1827 14106
rect 0 14048 1766 14104
rect 1822 14048 1827 14104
rect 0 14046 1827 14048
rect 0 14016 480 14046
rect 1761 14043 1827 14046
rect 16205 14106 16271 14109
rect 19520 14106 20000 14136
rect 16205 14104 20000 14106
rect 16205 14048 16210 14104
rect 16266 14048 20000 14104
rect 16205 14046 20000 14048
rect 16205 14043 16271 14046
rect 19520 14016 20000 14046
rect 0 13834 480 13864
rect 1853 13834 1919 13837
rect 0 13832 1919 13834
rect 0 13776 1858 13832
rect 1914 13776 1919 13832
rect 0 13774 1919 13776
rect 0 13744 480 13774
rect 1853 13771 1919 13774
rect 3049 13834 3115 13837
rect 3366 13834 3372 13836
rect 3049 13832 3372 13834
rect 3049 13776 3054 13832
rect 3110 13776 3372 13832
rect 3049 13774 3372 13776
rect 3049 13771 3115 13774
rect 3366 13772 3372 13774
rect 3436 13772 3442 13836
rect 15469 13834 15535 13837
rect 19520 13834 20000 13864
rect 15469 13832 20000 13834
rect 15469 13776 15474 13832
rect 15530 13776 20000 13832
rect 15469 13774 20000 13776
rect 15469 13771 15535 13774
rect 19520 13744 20000 13774
rect 6874 13632 7194 13633
rect 0 13562 480 13592
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 1853 13562 1919 13565
rect 0 13560 1919 13562
rect 0 13504 1858 13560
rect 1914 13504 1919 13560
rect 0 13502 1919 13504
rect 0 13472 480 13502
rect 1853 13499 1919 13502
rect 17585 13562 17651 13565
rect 19520 13562 20000 13592
rect 17585 13560 20000 13562
rect 17585 13504 17590 13560
rect 17646 13504 20000 13560
rect 17585 13502 20000 13504
rect 17585 13499 17651 13502
rect 19520 13472 20000 13502
rect 10542 13228 10548 13292
rect 10612 13290 10618 13292
rect 10961 13290 11027 13293
rect 10612 13288 11027 13290
rect 10612 13232 10966 13288
rect 11022 13232 11027 13288
rect 10612 13230 11027 13232
rect 10612 13228 10618 13230
rect 10961 13227 11027 13230
rect 0 13154 480 13184
rect 1945 13154 2011 13157
rect 0 13152 2011 13154
rect 0 13096 1950 13152
rect 2006 13096 2011 13152
rect 0 13094 2011 13096
rect 0 13064 480 13094
rect 1945 13091 2011 13094
rect 16205 13154 16271 13157
rect 19520 13154 20000 13184
rect 16205 13152 20000 13154
rect 16205 13096 16210 13152
rect 16266 13096 20000 13152
rect 16205 13094 20000 13096
rect 16205 13091 16271 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 19520 13064 20000 13094
rect 15770 13023 16090 13024
rect 0 12882 480 12912
rect 3325 12882 3391 12885
rect 0 12880 3391 12882
rect 0 12824 3330 12880
rect 3386 12824 3391 12880
rect 0 12822 3391 12824
rect 0 12792 480 12822
rect 3325 12819 3391 12822
rect 11145 12882 11211 12885
rect 19520 12882 20000 12912
rect 11145 12880 20000 12882
rect 11145 12824 11150 12880
rect 11206 12824 20000 12880
rect 11145 12822 20000 12824
rect 11145 12819 11211 12822
rect 19520 12792 20000 12822
rect 6874 12544 7194 12545
rect 0 12474 480 12504
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 4061 12474 4127 12477
rect 19520 12474 20000 12504
rect 0 12472 4127 12474
rect 0 12416 4066 12472
rect 4122 12416 4127 12472
rect 0 12414 4127 12416
rect 0 12384 480 12414
rect 4061 12411 4127 12414
rect 13310 12414 20000 12474
rect 2957 12338 3023 12341
rect 3233 12338 3299 12341
rect 2957 12336 3299 12338
rect 2957 12280 2962 12336
rect 3018 12280 3238 12336
rect 3294 12280 3299 12336
rect 2957 12278 3299 12280
rect 2957 12275 3023 12278
rect 3233 12275 3299 12278
rect 3693 12338 3759 12341
rect 4838 12338 4844 12340
rect 3693 12336 4844 12338
rect 3693 12280 3698 12336
rect 3754 12280 4844 12336
rect 3693 12278 4844 12280
rect 3693 12275 3759 12278
rect 4838 12276 4844 12278
rect 4908 12276 4914 12340
rect 5901 12338 5967 12341
rect 6729 12338 6795 12341
rect 8937 12338 9003 12341
rect 5901 12336 9003 12338
rect 5901 12280 5906 12336
rect 5962 12280 6734 12336
rect 6790 12280 8942 12336
rect 8998 12280 9003 12336
rect 5901 12278 9003 12280
rect 5901 12275 5967 12278
rect 6729 12275 6795 12278
rect 8937 12275 9003 12278
rect 10133 12338 10199 12341
rect 10358 12338 10364 12340
rect 10133 12336 10364 12338
rect 10133 12280 10138 12336
rect 10194 12280 10364 12336
rect 10133 12278 10364 12280
rect 10133 12275 10199 12278
rect 10358 12276 10364 12278
rect 10428 12276 10434 12340
rect 11421 12338 11487 12341
rect 13310 12338 13370 12414
rect 19520 12384 20000 12414
rect 11421 12336 13370 12338
rect 11421 12280 11426 12336
rect 11482 12280 13370 12336
rect 11421 12278 13370 12280
rect 11421 12275 11487 12278
rect 0 12202 480 12232
rect 3601 12202 3667 12205
rect 0 12200 3667 12202
rect 0 12144 3606 12200
rect 3662 12144 3667 12200
rect 0 12142 3667 12144
rect 0 12112 480 12142
rect 3601 12139 3667 12142
rect 5993 12202 6059 12205
rect 6453 12202 6519 12205
rect 9029 12202 9095 12205
rect 5993 12200 9095 12202
rect 5993 12144 5998 12200
rect 6054 12144 6458 12200
rect 6514 12144 9034 12200
rect 9090 12144 9095 12200
rect 5993 12142 9095 12144
rect 5993 12139 6059 12142
rect 6453 12139 6519 12142
rect 9029 12139 9095 12142
rect 9949 12202 10015 12205
rect 11237 12202 11303 12205
rect 19520 12202 20000 12232
rect 9949 12200 11303 12202
rect 9949 12144 9954 12200
rect 10010 12144 11242 12200
rect 11298 12144 11303 12200
rect 9949 12142 11303 12144
rect 9949 12139 10015 12142
rect 11237 12139 11303 12142
rect 15518 12142 20000 12202
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 10777 11930 10843 11933
rect 13997 11930 14063 11933
rect 10777 11928 14063 11930
rect 10777 11872 10782 11928
rect 10838 11872 14002 11928
rect 14058 11872 14063 11928
rect 10777 11870 14063 11872
rect 10777 11867 10843 11870
rect 13997 11867 14063 11870
rect 0 11794 480 11824
rect 3693 11794 3759 11797
rect 0 11792 3759 11794
rect 0 11736 3698 11792
rect 3754 11736 3759 11792
rect 0 11734 3759 11736
rect 0 11704 480 11734
rect 3693 11731 3759 11734
rect 5165 11794 5231 11797
rect 5533 11794 5599 11797
rect 5165 11792 5599 11794
rect 5165 11736 5170 11792
rect 5226 11736 5538 11792
rect 5594 11736 5599 11792
rect 5165 11734 5599 11736
rect 5165 11731 5231 11734
rect 5533 11731 5599 11734
rect 7833 11794 7899 11797
rect 11237 11794 11303 11797
rect 7833 11792 11303 11794
rect 7833 11736 7838 11792
rect 7894 11736 11242 11792
rect 11298 11736 11303 11792
rect 7833 11734 11303 11736
rect 7833 11731 7899 11734
rect 11237 11731 11303 11734
rect 15377 11794 15443 11797
rect 15518 11794 15578 12142
rect 19520 12112 20000 12142
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 15377 11792 15578 11794
rect 15377 11736 15382 11792
rect 15438 11736 15578 11792
rect 15377 11734 15578 11736
rect 16941 11794 17007 11797
rect 19520 11794 20000 11824
rect 16941 11792 20000 11794
rect 16941 11736 16946 11792
rect 17002 11736 20000 11792
rect 16941 11734 20000 11736
rect 15377 11731 15443 11734
rect 16941 11731 17007 11734
rect 19520 11704 20000 11734
rect 2773 11658 2839 11661
rect 8569 11658 8635 11661
rect 2773 11656 8635 11658
rect 2773 11600 2778 11656
rect 2834 11600 8574 11656
rect 8630 11600 8635 11656
rect 2773 11598 8635 11600
rect 2773 11595 2839 11598
rect 8569 11595 8635 11598
rect 10133 11658 10199 11661
rect 10593 11658 10659 11661
rect 10133 11656 10659 11658
rect 10133 11600 10138 11656
rect 10194 11600 10598 11656
rect 10654 11600 10659 11656
rect 10133 11598 10659 11600
rect 10133 11595 10199 11598
rect 10593 11595 10659 11598
rect 11697 11658 11763 11661
rect 12709 11658 12775 11661
rect 13353 11658 13419 11661
rect 16113 11658 16179 11661
rect 11697 11656 16179 11658
rect 11697 11600 11702 11656
rect 11758 11600 12714 11656
rect 12770 11600 13358 11656
rect 13414 11600 16118 11656
rect 16174 11600 16179 11656
rect 11697 11598 16179 11600
rect 11697 11595 11763 11598
rect 12709 11595 12775 11598
rect 13353 11595 13419 11598
rect 16113 11595 16179 11598
rect 0 11522 480 11552
rect 1301 11522 1367 11525
rect 0 11520 1367 11522
rect 0 11464 1306 11520
rect 1362 11464 1367 11520
rect 0 11462 1367 11464
rect 0 11432 480 11462
rect 1301 11459 1367 11462
rect 14917 11522 14983 11525
rect 19520 11522 20000 11552
rect 14917 11520 20000 11522
rect 14917 11464 14922 11520
rect 14978 11464 20000 11520
rect 14917 11462 20000 11464
rect 14917 11459 14983 11462
rect 6874 11456 7194 11457
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 19520 11432 20000 11462
rect 12805 11391 13125 11392
rect 6085 11386 6151 11389
rect 6453 11386 6519 11389
rect 6085 11384 6519 11386
rect 6085 11328 6090 11384
rect 6146 11328 6458 11384
rect 6514 11328 6519 11384
rect 6085 11326 6519 11328
rect 6085 11323 6151 11326
rect 6453 11323 6519 11326
rect 4981 11250 5047 11253
rect 5257 11250 5323 11253
rect 4981 11248 5323 11250
rect 4981 11192 4986 11248
rect 5042 11192 5262 11248
rect 5318 11192 5323 11248
rect 4981 11190 5323 11192
rect 4981 11187 5047 11190
rect 5257 11187 5323 11190
rect 9857 11250 9923 11253
rect 12249 11250 12315 11253
rect 9857 11248 12315 11250
rect 9857 11192 9862 11248
rect 9918 11192 12254 11248
rect 12310 11192 12315 11248
rect 9857 11190 12315 11192
rect 9857 11187 9923 11190
rect 12249 11187 12315 11190
rect 0 11114 480 11144
rect 2998 11114 3004 11116
rect 0 11054 3004 11114
rect 0 11024 480 11054
rect 2998 11052 3004 11054
rect 3068 11052 3074 11116
rect 7465 11114 7531 11117
rect 8477 11114 8543 11117
rect 3788 11112 8543 11114
rect 3788 11056 7470 11112
rect 7526 11056 8482 11112
rect 8538 11056 8543 11112
rect 3788 11054 8543 11056
rect 1485 10978 1551 10981
rect 3788 10978 3848 11054
rect 7465 11051 7531 11054
rect 8477 11051 8543 11054
rect 10501 11114 10567 11117
rect 12525 11114 12591 11117
rect 10501 11112 12591 11114
rect 10501 11056 10506 11112
rect 10562 11056 12530 11112
rect 12586 11056 12591 11112
rect 10501 11054 12591 11056
rect 10501 11051 10567 11054
rect 12525 11051 12591 11054
rect 16389 11114 16455 11117
rect 19520 11114 20000 11144
rect 16389 11112 20000 11114
rect 16389 11056 16394 11112
rect 16450 11056 20000 11112
rect 16389 11054 20000 11056
rect 16389 11051 16455 11054
rect 19520 11024 20000 11054
rect 1485 10976 3848 10978
rect 1485 10920 1490 10976
rect 1546 10920 3848 10976
rect 1485 10918 3848 10920
rect 1485 10915 1551 10918
rect 3909 10912 4229 10913
rect 0 10842 480 10872
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 7649 10842 7715 10845
rect 19520 10842 20000 10872
rect 0 10782 3848 10842
rect 0 10752 480 10782
rect 3788 10706 3848 10782
rect 5030 10840 7715 10842
rect 5030 10784 7654 10840
rect 7710 10784 7715 10840
rect 5030 10782 7715 10784
rect 5030 10706 5090 10782
rect 7649 10779 7715 10782
rect 16254 10782 20000 10842
rect 3788 10646 5090 10706
rect 5165 10706 5231 10709
rect 5901 10706 5967 10709
rect 5165 10704 5967 10706
rect 5165 10648 5170 10704
rect 5226 10648 5906 10704
rect 5962 10648 5967 10704
rect 5165 10646 5967 10648
rect 5165 10643 5231 10646
rect 5901 10643 5967 10646
rect 10041 10706 10107 10709
rect 13261 10706 13327 10709
rect 10041 10704 13327 10706
rect 10041 10648 10046 10704
rect 10102 10648 13266 10704
rect 13322 10648 13327 10704
rect 10041 10646 13327 10648
rect 10041 10643 10107 10646
rect 13261 10643 13327 10646
rect 14825 10706 14891 10709
rect 16254 10706 16314 10782
rect 19520 10752 20000 10782
rect 14825 10704 16314 10706
rect 14825 10648 14830 10704
rect 14886 10648 16314 10704
rect 14825 10646 16314 10648
rect 14825 10643 14891 10646
rect 8293 10570 8359 10573
rect 4064 10568 8359 10570
rect 4064 10512 8298 10568
rect 8354 10512 8359 10568
rect 4064 10510 8359 10512
rect 0 10434 480 10464
rect 3785 10434 3851 10437
rect 0 10432 3851 10434
rect 0 10376 3790 10432
rect 3846 10376 3851 10432
rect 0 10374 3851 10376
rect 0 10344 480 10374
rect 3785 10371 3851 10374
rect 4064 10298 4124 10510
rect 8293 10507 8359 10510
rect 12249 10570 12315 10573
rect 13169 10570 13235 10573
rect 14917 10570 14983 10573
rect 12249 10568 14983 10570
rect 12249 10512 12254 10568
rect 12310 10512 13174 10568
rect 13230 10512 14922 10568
rect 14978 10512 14983 10568
rect 12249 10510 14983 10512
rect 12249 10507 12315 10510
rect 13169 10507 13235 10510
rect 14917 10507 14983 10510
rect 4705 10434 4771 10437
rect 6085 10434 6151 10437
rect 4705 10432 6151 10434
rect 4705 10376 4710 10432
rect 4766 10376 6090 10432
rect 6146 10376 6151 10432
rect 4705 10374 6151 10376
rect 4705 10371 4771 10374
rect 6085 10371 6151 10374
rect 17309 10434 17375 10437
rect 19520 10434 20000 10464
rect 17309 10432 20000 10434
rect 17309 10376 17314 10432
rect 17370 10376 20000 10432
rect 17309 10374 20000 10376
rect 17309 10371 17375 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19520 10344 20000 10374
rect 12805 10303 13125 10304
rect 2822 10238 4124 10298
rect 7465 10298 7531 10301
rect 8477 10298 8543 10301
rect 7465 10296 8543 10298
rect 7465 10240 7470 10296
rect 7526 10240 8482 10296
rect 8538 10240 8543 10296
rect 7465 10238 8543 10240
rect 0 10162 480 10192
rect 2822 10165 2882 10238
rect 7465 10235 7531 10238
rect 8477 10235 8543 10238
rect 2822 10162 2931 10165
rect 0 10160 2931 10162
rect 0 10104 2870 10160
rect 2926 10104 2931 10160
rect 0 10102 2931 10104
rect 0 10072 480 10102
rect 2865 10099 2931 10102
rect 3049 10162 3115 10165
rect 11973 10162 12039 10165
rect 17401 10162 17467 10165
rect 3049 10160 17467 10162
rect 3049 10104 3054 10160
rect 3110 10104 11978 10160
rect 12034 10104 17406 10160
rect 17462 10104 17467 10160
rect 3049 10102 17467 10104
rect 3049 10099 3115 10102
rect 11973 10099 12039 10102
rect 17401 10099 17467 10102
rect 18137 10162 18203 10165
rect 19520 10162 20000 10192
rect 18137 10160 20000 10162
rect 18137 10104 18142 10160
rect 18198 10104 20000 10160
rect 18137 10102 20000 10104
rect 18137 10099 18203 10102
rect 19520 10072 20000 10102
rect 3049 10028 3115 10029
rect 2998 9964 3004 10028
rect 3068 10026 3115 10028
rect 3068 10024 3160 10026
rect 3110 9968 3160 10024
rect 3068 9966 3160 9968
rect 3068 9964 3115 9966
rect 3734 9964 3740 10028
rect 3804 10026 3810 10028
rect 3969 10026 4035 10029
rect 3804 10024 4035 10026
rect 3804 9968 3974 10024
rect 4030 9968 4035 10024
rect 3804 9966 4035 9968
rect 3804 9964 3810 9966
rect 3049 9963 3115 9964
rect 3969 9963 4035 9966
rect 4337 10026 4403 10029
rect 5717 10026 5783 10029
rect 6821 10026 6887 10029
rect 4337 10024 4538 10026
rect 4337 9968 4342 10024
rect 4398 9968 4538 10024
rect 4337 9966 4538 9968
rect 4337 9963 4403 9966
rect 0 9890 480 9920
rect 3693 9890 3759 9893
rect 0 9888 3759 9890
rect 0 9832 3698 9888
rect 3754 9832 3759 9888
rect 0 9830 3759 9832
rect 0 9800 480 9830
rect 3693 9827 3759 9830
rect 3909 9824 4229 9825
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 4337 9754 4403 9757
rect 4478 9754 4538 9966
rect 5717 10024 6887 10026
rect 5717 9968 5722 10024
rect 5778 9968 6826 10024
rect 6882 9968 6887 10024
rect 5717 9966 6887 9968
rect 5717 9963 5783 9966
rect 6821 9963 6887 9966
rect 10317 10026 10383 10029
rect 12801 10026 12867 10029
rect 10317 10024 12867 10026
rect 10317 9968 10322 10024
rect 10378 9968 12806 10024
rect 12862 9968 12867 10024
rect 10317 9966 12867 9968
rect 10317 9963 10383 9966
rect 12801 9963 12867 9966
rect 10358 9828 10364 9892
rect 10428 9890 10434 9892
rect 10501 9890 10567 9893
rect 15009 9890 15075 9893
rect 10428 9888 15075 9890
rect 10428 9832 10506 9888
rect 10562 9832 15014 9888
rect 15070 9832 15075 9888
rect 10428 9830 15075 9832
rect 10428 9828 10434 9830
rect 10501 9827 10567 9830
rect 15009 9827 15075 9830
rect 18229 9890 18295 9893
rect 19520 9890 20000 9920
rect 18229 9888 20000 9890
rect 18229 9832 18234 9888
rect 18290 9832 20000 9888
rect 18229 9830 20000 9832
rect 18229 9827 18295 9830
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19520 9800 20000 9830
rect 15770 9759 16090 9760
rect 10593 9756 10659 9757
rect 4337 9752 4538 9754
rect 4337 9696 4342 9752
rect 4398 9696 4538 9752
rect 4337 9694 4538 9696
rect 4337 9691 4403 9694
rect 10542 9692 10548 9756
rect 10612 9754 10659 9756
rect 12525 9754 12591 9757
rect 13813 9754 13879 9757
rect 10612 9752 10704 9754
rect 10654 9696 10704 9752
rect 10612 9694 10704 9696
rect 12525 9752 13879 9754
rect 12525 9696 12530 9752
rect 12586 9696 13818 9752
rect 13874 9696 13879 9752
rect 12525 9694 13879 9696
rect 10612 9692 10659 9694
rect 10593 9691 10659 9692
rect 12525 9691 12591 9694
rect 13813 9691 13879 9694
rect 1853 9618 1919 9621
rect 9489 9618 9555 9621
rect 1853 9616 9555 9618
rect 1853 9560 1858 9616
rect 1914 9560 9494 9616
rect 9550 9560 9555 9616
rect 1853 9558 9555 9560
rect 1853 9555 1919 9558
rect 9489 9555 9555 9558
rect 11237 9618 11303 9621
rect 12249 9618 12315 9621
rect 11237 9616 12315 9618
rect 11237 9560 11242 9616
rect 11298 9560 12254 9616
rect 12310 9560 12315 9616
rect 11237 9558 12315 9560
rect 11237 9555 11303 9558
rect 12249 9555 12315 9558
rect 0 9482 480 9512
rect 2129 9482 2195 9485
rect 10593 9482 10659 9485
rect 0 9480 10659 9482
rect 0 9424 2134 9480
rect 2190 9424 10598 9480
rect 10654 9424 10659 9480
rect 0 9422 10659 9424
rect 0 9392 480 9422
rect 2129 9419 2195 9422
rect 10593 9419 10659 9422
rect 18229 9482 18295 9485
rect 19520 9482 20000 9512
rect 18229 9480 20000 9482
rect 18229 9424 18234 9480
rect 18290 9424 20000 9480
rect 18229 9422 20000 9424
rect 18229 9419 18295 9422
rect 19520 9392 20000 9422
rect 6874 9280 7194 9281
rect 0 9210 480 9240
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 4705 9210 4771 9213
rect 6494 9210 6500 9212
rect 0 9208 4771 9210
rect 0 9152 4710 9208
rect 4766 9152 4771 9208
rect 0 9150 4771 9152
rect 0 9120 480 9150
rect 4705 9147 4771 9150
rect 5214 9150 6500 9210
rect 565 9074 631 9077
rect 5214 9074 5274 9150
rect 6494 9148 6500 9150
rect 6564 9210 6570 9212
rect 10041 9210 10107 9213
rect 10501 9210 10567 9213
rect 6564 9150 6792 9210
rect 6564 9148 6570 9150
rect 5533 9076 5599 9077
rect 5993 9076 6059 9077
rect 5533 9074 5580 9076
rect 565 9072 5274 9074
rect 565 9016 570 9072
rect 626 9016 5274 9072
rect 565 9014 5274 9016
rect 5488 9072 5580 9074
rect 5488 9016 5538 9072
rect 5488 9014 5580 9016
rect 565 9011 631 9014
rect 5533 9012 5580 9014
rect 5644 9012 5650 9076
rect 5942 9012 5948 9076
rect 6012 9074 6059 9076
rect 6732 9074 6792 9150
rect 10041 9208 10567 9210
rect 10041 9152 10046 9208
rect 10102 9152 10506 9208
rect 10562 9152 10567 9208
rect 10041 9150 10567 9152
rect 10041 9147 10107 9150
rect 10501 9147 10567 9150
rect 17585 9210 17651 9213
rect 19520 9210 20000 9240
rect 17585 9208 20000 9210
rect 17585 9152 17590 9208
rect 17646 9152 20000 9208
rect 17585 9150 20000 9152
rect 17585 9147 17651 9150
rect 19520 9120 20000 9150
rect 8201 9074 8267 9077
rect 11145 9074 11211 9077
rect 16113 9074 16179 9077
rect 16246 9074 16252 9076
rect 6012 9072 6104 9074
rect 6054 9016 6104 9072
rect 6012 9014 6104 9016
rect 6732 9072 8267 9074
rect 6732 9016 8206 9072
rect 8262 9016 8267 9072
rect 6732 9014 8267 9016
rect 6012 9012 6059 9014
rect 5533 9011 5599 9012
rect 5993 9011 6059 9012
rect 8201 9011 8267 9014
rect 9814 9072 16252 9074
rect 9814 9016 11150 9072
rect 11206 9016 16118 9072
rect 16174 9016 16252 9072
rect 9814 9014 16252 9016
rect 3969 8938 4035 8941
rect 7373 8938 7439 8941
rect 3969 8936 7439 8938
rect 3969 8880 3974 8936
rect 4030 8880 7378 8936
rect 7434 8880 7439 8936
rect 3969 8878 7439 8880
rect 3969 8875 4035 8878
rect 7373 8875 7439 8878
rect 8293 8938 8359 8941
rect 8845 8938 8911 8941
rect 9814 8938 9874 9014
rect 11145 9011 11211 9014
rect 16113 9011 16179 9014
rect 16246 9012 16252 9014
rect 16316 9012 16322 9076
rect 8293 8936 9874 8938
rect 8293 8880 8298 8936
rect 8354 8880 8850 8936
rect 8906 8880 9874 8936
rect 8293 8878 9874 8880
rect 10409 8938 10475 8941
rect 17033 8938 17099 8941
rect 10409 8936 17099 8938
rect 10409 8880 10414 8936
rect 10470 8880 17038 8936
rect 17094 8880 17099 8936
rect 10409 8878 17099 8880
rect 8293 8875 8359 8878
rect 8845 8875 8911 8878
rect 10409 8875 10475 8878
rect 17033 8875 17099 8878
rect 0 8802 480 8832
rect 4889 8804 4955 8805
rect 0 8742 3848 8802
rect 0 8712 480 8742
rect 0 8530 480 8560
rect 565 8530 631 8533
rect 0 8528 631 8530
rect 0 8472 570 8528
rect 626 8472 631 8528
rect 0 8470 631 8472
rect 3788 8530 3848 8742
rect 4838 8740 4844 8804
rect 4908 8802 4955 8804
rect 6545 8802 6611 8805
rect 4908 8800 6611 8802
rect 4950 8744 6550 8800
rect 6606 8744 6611 8800
rect 4908 8742 6611 8744
rect 4908 8740 4955 8742
rect 4889 8739 4955 8740
rect 6545 8739 6611 8742
rect 18321 8802 18387 8805
rect 19520 8802 20000 8832
rect 18321 8800 20000 8802
rect 18321 8744 18326 8800
rect 18382 8744 20000 8800
rect 18321 8742 20000 8744
rect 18321 8739 18387 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 19520 8712 20000 8742
rect 15770 8671 16090 8672
rect 10501 8666 10567 8669
rect 12893 8666 12959 8669
rect 10501 8664 12959 8666
rect 10501 8608 10506 8664
rect 10562 8608 12898 8664
rect 12954 8608 12959 8664
rect 10501 8606 12959 8608
rect 10501 8603 10567 8606
rect 12893 8603 12959 8606
rect 6269 8530 6335 8533
rect 3788 8528 6335 8530
rect 3788 8472 6274 8528
rect 6330 8472 6335 8528
rect 3788 8470 6335 8472
rect 0 8440 480 8470
rect 565 8467 631 8470
rect 6269 8467 6335 8470
rect 6545 8530 6611 8533
rect 15193 8530 15259 8533
rect 19520 8530 20000 8560
rect 6545 8528 15026 8530
rect 6545 8472 6550 8528
rect 6606 8472 15026 8528
rect 6545 8470 15026 8472
rect 6545 8467 6611 8470
rect 3509 8394 3575 8397
rect 4797 8394 4863 8397
rect 3509 8392 4863 8394
rect 3509 8336 3514 8392
rect 3570 8336 4802 8392
rect 4858 8336 4863 8392
rect 3509 8334 4863 8336
rect 3509 8331 3575 8334
rect 4797 8331 4863 8334
rect 6545 8394 6611 8397
rect 6821 8394 6887 8397
rect 6545 8392 6887 8394
rect 6545 8336 6550 8392
rect 6606 8336 6826 8392
rect 6882 8336 6887 8392
rect 6545 8334 6887 8336
rect 6545 8331 6611 8334
rect 6821 8331 6887 8334
rect 8201 8394 8267 8397
rect 14273 8394 14339 8397
rect 8201 8392 14339 8394
rect 8201 8336 8206 8392
rect 8262 8336 14278 8392
rect 14334 8336 14339 8392
rect 8201 8334 14339 8336
rect 14966 8394 15026 8470
rect 15193 8528 20000 8530
rect 15193 8472 15198 8528
rect 15254 8472 20000 8528
rect 15193 8470 20000 8472
rect 15193 8467 15259 8470
rect 19520 8440 20000 8470
rect 15377 8394 15443 8397
rect 16573 8394 16639 8397
rect 14966 8392 16639 8394
rect 14966 8336 15382 8392
rect 15438 8336 16578 8392
rect 16634 8336 16639 8392
rect 14966 8334 16639 8336
rect 8201 8331 8267 8334
rect 14273 8331 14339 8334
rect 15377 8331 15443 8334
rect 16573 8331 16639 8334
rect 10133 8258 10199 8261
rect 11145 8258 11211 8261
rect 10133 8256 11211 8258
rect 10133 8200 10138 8256
rect 10194 8200 11150 8256
rect 11206 8200 11211 8256
rect 10133 8198 11211 8200
rect 10133 8195 10199 8198
rect 11145 8195 11211 8198
rect 11421 8258 11487 8261
rect 11697 8258 11763 8261
rect 12525 8258 12591 8261
rect 11421 8256 12591 8258
rect 11421 8200 11426 8256
rect 11482 8200 11702 8256
rect 11758 8200 12530 8256
rect 12586 8200 12591 8256
rect 11421 8198 12591 8200
rect 11421 8195 11487 8198
rect 11697 8195 11763 8198
rect 12525 8195 12591 8198
rect 6874 8192 7194 8193
rect 0 8122 480 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 1209 8122 1275 8125
rect 0 8120 1275 8122
rect 0 8064 1214 8120
rect 1270 8064 1275 8120
rect 0 8062 1275 8064
rect 0 8032 480 8062
rect 1209 8059 1275 8062
rect 1393 8122 1459 8125
rect 5942 8122 5948 8124
rect 1393 8120 5948 8122
rect 1393 8064 1398 8120
rect 1454 8064 5948 8120
rect 1393 8062 5948 8064
rect 1393 8059 1459 8062
rect 5942 8060 5948 8062
rect 6012 8060 6018 8124
rect 9949 8122 10015 8125
rect 12065 8122 12131 8125
rect 9949 8120 12131 8122
rect 9949 8064 9954 8120
rect 10010 8064 12070 8120
rect 12126 8064 12131 8120
rect 9949 8062 12131 8064
rect 9949 8059 10015 8062
rect 12065 8059 12131 8062
rect 15377 8122 15443 8125
rect 19520 8122 20000 8152
rect 15377 8120 20000 8122
rect 15377 8064 15382 8120
rect 15438 8064 20000 8120
rect 15377 8062 20000 8064
rect 15377 8059 15443 8062
rect 19520 8032 20000 8062
rect 3734 7986 3740 7988
rect 2500 7926 3740 7986
rect 0 7850 480 7880
rect 2500 7850 2560 7926
rect 3734 7924 3740 7926
rect 3804 7924 3810 7988
rect 4705 7986 4771 7989
rect 10869 7986 10935 7989
rect 4705 7984 10935 7986
rect 4705 7928 4710 7984
rect 4766 7928 10874 7984
rect 10930 7928 10935 7984
rect 4705 7926 10935 7928
rect 4705 7923 4771 7926
rect 10869 7923 10935 7926
rect 12341 7984 12407 7989
rect 12341 7928 12346 7984
rect 12402 7928 12407 7984
rect 12341 7923 12407 7928
rect 0 7790 2560 7850
rect 4061 7850 4127 7853
rect 9622 7850 9628 7852
rect 4061 7848 9628 7850
rect 4061 7792 4066 7848
rect 4122 7792 9628 7848
rect 4061 7790 9628 7792
rect 0 7760 480 7790
rect 4061 7787 4127 7790
rect 9622 7788 9628 7790
rect 9692 7850 9698 7852
rect 12344 7850 12404 7923
rect 9692 7790 12404 7850
rect 12985 7850 13051 7853
rect 13353 7850 13419 7853
rect 12985 7848 13419 7850
rect 12985 7792 12990 7848
rect 13046 7792 13358 7848
rect 13414 7792 13419 7848
rect 12985 7790 13419 7792
rect 9692 7788 9698 7790
rect 12985 7787 13051 7790
rect 13353 7787 13419 7790
rect 15469 7850 15535 7853
rect 19520 7850 20000 7880
rect 15469 7848 20000 7850
rect 15469 7792 15474 7848
rect 15530 7792 20000 7848
rect 15469 7790 20000 7792
rect 15469 7787 15535 7790
rect 19520 7760 20000 7790
rect 12249 7714 12315 7717
rect 15285 7714 15351 7717
rect 12249 7712 15351 7714
rect 12249 7656 12254 7712
rect 12310 7656 15290 7712
rect 15346 7656 15351 7712
rect 12249 7654 15351 7656
rect 12249 7651 12315 7654
rect 15285 7651 15351 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 11881 7578 11947 7581
rect 13629 7578 13695 7581
rect 11881 7576 13695 7578
rect 11881 7520 11886 7576
rect 11942 7520 13634 7576
rect 13690 7520 13695 7576
rect 11881 7518 13695 7520
rect 11881 7515 11947 7518
rect 13629 7515 13695 7518
rect 0 7442 480 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 0 7352 480 7382
rect 1301 7379 1367 7382
rect 11789 7442 11855 7445
rect 14089 7442 14155 7445
rect 11789 7440 14155 7442
rect 11789 7384 11794 7440
rect 11850 7384 14094 7440
rect 14150 7384 14155 7440
rect 11789 7382 14155 7384
rect 11789 7379 11855 7382
rect 14089 7379 14155 7382
rect 15561 7442 15627 7445
rect 19520 7442 20000 7472
rect 15561 7440 20000 7442
rect 15561 7384 15566 7440
rect 15622 7384 20000 7440
rect 15561 7382 20000 7384
rect 15561 7379 15627 7382
rect 19520 7352 20000 7382
rect 2405 7306 2471 7309
rect 7557 7306 7623 7309
rect 2405 7304 7623 7306
rect 2405 7248 2410 7304
rect 2466 7248 7562 7304
rect 7618 7248 7623 7304
rect 2405 7246 7623 7248
rect 2405 7243 2471 7246
rect 7557 7243 7623 7246
rect 11789 7306 11855 7309
rect 12157 7306 12223 7309
rect 16573 7306 16639 7309
rect 11789 7304 16639 7306
rect 11789 7248 11794 7304
rect 11850 7248 12162 7304
rect 12218 7248 16578 7304
rect 16634 7248 16639 7304
rect 11789 7246 16639 7248
rect 11789 7243 11855 7246
rect 12157 7243 12223 7246
rect 16573 7243 16639 7246
rect 0 7170 480 7200
rect 5574 7170 5580 7172
rect 0 7110 5580 7170
rect 0 7080 480 7110
rect 5574 7108 5580 7110
rect 5644 7108 5650 7172
rect 7741 7170 7807 7173
rect 12157 7170 12223 7173
rect 7741 7168 12223 7170
rect 7741 7112 7746 7168
rect 7802 7112 12162 7168
rect 12218 7112 12223 7168
rect 7741 7110 12223 7112
rect 7741 7107 7807 7110
rect 12157 7107 12223 7110
rect 16481 7170 16547 7173
rect 19520 7170 20000 7200
rect 16481 7168 20000 7170
rect 16481 7112 16486 7168
rect 16542 7112 20000 7168
rect 16481 7110 20000 7112
rect 16481 7107 16547 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 19520 7080 20000 7110
rect 12805 7039 13125 7040
rect 2865 7034 2931 7037
rect 3182 7034 3188 7036
rect 2865 7032 3188 7034
rect 2865 6976 2870 7032
rect 2926 6976 3188 7032
rect 2865 6974 3188 6976
rect 2865 6971 2931 6974
rect 3182 6972 3188 6974
rect 3252 6972 3258 7036
rect 0 6898 480 6928
rect 2865 6898 2931 6901
rect 0 6896 2931 6898
rect 0 6840 2870 6896
rect 2926 6840 2931 6896
rect 0 6838 2931 6840
rect 0 6808 480 6838
rect 2865 6835 2931 6838
rect 3877 6898 3943 6901
rect 9581 6898 9647 6901
rect 3877 6896 9647 6898
rect 3877 6840 3882 6896
rect 3938 6840 9586 6896
rect 9642 6840 9647 6896
rect 3877 6838 9647 6840
rect 3877 6835 3943 6838
rect 9581 6835 9647 6838
rect 15377 6898 15443 6901
rect 19520 6898 20000 6928
rect 15377 6896 20000 6898
rect 15377 6840 15382 6896
rect 15438 6840 20000 6896
rect 15377 6838 20000 6840
rect 15377 6835 15443 6838
rect 19520 6808 20000 6838
rect 6269 6762 6335 6765
rect 6729 6762 6795 6765
rect 6269 6760 6795 6762
rect 6269 6704 6274 6760
rect 6330 6704 6734 6760
rect 6790 6704 6795 6760
rect 6269 6702 6795 6704
rect 6269 6699 6335 6702
rect 6729 6699 6795 6702
rect 13169 6626 13235 6629
rect 14273 6626 14339 6629
rect 13169 6624 14339 6626
rect 13169 6568 13174 6624
rect 13230 6568 14278 6624
rect 14334 6568 14339 6624
rect 13169 6566 14339 6568
rect 13169 6563 13235 6566
rect 14273 6563 14339 6566
rect 3909 6560 4229 6561
rect 0 6490 480 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 6637 6490 6703 6493
rect 0 6430 3802 6490
rect 0 6400 480 6430
rect 3742 6354 3802 6430
rect 4294 6488 6703 6490
rect 4294 6432 6642 6488
rect 6698 6432 6703 6488
rect 4294 6430 6703 6432
rect 4294 6354 4354 6430
rect 6637 6427 6703 6430
rect 10961 6490 11027 6493
rect 12617 6490 12683 6493
rect 10961 6488 12683 6490
rect 10961 6432 10966 6488
rect 11022 6432 12622 6488
rect 12678 6432 12683 6488
rect 10961 6430 12683 6432
rect 10961 6427 11027 6430
rect 12617 6427 12683 6430
rect 16205 6490 16271 6493
rect 19520 6490 20000 6520
rect 16205 6488 20000 6490
rect 16205 6432 16210 6488
rect 16266 6432 20000 6488
rect 16205 6430 20000 6432
rect 16205 6427 16271 6430
rect 19520 6400 20000 6430
rect 3742 6294 4354 6354
rect 4797 6354 4863 6357
rect 8569 6354 8635 6357
rect 4797 6352 8635 6354
rect 4797 6296 4802 6352
rect 4858 6296 8574 6352
rect 8630 6296 8635 6352
rect 4797 6294 8635 6296
rect 4797 6291 4863 6294
rect 8569 6291 8635 6294
rect 16246 6292 16252 6356
rect 16316 6354 16322 6356
rect 16389 6354 16455 6357
rect 16316 6352 16455 6354
rect 16316 6296 16394 6352
rect 16450 6296 16455 6352
rect 16316 6294 16455 6296
rect 16316 6292 16322 6294
rect 16389 6291 16455 6294
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 18321 6218 18387 6221
rect 19520 6218 20000 6248
rect 18321 6216 20000 6218
rect 18321 6160 18326 6216
rect 18382 6160 20000 6216
rect 18321 6158 20000 6160
rect 18321 6155 18387 6158
rect 19520 6128 20000 6158
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 1761 5946 1827 5949
rect 6637 5946 6703 5949
rect 1761 5944 6703 5946
rect 1761 5888 1766 5944
rect 1822 5888 6642 5944
rect 6698 5888 6703 5944
rect 1761 5886 6703 5888
rect 1761 5883 1827 5886
rect 6637 5883 6703 5886
rect 0 5810 480 5840
rect 2773 5810 2839 5813
rect 0 5808 2839 5810
rect 0 5752 2778 5808
rect 2834 5752 2839 5808
rect 0 5750 2839 5752
rect 0 5720 480 5750
rect 2773 5747 2839 5750
rect 4153 5810 4219 5813
rect 8385 5810 8451 5813
rect 4153 5808 8451 5810
rect 4153 5752 4158 5808
rect 4214 5752 8390 5808
rect 8446 5752 8451 5808
rect 4153 5750 8451 5752
rect 4153 5747 4219 5750
rect 8385 5747 8451 5750
rect 18413 5810 18479 5813
rect 19520 5810 20000 5840
rect 18413 5808 20000 5810
rect 18413 5752 18418 5808
rect 18474 5752 20000 5808
rect 18413 5750 20000 5752
rect 18413 5747 18479 5750
rect 19520 5720 20000 5750
rect 2865 5674 2931 5677
rect 6085 5674 6151 5677
rect 2865 5672 6151 5674
rect 2865 5616 2870 5672
rect 2926 5616 6090 5672
rect 6146 5616 6151 5672
rect 2865 5614 6151 5616
rect 2865 5611 2931 5614
rect 6085 5611 6151 5614
rect 0 5538 480 5568
rect 3693 5538 3759 5541
rect 0 5536 3759 5538
rect 0 5480 3698 5536
rect 3754 5480 3759 5536
rect 0 5478 3759 5480
rect 0 5448 480 5478
rect 3693 5475 3759 5478
rect 4981 5538 5047 5541
rect 6545 5538 6611 5541
rect 8477 5538 8543 5541
rect 4981 5536 8543 5538
rect 4981 5480 4986 5536
rect 5042 5480 6550 5536
rect 6606 5480 8482 5536
rect 8538 5480 8543 5536
rect 4981 5478 8543 5480
rect 4981 5475 5047 5478
rect 6545 5475 6611 5478
rect 8477 5475 8543 5478
rect 18229 5538 18295 5541
rect 19520 5538 20000 5568
rect 18229 5536 20000 5538
rect 18229 5480 18234 5536
rect 18290 5480 20000 5536
rect 18229 5478 20000 5480
rect 18229 5475 18295 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 19520 5448 20000 5478
rect 15770 5407 16090 5408
rect 1669 5402 1735 5405
rect 1669 5400 3434 5402
rect 1669 5344 1674 5400
rect 1730 5344 3434 5400
rect 1669 5342 3434 5344
rect 1669 5339 1735 5342
rect 3233 5266 3299 5269
rect 1350 5264 3299 5266
rect 1350 5208 3238 5264
rect 3294 5208 3299 5264
rect 1350 5206 3299 5208
rect 3374 5266 3434 5342
rect 3693 5266 3759 5269
rect 3374 5264 3759 5266
rect 3374 5208 3698 5264
rect 3754 5208 3759 5264
rect 3374 5206 3759 5208
rect 0 5130 480 5160
rect 1350 5130 1410 5206
rect 3233 5203 3299 5206
rect 3693 5203 3759 5206
rect 0 5070 1410 5130
rect 0 5040 480 5070
rect 3734 5068 3740 5132
rect 3804 5130 3810 5132
rect 4153 5130 4219 5133
rect 3804 5128 4219 5130
rect 3804 5072 4158 5128
rect 4214 5072 4219 5128
rect 3804 5070 4219 5072
rect 3804 5068 3810 5070
rect 4153 5067 4219 5070
rect 16481 5130 16547 5133
rect 19520 5130 20000 5160
rect 16481 5128 20000 5130
rect 16481 5072 16486 5128
rect 16542 5072 20000 5128
rect 16481 5070 20000 5072
rect 16481 5067 16547 5070
rect 19520 5040 20000 5070
rect 1301 4994 1367 4997
rect 6453 4994 6519 4997
rect 1301 4992 6519 4994
rect 1301 4936 1306 4992
rect 1362 4936 6458 4992
rect 6514 4936 6519 4992
rect 1301 4934 6519 4936
rect 1301 4931 1367 4934
rect 6453 4931 6519 4934
rect 14457 4994 14523 4997
rect 17401 4994 17467 4997
rect 14457 4992 17467 4994
rect 14457 4936 14462 4992
rect 14518 4936 17406 4992
rect 17462 4936 17467 4992
rect 14457 4934 17467 4936
rect 14457 4931 14523 4934
rect 17401 4931 17467 4934
rect 6874 4928 7194 4929
rect 0 4858 480 4888
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 4245 4858 4311 4861
rect 0 4856 4311 4858
rect 0 4800 4250 4856
rect 4306 4800 4311 4856
rect 0 4798 4311 4800
rect 0 4768 480 4798
rect 4245 4795 4311 4798
rect 17861 4858 17927 4861
rect 19520 4858 20000 4888
rect 17861 4856 20000 4858
rect 17861 4800 17866 4856
rect 17922 4800 20000 4856
rect 17861 4798 20000 4800
rect 17861 4795 17927 4798
rect 19520 4768 20000 4798
rect 5533 4724 5599 4725
rect 5533 4722 5580 4724
rect 5452 4720 5580 4722
rect 5644 4722 5650 4724
rect 7741 4722 7807 4725
rect 5644 4720 7807 4722
rect 5452 4664 5538 4720
rect 5644 4664 7746 4720
rect 7802 4664 7807 4720
rect 5452 4662 5580 4664
rect 5533 4660 5580 4662
rect 5644 4662 7807 4664
rect 5644 4660 5650 4662
rect 5533 4659 5599 4660
rect 7741 4659 7807 4662
rect 10041 4722 10107 4725
rect 16481 4722 16547 4725
rect 10041 4720 16547 4722
rect 10041 4664 10046 4720
rect 10102 4664 16486 4720
rect 16542 4664 16547 4720
rect 10041 4662 16547 4664
rect 10041 4659 10107 4662
rect 16481 4659 16547 4662
rect 3509 4586 3575 4589
rect 2454 4584 3575 4586
rect 2454 4528 3514 4584
rect 3570 4528 3575 4584
rect 2454 4526 3575 4528
rect 0 4450 480 4480
rect 2454 4450 2514 4526
rect 3509 4523 3575 4526
rect 4245 4586 4311 4589
rect 9581 4586 9647 4589
rect 4245 4584 9647 4586
rect 4245 4528 4250 4584
rect 4306 4528 9586 4584
rect 9642 4528 9647 4584
rect 4245 4526 9647 4528
rect 4245 4523 4311 4526
rect 9581 4523 9647 4526
rect 11329 4586 11395 4589
rect 17033 4586 17099 4589
rect 11329 4584 17099 4586
rect 11329 4528 11334 4584
rect 11390 4528 17038 4584
rect 17094 4528 17099 4584
rect 11329 4526 17099 4528
rect 11329 4523 11395 4526
rect 17033 4523 17099 4526
rect 0 4390 2514 4450
rect 5717 4450 5783 4453
rect 5942 4450 5948 4452
rect 5717 4448 5948 4450
rect 5717 4392 5722 4448
rect 5778 4392 5948 4448
rect 5717 4390 5948 4392
rect 0 4360 480 4390
rect 5717 4387 5783 4390
rect 5942 4388 5948 4390
rect 6012 4450 6018 4452
rect 7925 4450 7991 4453
rect 6012 4448 7991 4450
rect 6012 4392 7930 4448
rect 7986 4392 7991 4448
rect 6012 4390 7991 4392
rect 6012 4388 6018 4390
rect 7925 4387 7991 4390
rect 18321 4450 18387 4453
rect 19520 4450 20000 4480
rect 18321 4448 20000 4450
rect 18321 4392 18326 4448
rect 18382 4392 20000 4448
rect 18321 4390 20000 4392
rect 18321 4387 18387 4390
rect 3909 4384 4229 4385
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19520 4360 20000 4390
rect 15770 4319 16090 4320
rect 5901 4314 5967 4317
rect 7465 4314 7531 4317
rect 5901 4312 7531 4314
rect 5901 4256 5906 4312
rect 5962 4256 7470 4312
rect 7526 4256 7531 4312
rect 5901 4254 7531 4256
rect 5901 4251 5967 4254
rect 7465 4251 7531 4254
rect 0 4178 480 4208
rect 3049 4178 3115 4181
rect 0 4176 3115 4178
rect 0 4120 3054 4176
rect 3110 4120 3115 4176
rect 0 4118 3115 4120
rect 0 4088 480 4118
rect 3049 4115 3115 4118
rect 4061 4178 4127 4181
rect 4705 4178 4771 4181
rect 6545 4180 6611 4181
rect 4061 4176 4771 4178
rect 4061 4120 4066 4176
rect 4122 4120 4710 4176
rect 4766 4120 4771 4176
rect 4061 4118 4771 4120
rect 4061 4115 4127 4118
rect 4705 4115 4771 4118
rect 6494 4116 6500 4180
rect 6564 4178 6611 4180
rect 7005 4178 7071 4181
rect 8293 4178 8359 4181
rect 6564 4176 6656 4178
rect 6606 4120 6656 4176
rect 6564 4118 6656 4120
rect 7005 4176 8359 4178
rect 7005 4120 7010 4176
rect 7066 4120 8298 4176
rect 8354 4120 8359 4176
rect 7005 4118 8359 4120
rect 6564 4116 6611 4118
rect 6545 4115 6611 4116
rect 7005 4115 7071 4118
rect 8293 4115 8359 4118
rect 18229 4178 18295 4181
rect 19520 4178 20000 4208
rect 18229 4176 20000 4178
rect 18229 4120 18234 4176
rect 18290 4120 20000 4176
rect 18229 4118 20000 4120
rect 18229 4115 18295 4118
rect 19520 4088 20000 4118
rect 6177 4044 6243 4045
rect 6126 3980 6132 4044
rect 6196 4042 6243 4044
rect 7649 4042 7715 4045
rect 12157 4042 12223 4045
rect 6196 4040 6288 4042
rect 6238 3984 6288 4040
rect 6196 3982 6288 3984
rect 6456 3982 7482 4042
rect 6196 3980 6243 3982
rect 6177 3979 6243 3980
rect 3366 3844 3372 3908
rect 3436 3906 3442 3908
rect 6456 3906 6516 3982
rect 3436 3846 6516 3906
rect 7422 3906 7482 3982
rect 7649 4040 12223 4042
rect 7649 3984 7654 4040
rect 7710 3984 12162 4040
rect 12218 3984 12223 4040
rect 7649 3982 12223 3984
rect 7649 3979 7715 3982
rect 12157 3979 12223 3982
rect 12433 3906 12499 3909
rect 7422 3904 12499 3906
rect 7422 3848 12438 3904
rect 12494 3848 12499 3904
rect 7422 3846 12499 3848
rect 3436 3844 3442 3846
rect 12433 3843 12499 3846
rect 6874 3840 7194 3841
rect 0 3770 480 3800
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 5901 3770 5967 3773
rect 0 3768 5967 3770
rect 0 3712 5906 3768
rect 5962 3712 5967 3768
rect 0 3710 5967 3712
rect 0 3680 480 3710
rect 5901 3707 5967 3710
rect 18229 3770 18295 3773
rect 19520 3770 20000 3800
rect 18229 3768 20000 3770
rect 18229 3712 18234 3768
rect 18290 3712 20000 3768
rect 18229 3710 20000 3712
rect 18229 3707 18295 3710
rect 19520 3680 20000 3710
rect 1669 3634 1735 3637
rect 17033 3634 17099 3637
rect 1669 3632 17099 3634
rect 1669 3576 1674 3632
rect 1730 3576 17038 3632
rect 17094 3576 17099 3632
rect 1669 3574 17099 3576
rect 1669 3571 1735 3574
rect 17033 3571 17099 3574
rect 0 3498 480 3528
rect 3509 3498 3575 3501
rect 0 3496 3575 3498
rect 0 3440 3514 3496
rect 3570 3440 3575 3496
rect 0 3438 3575 3440
rect 0 3408 480 3438
rect 3509 3435 3575 3438
rect 5901 3498 5967 3501
rect 6126 3498 6132 3500
rect 5901 3496 6132 3498
rect 5901 3440 5906 3496
rect 5962 3440 6132 3496
rect 5901 3438 6132 3440
rect 5901 3435 5967 3438
rect 6126 3436 6132 3438
rect 6196 3436 6202 3500
rect 10593 3498 10659 3501
rect 16113 3498 16179 3501
rect 10593 3496 16179 3498
rect 10593 3440 10598 3496
rect 10654 3440 16118 3496
rect 16174 3440 16179 3496
rect 10593 3438 16179 3440
rect 10593 3435 10659 3438
rect 16113 3435 16179 3438
rect 16297 3498 16363 3501
rect 19520 3498 20000 3528
rect 16297 3496 20000 3498
rect 16297 3440 16302 3496
rect 16358 3440 20000 3496
rect 16297 3438 20000 3440
rect 16297 3435 16363 3438
rect 19520 3408 20000 3438
rect 3909 3296 4229 3297
rect 0 3226 480 3256
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 3417 3226 3483 3229
rect 0 3224 3483 3226
rect 0 3168 3422 3224
rect 3478 3168 3483 3224
rect 0 3166 3483 3168
rect 0 3136 480 3166
rect 3417 3163 3483 3166
rect 10593 3226 10659 3229
rect 14825 3226 14891 3229
rect 10593 3224 14891 3226
rect 10593 3168 10598 3224
rect 10654 3168 14830 3224
rect 14886 3168 14891 3224
rect 10593 3166 14891 3168
rect 10593 3163 10659 3166
rect 14825 3163 14891 3166
rect 16573 3226 16639 3229
rect 19520 3226 20000 3256
rect 16573 3224 20000 3226
rect 16573 3168 16578 3224
rect 16634 3168 20000 3224
rect 16573 3166 20000 3168
rect 16573 3163 16639 3166
rect 19520 3136 20000 3166
rect 3182 3028 3188 3092
rect 3252 3090 3258 3092
rect 3417 3090 3483 3093
rect 3252 3088 3483 3090
rect 3252 3032 3422 3088
rect 3478 3032 3483 3088
rect 3252 3030 3483 3032
rect 3252 3028 3258 3030
rect 3417 3027 3483 3030
rect 6361 3090 6427 3093
rect 9622 3090 9628 3092
rect 6361 3088 9628 3090
rect 6361 3032 6366 3088
rect 6422 3032 9628 3088
rect 6361 3030 9628 3032
rect 6361 3027 6427 3030
rect 9622 3028 9628 3030
rect 9692 3090 9698 3092
rect 10869 3090 10935 3093
rect 9692 3088 10935 3090
rect 9692 3032 10874 3088
rect 10930 3032 10935 3088
rect 9692 3030 10935 3032
rect 9692 3028 9698 3030
rect 10869 3027 10935 3030
rect 5165 2954 5231 2957
rect 16665 2954 16731 2957
rect 5165 2952 16731 2954
rect 5165 2896 5170 2952
rect 5226 2896 16670 2952
rect 16726 2896 16731 2952
rect 5165 2894 16731 2896
rect 5165 2891 5231 2894
rect 16665 2891 16731 2894
rect 0 2818 480 2848
rect 1577 2818 1643 2821
rect 0 2816 1643 2818
rect 0 2760 1582 2816
rect 1638 2760 1643 2816
rect 0 2758 1643 2760
rect 0 2728 480 2758
rect 1577 2755 1643 2758
rect 7557 2818 7623 2821
rect 10501 2818 10567 2821
rect 7557 2816 10567 2818
rect 7557 2760 7562 2816
rect 7618 2760 10506 2816
rect 10562 2760 10567 2816
rect 7557 2758 10567 2760
rect 7557 2755 7623 2758
rect 10501 2755 10567 2758
rect 16849 2818 16915 2821
rect 19520 2818 20000 2848
rect 16849 2816 20000 2818
rect 16849 2760 16854 2816
rect 16910 2760 20000 2816
rect 16849 2758 20000 2760
rect 16849 2755 16915 2758
rect 6874 2752 7194 2753
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 19520 2728 20000 2758
rect 12805 2687 13125 2688
rect 0 2546 480 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 480 2486
rect 4061 2483 4127 2486
rect 17401 2546 17467 2549
rect 19520 2546 20000 2576
rect 17401 2544 20000 2546
rect 17401 2488 17406 2544
rect 17462 2488 20000 2544
rect 17401 2486 20000 2488
rect 17401 2483 17467 2486
rect 19520 2456 20000 2486
rect 3909 2208 4229 2209
rect 0 2138 480 2168
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2143 16090 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 2048 480 2078
rect 2865 2075 2931 2078
rect 16389 2138 16455 2141
rect 19520 2138 20000 2168
rect 16389 2136 20000 2138
rect 16389 2080 16394 2136
rect 16450 2080 20000 2136
rect 16389 2078 20000 2080
rect 16389 2075 16455 2078
rect 19520 2048 20000 2078
rect 0 1866 480 1896
rect 2957 1866 3023 1869
rect 0 1864 3023 1866
rect 0 1808 2962 1864
rect 3018 1808 3023 1864
rect 0 1806 3023 1808
rect 0 1776 480 1806
rect 2957 1803 3023 1806
rect 17125 1866 17191 1869
rect 19520 1866 20000 1896
rect 17125 1864 20000 1866
rect 17125 1808 17130 1864
rect 17186 1808 20000 1864
rect 17125 1806 20000 1808
rect 17125 1803 17191 1806
rect 19520 1776 20000 1806
rect 0 1458 480 1488
rect 3601 1458 3667 1461
rect 0 1456 3667 1458
rect 0 1400 3606 1456
rect 3662 1400 3667 1456
rect 0 1398 3667 1400
rect 0 1368 480 1398
rect 3601 1395 3667 1398
rect 16757 1458 16823 1461
rect 19520 1458 20000 1488
rect 16757 1456 20000 1458
rect 16757 1400 16762 1456
rect 16818 1400 20000 1456
rect 16757 1398 20000 1400
rect 16757 1395 16823 1398
rect 19520 1368 20000 1398
rect 0 1186 480 1216
rect 3509 1186 3575 1189
rect 0 1184 3575 1186
rect 0 1128 3514 1184
rect 3570 1128 3575 1184
rect 0 1126 3575 1128
rect 0 1096 480 1126
rect 3509 1123 3575 1126
rect 17033 1186 17099 1189
rect 19520 1186 20000 1216
rect 17033 1184 20000 1186
rect 17033 1128 17038 1184
rect 17094 1128 20000 1184
rect 17033 1126 20000 1128
rect 17033 1123 17099 1126
rect 19520 1096 20000 1126
rect 0 778 480 808
rect 8109 778 8175 781
rect 0 776 8175 778
rect 0 720 8114 776
rect 8170 720 8175 776
rect 0 718 8175 720
rect 0 688 480 718
rect 8109 715 8175 718
rect 18045 778 18111 781
rect 19520 778 20000 808
rect 18045 776 20000 778
rect 18045 720 18050 776
rect 18106 720 20000 776
rect 18045 718 20000 720
rect 18045 715 18111 718
rect 19520 688 20000 718
rect 0 506 480 536
rect 3141 506 3207 509
rect 0 504 3207 506
rect 0 448 3146 504
rect 3202 448 3207 504
rect 0 446 3207 448
rect 0 416 480 446
rect 3141 443 3207 446
rect 17769 506 17835 509
rect 19520 506 20000 536
rect 17769 504 20000 506
rect 17769 448 17774 504
rect 17830 448 20000 504
rect 17769 446 20000 448
rect 17769 443 17835 446
rect 19520 416 20000 446
rect 0 234 480 264
rect 3417 234 3483 237
rect 0 232 3483 234
rect 0 176 3422 232
rect 3478 176 3483 232
rect 0 174 3483 176
rect 0 144 480 174
rect 3417 171 3483 174
rect 16481 234 16547 237
rect 19520 234 20000 264
rect 16481 232 20000 234
rect 16481 176 16486 232
rect 16542 176 20000 232
rect 16481 174 20000 176
rect 16481 171 16547 174
rect 19520 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 3372 13772 3436 13836
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 10548 13228 10612 13292
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 4844 12276 4908 12340
rect 10364 12276 10428 12340
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3004 11052 3068 11116
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3004 10024 3068 10028
rect 3004 9968 3054 10024
rect 3054 9968 3068 10024
rect 3004 9964 3068 9968
rect 3740 9964 3804 10028
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 10364 9828 10428 9892
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 10548 9752 10612 9756
rect 10548 9696 10598 9752
rect 10598 9696 10612 9752
rect 10548 9692 10612 9696
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 6500 9148 6564 9212
rect 5580 9072 5644 9076
rect 5580 9016 5594 9072
rect 5594 9016 5644 9072
rect 5580 9012 5644 9016
rect 5948 9072 6012 9076
rect 5948 9016 5998 9072
rect 5998 9016 6012 9072
rect 5948 9012 6012 9016
rect 16252 9012 16316 9076
rect 4844 8800 4908 8804
rect 4844 8744 4894 8800
rect 4894 8744 4908 8800
rect 4844 8740 4908 8744
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 5948 8060 6012 8124
rect 3740 7924 3804 7988
rect 9628 7788 9692 7852
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 5580 7108 5644 7172
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3188 6972 3252 7036
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 16252 6292 16316 6356
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 3740 5068 3804 5132
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 5580 4720 5644 4724
rect 5580 4664 5594 4720
rect 5594 4664 5644 4720
rect 5580 4660 5644 4664
rect 5948 4388 6012 4452
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6500 4176 6564 4180
rect 6500 4120 6550 4176
rect 6550 4120 6564 4176
rect 6500 4116 6564 4120
rect 6132 4040 6196 4044
rect 6132 3984 6182 4040
rect 6182 3984 6196 4040
rect 6132 3980 6196 3984
rect 3372 3844 3436 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 6132 3436 6196 3500
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 3188 3028 3252 3092
rect 9628 3028 9692 3092
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3371 13836 3437 13837
rect 3371 13772 3372 13836
rect 3436 13772 3437 13836
rect 3371 13771 3437 13772
rect 3003 11116 3069 11117
rect 3003 11052 3004 11116
rect 3068 11052 3069 11116
rect 3003 11051 3069 11052
rect 3006 10029 3066 11051
rect 3003 10028 3069 10029
rect 3003 9964 3004 10028
rect 3068 9964 3069 10028
rect 3003 9963 3069 9964
rect 3187 7036 3253 7037
rect 3187 6972 3188 7036
rect 3252 6972 3253 7036
rect 3187 6971 3253 6972
rect 3190 3093 3250 6971
rect 3374 3909 3434 13771
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 4843 12340 4909 12341
rect 4843 12276 4844 12340
rect 4908 12276 4909 12340
rect 4843 12275 4909 12276
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3739 10028 3805 10029
rect 3739 9964 3740 10028
rect 3804 9964 3805 10028
rect 3739 9963 3805 9964
rect 3742 7989 3802 9963
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 4846 8805 4906 12275
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6499 9212 6565 9213
rect 6499 9148 6500 9212
rect 6564 9148 6565 9212
rect 6499 9147 6565 9148
rect 5579 9076 5645 9077
rect 5579 9012 5580 9076
rect 5644 9012 5645 9076
rect 5579 9011 5645 9012
rect 5947 9076 6013 9077
rect 5947 9012 5948 9076
rect 6012 9012 6013 9076
rect 5947 9011 6013 9012
rect 4843 8804 4909 8805
rect 4843 8740 4844 8804
rect 4908 8740 4909 8804
rect 4843 8739 4909 8740
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3739 7988 3805 7989
rect 3739 7924 3740 7988
rect 3804 7924 3805 7988
rect 3739 7923 3805 7924
rect 3742 5133 3802 7923
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 5582 7173 5642 9011
rect 5950 8125 6010 9011
rect 5947 8124 6013 8125
rect 5947 8060 5948 8124
rect 6012 8060 6013 8124
rect 5947 8059 6013 8060
rect 5579 7172 5645 7173
rect 5579 7108 5580 7172
rect 5644 7108 5645 7172
rect 5579 7107 5645 7108
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3739 5132 3805 5133
rect 3739 5068 3740 5132
rect 3804 5068 3805 5132
rect 3739 5067 3805 5068
rect 3909 4384 4229 5408
rect 5582 4725 5642 7107
rect 5579 4724 5645 4725
rect 5579 4660 5580 4724
rect 5644 4660 5645 4724
rect 5579 4659 5645 4660
rect 5950 4453 6010 8059
rect 5947 4452 6013 4453
rect 5947 4388 5948 4452
rect 6012 4388 6013 4452
rect 5947 4387 6013 4388
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3371 3908 3437 3909
rect 3371 3844 3372 3908
rect 3436 3844 3437 3908
rect 3371 3843 3437 3844
rect 3909 3296 4229 4320
rect 6502 4181 6562 9147
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 10547 13292 10613 13293
rect 10547 13228 10548 13292
rect 10612 13228 10613 13292
rect 10547 13227 10613 13228
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 10363 12340 10429 12341
rect 10363 12276 10364 12340
rect 10428 12276 10429 12340
rect 10363 12275 10429 12276
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 10366 9893 10426 12275
rect 10363 9892 10429 9893
rect 10363 9828 10364 9892
rect 10428 9828 10429 9892
rect 10363 9827 10429 9828
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 10550 9757 10610 13227
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 10547 9756 10613 9757
rect 10547 9692 10548 9756
rect 10612 9692 10613 9756
rect 10547 9691 10613 9692
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6499 4180 6565 4181
rect 6499 4116 6500 4180
rect 6564 4116 6565 4180
rect 6499 4115 6565 4116
rect 6131 4044 6197 4045
rect 6131 3980 6132 4044
rect 6196 3980 6197 4044
rect 6131 3979 6197 3980
rect 6134 3501 6194 3979
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6131 3500 6197 3501
rect 6131 3436 6132 3500
rect 6196 3436 6197 3500
rect 6131 3435 6197 3436
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3187 3092 3253 3093
rect 3187 3028 3188 3092
rect 3252 3028 3253 3092
rect 3187 3027 3253 3028
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 2752 7195 3776
rect 9630 3093 9690 7787
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 8736 16090 9760
rect 16251 9076 16317 9077
rect 16251 9012 16252 9076
rect 16316 9012 16317 9076
rect 16251 9011 16317 9012
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 16254 6357 16314 9011
rect 16251 6356 16317 6357
rect 16251 6292 16252 6356
rect 16316 6292 16317 6356
rect 16251 6291 16317 6292
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 2208 16090 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1656 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1656 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2668 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4232 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1606821651
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1606821651
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1606821651
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1606821651
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1606821651
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1606821651
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1606821651
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71
timestamp 1606821651
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7544 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7084 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1606821651
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1606821651
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8556 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7912 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10028 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10580 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9568 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606821651
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1606821651
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1606821651
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1606821651
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1606821651
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11040 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11592 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606821651
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14444 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_131 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_143
timestamp 1606821651
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1606821651
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1606821651
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15180 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1606821651
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1606821651
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1606821651
transform 1 0 16744 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1606821651
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1606821651
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1606821651
transform 1 0 17480 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_S_FTB01
timestamp 1606821651
transform 1 0 17204 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606821651
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1606821651
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2116 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1606821651
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_20
timestamp 1606821651
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4600 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3128 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1606821651
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1606821651
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp 1606821651
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7636 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_top_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1606821651
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1606821651
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1606821651
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1606821651
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10948 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11960 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_106
timestamp 1606821651
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1606821651
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13892 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12972 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_127
timestamp 1606821651
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1606821651
transform 1 0 13524 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_S_FTB01
timestamp 1606821651
transform 1 0 16284 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1606821651
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1606821651
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1606821651
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_164
timestamp 1606821651
transform 1 0 16192 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_N_FTB01
timestamp 1606821651
transform 1 0 17756 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1606821651
transform 1 0 17020 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1606821651
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_179
timestamp 1606821651
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1606821651
transform 1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1606821651
transform 1 0 2852 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 3956 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3220 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1606821651
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5612 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1606821651
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1606821651
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 7820 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8372 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1606821651
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1606821651
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10488 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1606821651
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1606821651
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1606821651
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 14260 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1606821651
transform 1 0 13892 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1606821651
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_170
timestamp 1606821651
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606821651
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1606821651
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1932 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1606821651
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1606821651
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1606821651
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1606821651
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6348 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 6072 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1606821651
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 8004 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_73
timestamp 1606821651
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1606821651
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10488 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606821651
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1606821651
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12604 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11500 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_111
timestamp 1606821651
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_122
timestamp 1606821651
transform 1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1606821651
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1606821651
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 18032 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1606821651
transform 1 0 17020 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_171
timestamp 1606821651
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_182
timestamp 1606821651
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1606821651
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2300 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1606821651
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4140 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1606821651
transform 1 0 3772 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606821651
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1606821651
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_82
timestamp 1606821651
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 8924 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1606821651
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1606821651
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606821651
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 13064 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1606821651
transform 1 0 12696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14996 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 14720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1606821651
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1606821651
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_171
timestamp 1606821651
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606821651
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1606821651
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_8
timestamp 1606821651
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606821651
transform 1 0 1472 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 1656 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1606821651
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1606821651
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2024 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2208 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606821651
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 4784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1606821651
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_37
timestamp 1606821651
transform 1 0 4508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 6532 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5888 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 5060 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1606821651
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606821651
transform 1 0 8556 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6992 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7912 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_63
timestamp 1606821651
transform 1 0 6900 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1606821651
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_83
timestamp 1606821651
transform 1 0 8740 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606821651
transform 1 0 10488 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606821651
transform 1 0 8924 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8832 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1606821651
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1606821651
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1606821651
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1606821651
transform 1 0 12328 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_105
timestamp 1606821651
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 12696 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13248 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12788 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13800 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_130
timestamp 1606821651
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1606821651
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15824 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1606821651
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1606821651
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1606821651
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 1606821651
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1606821651
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606821651
transform 1 0 18124 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16468 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16836 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_183
timestamp 1606821651
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1606821651
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp 1606821651
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_188
timestamp 1606821651
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1606821651
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1656 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4508 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1606821651
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1606821651
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_35
timestamp 1606821651
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6256 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 1606821651
transform 1 0 5980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8096 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_72
timestamp 1606821651
transform 1 0 7728 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1606821651
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1606821651
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10856 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_122
timestamp 1606821651
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13524 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1606821651
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15732 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606821651
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1606821651
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1606821651
transform 1 0 17388 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_175
timestamp 1606821651
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1606821651
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1656 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2668 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4692 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1606821651
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1606821651
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_55
timestamp 1606821651
transform 1 0 6164 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606821651
transform 1 0 7820 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1606821651
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_77
timestamp 1606821651
transform 1 0 8188 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_top_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8924 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11040 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp 1606821651
transform 1 0 10764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606821651
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 14260 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 12696 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_130
timestamp 1606821651
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1606821651
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 14812 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_147
timestamp 1606821651
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1606821651
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606821651
transform 1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1606821651
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606821651
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1606821651
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1606821651
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1606821651
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4232 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606821651
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1606821651
transform 1 0 5244 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1606821651
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp 1606821651
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_54
timestamp 1606821651
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606821651
transform 1 0 7268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7820 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1606821651
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_71
timestamp 1606821651
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10304 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1606821651
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_96
timestamp 1606821651
transform 1 0 9936 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1606821651
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12972 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1606821651
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1606821651
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16376 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15364 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606821651
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1606821651
transform 1 0 16192 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17388 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_175
timestamp 1606821651
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1606821651
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2392 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_12
timestamp 1606821651
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606821651
transform 1 0 4048 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1606821651
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_36
timestamp 1606821651
transform 1 0 4416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1606821651
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1606821651
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8280 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1606821651
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1606821651
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9292 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10304 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_87
timestamp 1606821651
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1606821651
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1606821651
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13800 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1606821651
transform 1 0 13432 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14812 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_147
timestamp 1606821651
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_165
timestamp 1606821651
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606821651
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16468 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1606821651
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606821651
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1606821651
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1606821651
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606821651
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_25
timestamp 1606821651
transform 1 0 3404 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5980 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1606821651
transform 1 0 5520 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_52
timestamp 1606821651
transform 1 0 5888 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7912 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1606821651
transform 1 0 7452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1606821651
transform 1 0 7820 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10672 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1606821651
transform 1 0 12144 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1606821651
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15456 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606821651
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1606821651
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16468 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_183
timestamp 1606821651
transform 1 0 17940 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1606821651
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1748 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1606821651
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1606821651
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_25
timestamp 1606821651
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_23
timestamp 1606821651
transform 1 0 3220 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606821651
transform 1 0 3036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1606821651
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_36
timestamp 1606821651
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4600 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606821651
transform 1 0 5060 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5704 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1606821651
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1606821651
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606821651
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1606821651
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_66
timestamp 1606821651
transform 1 0 7176 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1606821651
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9844 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1606821651
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_104
timestamp 1606821651
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11592 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 11316 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 10856 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1606821651
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606821651
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1606821651
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1606821651
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 13248 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1606821651
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1606821651
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1606821651
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606821651
transform 1 0 13708 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1606821651
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15548 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_154
timestamp 1606821651
transform 1 0 15272 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606821651
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1606821651
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_173
timestamp 1606821651
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1606821651
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606821651
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 17940 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_187
timestamp 1606821651
transform 1 0 18308 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1606821651
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606821651
transform 1 0 1472 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1606821651
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1606821651
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4232 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1606821651
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5244 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 1606821651
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1606821651
transform 1 0 6072 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606821651
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7360 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10212 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_84
timestamp 1606821651
transform 1 0 8832 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1606821651
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1606821651
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606821651
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14352 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_top_ipin_0.prog_clk
timestamp 1606821651
transform 1 0 14076 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1606821651
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1606821651
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1606821651
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16560 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1606821651
transform 1 0 17388 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1606821651
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1606821651
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1606821651
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606821651
transform 1 0 3036 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_24
timestamp 1606821651
transform 1 0 3312 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1606821651
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1606821651
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_59
timestamp 1606821651
transform 1 0 6532 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_67
timestamp 1606821651
transform 1 0 7268 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1606821651
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11868 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10856 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_115
timestamp 1606821651
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1606821651
transform 1 0 12696 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15640 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1606821651
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606821651
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17296 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1606821651
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1606821651
transform 1 0 18124 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1606821651
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2024 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1606821651
transform 1 0 1932 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_26
timestamp 1606821651
transform 1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_38
timestamp 1606821651
transform 1 0 4600 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_42
timestamp 1606821651
transform 1 0 4968 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8464 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1606821651
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1606821651
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606821651
transform 1 0 11776 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1606821651
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1606821651
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14352 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13340 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1606821651
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1606821651
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1606821651
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_171
timestamp 1606821651
transform 1 0 16836 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1606821651
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1606821651
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1606821651
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5060 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1606821651
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606821651
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_63
timestamp 1606821651
transform 1 0 6900 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_72
timestamp 1606821651
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1606821651
transform 1 0 10304 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1606821651
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1606821651
transform 1 0 10212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11316 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1606821651
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_120
timestamp 1606821651
transform 1 0 12144 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_132
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1606821651
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15732 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1606821651
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1606821651
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606821651
transform 1 0 18124 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1606821651
transform 1 0 17112 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_168
timestamp 1606821651
transform 1 0 16560 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1606821651
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1606821651
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_10
timestamp 1606821651
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1606821651
transform 1 0 1564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 1656 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1606821651
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606821651
transform 1 0 2300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_17
timestamp 1606821651
transform 1 0 2668 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 3220 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4324 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4876 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1606821651
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_32
timestamp 1606821651
transform 1 0 4048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1606821651
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5888 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_44
timestamp 1606821651
transform 1 0 5152 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606821651
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_50
timestamp 1606821651
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1606821651
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8372 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7912 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_71
timestamp 1606821651
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_83
timestamp 1606821651
transform 1 0 8740 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_72
timestamp 1606821651
transform 1 0 7728 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_78
timestamp 1606821651
transform 1 0 8280 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9844 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10488 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1606821651
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1606821651
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1606821651
transform 1 0 10396 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1606821651
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606821651
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1606821651
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1606821651
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606821651
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_135
timestamp 1606821651
transform 1 0 13524 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1606821651
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1606821651
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_147
timestamp 1606821651
transform 1 0 14628 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606821651
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1606821651
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606821651
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1606821651
transform 1 0 2300 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1606821651
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1606821651
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1606821651
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 3864 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606821651
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1606821651
transform 1 0 3404 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_29
timestamp 1606821651
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_34
timestamp 1606821651
transform 1 0 4232 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1606821651
transform 1 0 5336 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606821651
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_1_N_FTB01
timestamp 1606821651
transform 1 0 8004 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1606821651
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1606821651
transform 1 0 8556 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1606821651
transform 1 0 9660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_105
timestamp 1606821651
transform 1 0 10764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1606821651
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606821651
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1606821651
transform 1 0 14076 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_135
timestamp 1606821651
transform 1 0 13524 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1606821651
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1606821651
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606821651
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606821651
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1606821651
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606821651
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1606821651
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606821651
transform 1 0 2300 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1606821651
transform 1 0 1564 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1606821651
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_17
timestamp 1606821651
transform 1 0 2668 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1606821651
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_40
timestamp 1606821651
transform 1 0 4784 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606821651
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_49
timestamp 1606821651
transform 1 0 5612 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1606821651
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1606821651
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606821651
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1606821651
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1606821651
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1606821651
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1606821651
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1606821651
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606821651
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1606821651
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1606821651
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1606821651
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_180
timestamp 1606821651
transform 1 0 17664 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606821651
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 18234 16520 18290 17000 6 REGIN_FEEDTHROUGH
port 0 nsew default input
rlabel metal3 s 0 16736 480 16856 6 REGOUT_FEEDTHROUGH
port 1 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 SC_IN_BOT
port 2 nsew default input
rlabel metal2 s 1674 16520 1730 17000 6 SC_IN_TOP
port 3 nsew default input
rlabel metal2 s 17590 0 17646 480 6 SC_OUT_BOT
port 4 nsew default tristate
rlabel metal2 s 4986 16520 5042 17000 6 SC_OUT_TOP
port 5 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal2 s 11242 0 11298 480 6 bottom_grid_pin_10_
port 7 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 bottom_grid_pin_11_
port 8 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 bottom_grid_pin_13_
port 10 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 bottom_grid_pin_14_
port 11 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 bottom_grid_pin_15_
port 12 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 bottom_grid_pin_1_
port 13 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 bottom_grid_pin_2_
port 14 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_3_
port 15 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 bottom_grid_pin_4_
port 16 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 bottom_grid_pin_5_
port 17 nsew default tristate
rlabel metal2 s 7562 0 7618 480 6 bottom_grid_pin_6_
port 18 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 bottom_grid_pin_7_
port 19 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 bottom_grid_pin_8_
port 20 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 bottom_grid_pin_9_
port 21 nsew default tristate
rlabel metal2 s 386 0 442 480 6 ccff_head
port 22 nsew default input
rlabel metal2 s 1214 0 1270 480 6 ccff_tail
port 23 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[0]
port 24 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[10]
port 25 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[11]
port 26 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[12]
port 27 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[13]
port 28 nsew default input
rlabel metal3 s 0 11432 480 11552 6 chanx_left_in[14]
port 29 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[15]
port 30 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[16]
port 31 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[17]
port 32 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[18]
port 33 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[19]
port 34 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[1]
port 35 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_left_in[2]
port 36 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[3]
port 37 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[4]
port 38 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[5]
port 39 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[6]
port 40 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[7]
port 41 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[8]
port 42 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[9]
port 43 nsew default input
rlabel metal3 s 0 144 480 264 6 chanx_left_out[0]
port 44 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[10]
port 45 nsew default tristate
rlabel metal3 s 0 3680 480 3800 6 chanx_left_out[11]
port 46 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 chanx_left_out[12]
port 47 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[13]
port 48 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[14]
port 49 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[15]
port 50 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[16]
port 51 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 chanx_left_out[17]
port 52 nsew default tristate
rlabel metal3 s 0 6128 480 6248 6 chanx_left_out[18]
port 53 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 chanx_left_out[19]
port 54 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_out[1]
port 55 nsew default tristate
rlabel metal3 s 0 688 480 808 6 chanx_left_out[2]
port 56 nsew default tristate
rlabel metal3 s 0 1096 480 1216 6 chanx_left_out[3]
port 57 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[4]
port 58 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[5]
port 59 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[6]
port 60 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 chanx_left_out[7]
port 61 nsew default tristate
rlabel metal3 s 0 2728 480 2848 6 chanx_left_out[8]
port 62 nsew default tristate
rlabel metal3 s 0 3136 480 3256 6 chanx_left_out[9]
port 63 nsew default tristate
rlabel metal3 s 19520 10344 20000 10464 6 chanx_right_in[0]
port 64 nsew default input
rlabel metal3 s 19520 13744 20000 13864 6 chanx_right_in[10]
port 65 nsew default input
rlabel metal3 s 19520 14016 20000 14136 6 chanx_right_in[11]
port 66 nsew default input
rlabel metal3 s 19520 14424 20000 14544 6 chanx_right_in[12]
port 67 nsew default input
rlabel metal3 s 19520 14696 20000 14816 6 chanx_right_in[13]
port 68 nsew default input
rlabel metal3 s 19520 15104 20000 15224 6 chanx_right_in[14]
port 69 nsew default input
rlabel metal3 s 19520 15376 20000 15496 6 chanx_right_in[15]
port 70 nsew default input
rlabel metal3 s 19520 15784 20000 15904 6 chanx_right_in[16]
port 71 nsew default input
rlabel metal3 s 19520 16056 20000 16176 6 chanx_right_in[17]
port 72 nsew default input
rlabel metal3 s 19520 16464 20000 16584 6 chanx_right_in[18]
port 73 nsew default input
rlabel metal3 s 19520 16736 20000 16856 6 chanx_right_in[19]
port 74 nsew default input
rlabel metal3 s 19520 10752 20000 10872 6 chanx_right_in[1]
port 75 nsew default input
rlabel metal3 s 19520 11024 20000 11144 6 chanx_right_in[2]
port 76 nsew default input
rlabel metal3 s 19520 11432 20000 11552 6 chanx_right_in[3]
port 77 nsew default input
rlabel metal3 s 19520 11704 20000 11824 6 chanx_right_in[4]
port 78 nsew default input
rlabel metal3 s 19520 12112 20000 12232 6 chanx_right_in[5]
port 79 nsew default input
rlabel metal3 s 19520 12384 20000 12504 6 chanx_right_in[6]
port 80 nsew default input
rlabel metal3 s 19520 12792 20000 12912 6 chanx_right_in[7]
port 81 nsew default input
rlabel metal3 s 19520 13064 20000 13184 6 chanx_right_in[8]
port 82 nsew default input
rlabel metal3 s 19520 13472 20000 13592 6 chanx_right_in[9]
port 83 nsew default input
rlabel metal3 s 19520 3680 20000 3800 6 chanx_right_out[0]
port 84 nsew default tristate
rlabel metal3 s 19520 7080 20000 7200 6 chanx_right_out[10]
port 85 nsew default tristate
rlabel metal3 s 19520 7352 20000 7472 6 chanx_right_out[11]
port 86 nsew default tristate
rlabel metal3 s 19520 7760 20000 7880 6 chanx_right_out[12]
port 87 nsew default tristate
rlabel metal3 s 19520 8032 20000 8152 6 chanx_right_out[13]
port 88 nsew default tristate
rlabel metal3 s 19520 8440 20000 8560 6 chanx_right_out[14]
port 89 nsew default tristate
rlabel metal3 s 19520 8712 20000 8832 6 chanx_right_out[15]
port 90 nsew default tristate
rlabel metal3 s 19520 9120 20000 9240 6 chanx_right_out[16]
port 91 nsew default tristate
rlabel metal3 s 19520 9392 20000 9512 6 chanx_right_out[17]
port 92 nsew default tristate
rlabel metal3 s 19520 9800 20000 9920 6 chanx_right_out[18]
port 93 nsew default tristate
rlabel metal3 s 19520 10072 20000 10192 6 chanx_right_out[19]
port 94 nsew default tristate
rlabel metal3 s 19520 4088 20000 4208 6 chanx_right_out[1]
port 95 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 chanx_right_out[2]
port 96 nsew default tristate
rlabel metal3 s 19520 4768 20000 4888 6 chanx_right_out[3]
port 97 nsew default tristate
rlabel metal3 s 19520 5040 20000 5160 6 chanx_right_out[4]
port 98 nsew default tristate
rlabel metal3 s 19520 5448 20000 5568 6 chanx_right_out[5]
port 99 nsew default tristate
rlabel metal3 s 19520 5720 20000 5840 6 chanx_right_out[6]
port 100 nsew default tristate
rlabel metal3 s 19520 6128 20000 6248 6 chanx_right_out[7]
port 101 nsew default tristate
rlabel metal3 s 19520 6400 20000 6520 6 chanx_right_out[8]
port 102 nsew default tristate
rlabel metal3 s 19520 6808 20000 6928 6 chanx_right_out[9]
port 103 nsew default tristate
rlabel metal3 s 19520 3408 20000 3528 6 clk_1_E_in
port 104 nsew default input
rlabel metal2 s 8298 16520 8354 17000 6 clk_1_N_out
port 105 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 clk_1_S_out
port 106 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 clk_1_W_in
port 107 nsew default input
rlabel metal3 s 19520 3136 20000 3256 6 clk_2_E_in
port 108 nsew default input
rlabel metal3 s 19520 1368 20000 1488 6 clk_2_E_out
port 109 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 clk_2_W_in
port 110 nsew default input
rlabel metal3 s 0 14424 480 14544 6 clk_2_W_out
port 111 nsew default tristate
rlabel metal3 s 19520 2728 20000 2848 6 clk_3_E_in
port 112 nsew default input
rlabel metal3 s 19520 1096 20000 1216 6 clk_3_E_out
port 113 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 clk_3_W_in
port 114 nsew default input
rlabel metal3 s 0 14016 480 14136 6 clk_3_W_out
port 115 nsew default tristate
rlabel metal2 s 11610 16520 11666 17000 6 prog_clk_0_N_in
port 116 nsew default input
rlabel metal2 s 14922 16520 14978 17000 6 prog_clk_0_W_out
port 117 nsew default tristate
rlabel metal3 s 19520 2456 20000 2576 6 prog_clk_1_E_in
port 118 nsew default input
rlabel metal3 s 19520 688 20000 808 6 prog_clk_1_N_out
port 119 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 prog_clk_1_S_out
port 120 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 prog_clk_1_W_in
port 121 nsew default input
rlabel metal3 s 19520 2048 20000 2168 6 prog_clk_2_E_in
port 122 nsew default input
rlabel metal3 s 19520 416 20000 536 6 prog_clk_2_E_out
port 123 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 prog_clk_2_W_in
port 124 nsew default input
rlabel metal3 s 0 13744 480 13864 6 prog_clk_2_W_out
port 125 nsew default tristate
rlabel metal3 s 19520 1776 20000 1896 6 prog_clk_3_E_in
port 126 nsew default input
rlabel metal3 s 19520 144 20000 264 6 prog_clk_3_E_out
port 127 nsew default tristate
rlabel metal3 s 0 14696 480 14816 6 prog_clk_3_W_in
port 128 nsew default input
rlabel metal3 s 0 13472 480 13592 6 prog_clk_3_W_out
port 129 nsew default tristate
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 130 nsew default input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 131 nsew default input
<< properties >>
string FIXED_BBOX 0 0 20000 17000
<< end >>
