* NGSPICE file created from sb_2__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_2__1_ bottom_left_grid_pin_42_ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_
+ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_
+ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ prog_clk_0_N_in top_left_grid_pin_42_ top_left_grid_pin_43_
+ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_
+ top_left_grid_pin_48_ top_left_grid_pin_49_ top_right_grid_pin_1_ VPWR VGND
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_44_ bottom_left_grid_pin_42_
+ mux_bottom_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_062_ VGND VGND VPWR VPWR _062_/HI _062_/LO sky130_fd_sc_hd__conb_1
X_114_ _114_/A VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_061_ VGND VGND VPWR VPWR _061_/HI _061_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _070_/A sky130_fd_sc_hd__buf_4
X_113_ chany_bottom_in[6] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_4
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_35.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_7.mux_l1_in_3_ _045_/HI left_bottom_grid_pin_41_ mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__buf_4
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_15.mux_l3_in_0_ mux_left_track_15.mux_l2_in_1_/X mux_left_track_15.mux_l2_in_0_/X
+ mux_left_track_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l2_in_3_ _047_/HI chanx_left_in[14] mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_mem_bottom_track_1.prog_clk clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_15.mux_l2_in_1_ _064_/HI left_bottom_grid_pin_37_ mux_left_track_15.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_060_ VGND VGND VPWR VPWR _060_/HI _060_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_112_ chany_bottom_in[5] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_7.mux_l2_in_1_ mux_left_track_7.mux_l1_in_3_/X mux_left_track_7.mux_l1_in_2_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_7.mux_l1_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[7] chanx_left_in[0] mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l2_in_0_ chany_bottom_in[19] mux_left_track_15.mux_l1_in_0_/X
+ mux_left_track_15.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_111_ chany_bottom_in[4] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l1_in_1_ left_bottom_grid_pin_35_ chany_bottom_in[6] mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ chany_bottom_in[12] mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[2] top_right_grid_pin_1_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _114_/A sky130_fd_sc_hd__buf_4
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l1_in_0_ chany_bottom_in[12] chany_top_in[12] mux_left_track_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_110_ _110_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_9.mux_l2_in_3_ _060_/HI chanx_left_in[18] mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__buf_4
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_7.mux_l1_in_0_ chany_bottom_in[3] chany_top_in[6] mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ mux_bottom_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_21.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[4] mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_39.mux_l2_in_0_ _043_/HI mux_left_track_39.mux_l1_in_0_/X ccff_tail
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l2_in_1_ _056_/HI mux_bottom_track_25.mux_l1_in_2_/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ chany_top_in[12] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l2_in_1_ bottom_left_grid_pin_49_ bottom_left_grid_pin_45_
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_2_ chanx_left_in[13] chanx_left_in[6] mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_39.mux_l1_in_0_ left_bottom_grid_pin_41_ chany_top_in[1] mux_left_track_39.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
X_098_ _098_/A VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_9.mux_l2_in_0_ bottom_right_grid_pin_1_ mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_43_
+ mux_bottom_track_25.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_3_ _048_/HI chanx_left_in[17] mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _068_/A sky130_fd_sc_hd__buf_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__buf_4
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l1_in_3_ _038_/HI left_bottom_grid_pin_41_ mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_11.mux_l3_in_0_ mux_left_track_11.mux_l2_in_1_/X mux_left_track_11.mux_l2_in_0_/X
+ mux_left_track_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l2_in_1_ mux_top_track_16.mux_l1_in_3_/X mux_top_track_16.mux_l1_in_2_/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_097_ chany_top_in[10] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_1_ _062_/HI left_bottom_grid_pin_35_ mux_left_track_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_ chanx_left_in[10] chanx_left_in[3] mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _090_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_13.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l1_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_096_ chany_top_in[9] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_6_ chanx_left_in[17] chanx_left_in[10] mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_079_ left_bottom_grid_pin_35_ VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__buf_4
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_ chany_bottom_in[11] mux_left_track_11.mux_l1_in_0_/X
+ mux_left_track_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[17] chany_bottom_in[8] mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_1_ left_bottom_grid_pin_35_ chany_bottom_in[4] mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_095_ chany_top_in[8] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_5_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
X_078_ _078_/A VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l1_in_0_ top_left_grid_pin_47_ top_left_grid_pin_43_ mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ chany_bottom_in[9] chany_top_in[9] mux_left_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_23.mux_l2_in_0_ mux_left_track_23.mux_l1_in_1_/X mux_left_track_23.mux_l1_in_0_/X
+ mux_left_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_3_ _059_/HI mux_bottom_track_5.mux_l1_in_6_/X mux_bottom_track_5.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_23.mux_l1_in_1_ _035_/HI left_bottom_grid_pin_41_ mux_left_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_0_ chany_bottom_in[0] chany_top_in[4] mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_19.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_094_ _094_/A VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_4_ bottom_left_grid_pin_48_ bottom_left_grid_pin_47_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_4_/X
+ sky130_fd_sc_hd__mux2_1
X_077_ _077_/A VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ mux_bottom_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_2_ mux_bottom_track_5.mux_l1_in_5_/X mux_bottom_track_5.mux_l1_in_4_/X
+ mux_bottom_track_5.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_23.mux_l1_in_0_ chany_bottom_in[17] chany_top_in[17] mux_left_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_093_ chany_top_in[6] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xmux_left_track_35.mux_l2_in_0_ _041_/HI mux_left_track_35.mux_l1_in_0_/X mux_left_track_35.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_3_ bottom_left_grid_pin_46_ bottom_left_grid_pin_45_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_076_ _076_/A VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_31.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_059_ VGND VGND VPWR VPWR _059_/HI _059_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__buf_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ chany_top_in[5] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_44_ bottom_left_grid_pin_43_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
X_075_ _075_/A VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_29.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_35.mux_l1_in_0_ left_bottom_grid_pin_39_ chany_top_in[7] mux_left_track_35.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ VGND VGND VPWR VPWR _058_/HI _058_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ mux_bottom_track_33.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_37.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _066_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l2_in_1_ _058_/HI mux_bottom_track_33.mux_l1_in_2_/X mux_bottom_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_091_ chany_top_in[4] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ _074_/A VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l1_in_2_ chanx_left_in[14] chanx_left_in[7] mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_42_ bottom_right_grid_pin_1_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ VGND VGND VPWR VPWR _057_/HI _057_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_109_ chany_bottom_in[2] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_35.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__buf_4
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_090_ _090_/A VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__buf_4
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_1_ chanx_left_in[0] bottom_left_grid_pin_48_ mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_073_ _073_/A VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_125_ chany_bottom_in[18] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
X_056_ VGND VGND VPWR VPWR _056_/HI _056_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l1_in_3_ _050_/HI chanx_left_in[16] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
X_108_ _108_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_6_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_2.mux_l2_in_3_ _049_/HI chanx_left_in[13] mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l2_in_1_ mux_top_track_24.mux_l1_in_3_/X mux_top_track_24.mux_l1_in_2_/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_0_ bottom_left_grid_pin_44_ chany_top_in[10] mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_072_ _072_/A VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ chany_bottom_in[17] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ mux_top_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l1_in_2_ chanx_left_in[9] chanx_left_in[2] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_107_ _107_/A VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_1_ _046_/HI left_bottom_grid_pin_34_ mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[13] mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_23.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ _071_/A VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_123_ chany_bottom_in[16] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l1_in_1_ chany_bottom_in[18] chany_bottom_in[9] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_106_ _106_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_1_ _065_/HI left_bottom_grid_pin_38_ mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l2_in_3_ _054_/HI chanx_left_in[15] mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_9.mux_l2_in_0_ chany_bottom_in[8] mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ mux_bottom_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_2.mux_l2_in_1_ chany_bottom_in[4] top_left_grid_pin_49_ mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_070_ _070_/A VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _118_/A sky130_fd_sc_hd__buf_4
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_122_ _122_/A VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l1_in_0_ top_left_grid_pin_48_ top_left_grid_pin_44_ mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_29.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_105_ chany_top_in[18] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_2_ chanx_left_in[8] chanx_left_in[1] mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chany_bottom_in[13] chany_top_in[13] mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_29.mux_l2_in_0_ _037_/HI mux_left_track_29.mux_l1_in_0_/X mux_left_track_29.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_31.mux_l2_in_0_ _039_/HI mux_left_track_31.mux_l1_in_0_/X mux_left_track_31.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l1_in_0_ chany_bottom_in[7] chany_top_in[8] mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_2.mux_l2_in_0_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_121_ chany_bottom_in[14] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_104_ chany_top_in[17] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_1_ bottom_left_grid_pin_49_ mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_29.mux_l1_in_0_ left_bottom_grid_pin_36_ chany_top_in[19] mux_left_track_29.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_31.mux_l1_in_0_ left_bottom_grid_pin_37_ chany_top_in[15] mux_left_track_31.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_120_ chany_bottom_in[13] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
X_103_ chany_top_in[16] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_43_ bottom_right_grid_pin_1_
+ mux_bottom_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_15.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__buf_4
X_102_ _102_/A VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_15.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_101_ chany_top_in[14] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_5.mux_l1_in_3_ _044_/HI left_bottom_grid_pin_40_ mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_13.mux_l3_in_0_ mux_left_track_13.mux_l2_in_1_/X mux_left_track_13.mux_l2_in_0_/X
+ mux_left_track_13.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__buf_4
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_13.mux_l2_in_1_ _063_/HI left_bottom_grid_pin_36_ mux_left_track_13.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_13.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ chany_top_in[13] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_3_ _053_/HI chanx_left_in[18] mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_13.mux_l2_in_0_ chany_bottom_in[15] mux_left_track_13.mux_l1_in_0_/X
+ mux_left_track_13.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_32.mux_l2_in_1_ _051_/HI mux_top_track_32.mux_l1_in_2_/X mux_top_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ mux_top_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_32.mux_l1_in_2_ chanx_left_in[15] chanx_left_in[8] mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_5.mux_l1_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[5] mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_33.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[4] mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_13.mux_l1_in_0_ chany_bottom_in[10] chany_top_in[10] mux_left_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_32.mux_l1_in_1_ chanx_left_in[1] chany_bottom_in[10] mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_0_ chany_bottom_in[1] chany_top_in[5] mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l1_in_1_ _036_/HI left_bottom_grid_pin_34_ mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ chany_top_in[2] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_31.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_1_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_39.mux_l1_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l1_in_0_ top_left_grid_pin_49_ top_left_grid_pin_45_ mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_0_ chany_bottom_in[18] chany_top_in[18] mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_088_ _088_/A VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_37.mux_l2_in_0_ _042_/HI mux_left_track_37.mux_l1_in_0_/X mux_left_track_37.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.mux_l2_in_0_ top_right_grid_pin_1_ mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _098_/A sky130_fd_sc_hd__buf_4
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_37.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _110_/A sky130_fd_sc_hd__buf_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_087_ _087_/A VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_37.mux_l1_in_0_ left_bottom_grid_pin_40_ chany_top_in[3] mux_left_track_37.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ top_left_grid_pin_46_ top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ _086_/A VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _067_/A sky130_fd_sc_hd__buf_4
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ _069_/A VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_6_ chanx_left_in[19] chanx_left_in[12] mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_3_ _061_/HI left_bottom_grid_pin_40_ mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__buf_4
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_085_ _085_/A VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_068_ _068_/A VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_5_ chanx_left_in[5] chany_bottom_in[14] mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XFILLER_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l2_in_3_ _052_/HI mux_top_track_4.mux_l1_in_6_/X mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__buf_4
X_067_ _067_/A VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_119_ chany_bottom_in[12] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xmux_top_track_4.mux_l1_in_4_ chany_bottom_in[5] top_right_grid_pin_1_ mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ mux_top_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[2] mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_083_ _083_/A VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l2_in_2_ mux_top_track_4.mux_l1_in_5_/X mux_top_track_4.mux_l1_in_4_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_066_ _066_/A VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_28_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_118_ _118_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xmux_left_track_19.mux_l2_in_0_ mux_left_track_19.mux_l1_in_1_/X mux_left_track_19.mux_l1_in_0_/X
+ mux_left_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_3_ top_left_grid_pin_49_ top_left_grid_pin_48_ mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_21.mux_l2_in_0_ mux_left_track_21.mux_l1_in_1_/X mux_left_track_21.mux_l1_in_0_/X
+ mux_left_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_19.mux_l1_in_1_ _033_/HI left_bottom_grid_pin_39_ mux_left_track_19.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_3_ _057_/HI chanx_left_in[16] mux_bottom_track_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.mux_l1_in_1_ _034_/HI left_bottom_grid_pin_40_ mux_left_track_21.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[2] chany_top_in[0] mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_082_ _082_/A VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _122_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ mux_bottom_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_065_ VGND VGND VPWR VPWR _065_/HI _065_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_3_5_0_mem_bottom_track_1.prog_clk clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_117_ chany_bottom_in[10] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xmux_top_track_4.mux_l1_in_2_ top_left_grid_pin_47_ top_left_grid_pin_46_ mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_11.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_3_ _055_/HI chanx_left_in[19] mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.mux_l1_in_0_ chany_bottom_in[14] chany_top_in[14] mux_left_track_19.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_2_ chanx_left_in[9] chanx_left_in[2] mux_bottom_track_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.mux_l1_in_0_ chany_bottom_in[16] chany_top_in[16] mux_left_track_21.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l2_in_0_ _040_/HI mux_left_track_33.mux_l1_in_0_/X mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_081_ _081_/A VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__buf_4
X_064_ VGND VGND VPWR VPWR _064_/HI _064_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_1_ mux_bottom_track_17.mux_l1_in_3_/X mux_bottom_track_17.mux_l1_in_2_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_45_ top_left_grid_pin_44_ mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_116_ chany_bottom_in[9] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_2_ chanx_left_in[12] chanx_left_in[5] mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ bottom_left_grid_pin_48_ bottom_left_grid_pin_46_
+ mux_bottom_track_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_080_ _080_/A VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l1_in_0_ left_bottom_grid_pin_38_ chany_top_in[11] mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_063_ VGND VGND VPWR VPWR _063_/HI _063_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_43_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ chany_bottom_in[8] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_42_
+ mux_bottom_track_17.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

