magic
tech sky130A
magscale 1 2
timestamp 1605014177
<< locali >>
rect 7665 33439 7699 33541
rect 12449 31127 12483 31297
rect 4261 29019 4295 29257
rect 10149 23511 10183 23817
rect 10057 12155 10091 12325
rect 6193 9027 6227 9129
rect 6469 6239 6503 6341
<< viali >>
rect 4445 36329 4479 36363
rect 5549 36329 5583 36363
rect 4261 36193 4295 36227
rect 5365 36193 5399 36227
rect 1593 35785 1627 35819
rect 2697 35785 2731 35819
rect 4445 35785 4479 35819
rect 5825 35785 5859 35819
rect 7021 35785 7055 35819
rect 8125 35717 8159 35751
rect 1409 35581 1443 35615
rect 2513 35581 2547 35615
rect 3065 35581 3099 35615
rect 4261 35581 4295 35615
rect 5641 35581 5675 35615
rect 6837 35581 6871 35615
rect 7941 35581 7975 35615
rect 9045 35581 9079 35615
rect 9689 35581 9723 35615
rect 4169 35513 4203 35547
rect 2053 35445 2087 35479
rect 4813 35445 4847 35479
rect 5457 35445 5491 35479
rect 6193 35445 6227 35479
rect 7481 35445 7515 35479
rect 8493 35445 8527 35479
rect 9229 35445 9263 35479
rect 1593 35241 1627 35275
rect 2697 35241 2731 35275
rect 4261 35241 4295 35275
rect 6009 35241 6043 35275
rect 7113 35241 7147 35275
rect 10609 35241 10643 35275
rect 1409 35105 1443 35139
rect 2513 35105 2547 35139
rect 4077 35105 4111 35139
rect 5825 35105 5859 35139
rect 6929 35105 6963 35139
rect 7573 35105 7607 35139
rect 8401 35105 8435 35139
rect 10517 35105 10551 35139
rect 8493 35037 8527 35071
rect 8677 35037 8711 35071
rect 10793 35037 10827 35071
rect 7941 34969 7975 35003
rect 2053 34901 2087 34935
rect 3525 34901 3559 34935
rect 8033 34901 8067 34935
rect 9045 34901 9079 34935
rect 10057 34901 10091 34935
rect 10149 34901 10183 34935
rect 3341 34697 3375 34731
rect 7573 34697 7607 34731
rect 9597 34697 9631 34731
rect 2237 34629 2271 34663
rect 8493 34629 8527 34663
rect 10057 34629 10091 34663
rect 11069 34629 11103 34663
rect 1593 34561 1627 34595
rect 8953 34561 8987 34595
rect 9045 34561 9079 34595
rect 10701 34561 10735 34595
rect 1409 34493 1443 34527
rect 2513 34493 2547 34527
rect 3433 34493 3467 34527
rect 5917 34493 5951 34527
rect 7389 34493 7423 34527
rect 7941 34493 7975 34527
rect 8401 34493 8435 34527
rect 8861 34493 8895 34527
rect 9873 34493 9907 34527
rect 10425 34493 10459 34527
rect 10517 34493 10551 34527
rect 11805 34493 11839 34527
rect 3700 34425 3734 34459
rect 4813 34357 4847 34391
rect 7113 34357 7147 34391
rect 11437 34357 11471 34391
rect 2881 34153 2915 34187
rect 5549 34153 5583 34187
rect 8953 34153 8987 34187
rect 11253 34153 11287 34187
rect 1685 34085 1719 34119
rect 4436 34085 4470 34119
rect 6898 34085 6932 34119
rect 8677 34085 8711 34119
rect 10140 34085 10174 34119
rect 1409 34017 1443 34051
rect 2697 34017 2731 34051
rect 4169 34017 4203 34051
rect 6653 33949 6687 33983
rect 9873 33949 9907 33983
rect 3525 33813 3559 33847
rect 6469 33813 6503 33847
rect 8033 33813 8067 33847
rect 1961 33609 1995 33643
rect 5641 33609 5675 33643
rect 8677 33609 8711 33643
rect 10241 33609 10275 33643
rect 1593 33541 1627 33575
rect 7665 33541 7699 33575
rect 7941 33541 7975 33575
rect 2421 33473 2455 33507
rect 7389 33473 7423 33507
rect 8217 33473 8251 33507
rect 11345 33473 11379 33507
rect 1777 33405 1811 33439
rect 2973 33405 3007 33439
rect 5457 33405 5491 33439
rect 6009 33405 6043 33439
rect 7205 33405 7239 33439
rect 7665 33405 7699 33439
rect 8861 33405 8895 33439
rect 9117 33405 9151 33439
rect 3218 33337 3252 33371
rect 7297 33337 7331 33371
rect 10793 33337 10827 33371
rect 2789 33269 2823 33303
rect 4353 33269 4387 33303
rect 4905 33269 4939 33303
rect 5365 33269 5399 33303
rect 6561 33269 6595 33303
rect 6837 33269 6871 33303
rect 3801 33065 3835 33099
rect 4813 33065 4847 33099
rect 6745 33065 6779 33099
rect 7297 33065 7331 33099
rect 10149 33065 10183 33099
rect 10609 32997 10643 33031
rect 4629 32929 4663 32963
rect 8953 32929 8987 32963
rect 9965 32929 9999 32963
rect 10517 32929 10551 32963
rect 7389 32861 7423 32895
rect 7573 32861 7607 32895
rect 10701 32861 10735 32895
rect 3065 32725 3099 32759
rect 3433 32725 3467 32759
rect 4537 32725 4571 32759
rect 5273 32725 5307 32759
rect 5549 32725 5583 32759
rect 6929 32725 6963 32759
rect 9321 32725 9355 32759
rect 12541 32725 12575 32759
rect 6285 32521 6319 32555
rect 7113 32521 7147 32555
rect 8861 32521 8895 32555
rect 10885 32521 10919 32555
rect 3249 32453 3283 32487
rect 8677 32453 8711 32487
rect 10241 32453 10275 32487
rect 10609 32453 10643 32487
rect 1593 32385 1627 32419
rect 3801 32385 3835 32419
rect 3985 32385 4019 32419
rect 5365 32385 5399 32419
rect 5457 32385 5491 32419
rect 6653 32385 6687 32419
rect 7941 32385 7975 32419
rect 9505 32385 9539 32419
rect 12909 32385 12943 32419
rect 13093 32385 13127 32419
rect 1409 32317 1443 32351
rect 5273 32317 5307 32351
rect 9229 32317 9263 32351
rect 12265 32317 12299 32351
rect 2881 32249 2915 32283
rect 3709 32249 3743 32283
rect 7757 32249 7791 32283
rect 8401 32249 8435 32283
rect 11897 32249 11931 32283
rect 12817 32249 12851 32283
rect 2237 32181 2271 32215
rect 3341 32181 3375 32215
rect 4629 32181 4663 32215
rect 4905 32181 4939 32215
rect 7297 32181 7331 32215
rect 7665 32181 7699 32215
rect 9321 32181 9355 32215
rect 12449 32181 12483 32215
rect 2881 31977 2915 32011
rect 5273 31977 5307 32011
rect 6377 31977 6411 32011
rect 6837 31977 6871 32011
rect 10517 31977 10551 32011
rect 13461 31977 13495 32011
rect 7297 31909 7331 31943
rect 8861 31909 8895 31943
rect 2789 31841 2823 31875
rect 5641 31841 5675 31875
rect 7205 31841 7239 31875
rect 10425 31841 10459 31875
rect 10885 31841 10919 31875
rect 12348 31841 12382 31875
rect 2973 31773 3007 31807
rect 5733 31773 5767 31807
rect 5917 31773 5951 31807
rect 7481 31773 7515 31807
rect 10977 31773 11011 31807
rect 11069 31773 11103 31807
rect 11989 31773 12023 31807
rect 12081 31773 12115 31807
rect 4997 31705 5031 31739
rect 2421 31637 2455 31671
rect 4537 31637 4571 31671
rect 6745 31637 6779 31671
rect 7849 31637 7883 31671
rect 8493 31637 8527 31671
rect 11529 31637 11563 31671
rect 2513 31433 2547 31467
rect 3341 31433 3375 31467
rect 4905 31433 4939 31467
rect 6653 31433 6687 31467
rect 8217 31433 8251 31467
rect 8401 31433 8435 31467
rect 12541 31433 12575 31467
rect 7849 31365 7883 31399
rect 1593 31297 1627 31331
rect 3249 31297 3283 31331
rect 3985 31297 4019 31331
rect 4445 31297 4479 31331
rect 5549 31297 5583 31331
rect 7389 31297 7423 31331
rect 8953 31297 8987 31331
rect 9873 31297 9907 31331
rect 11437 31297 11471 31331
rect 12265 31297 12299 31331
rect 12449 31297 12483 31331
rect 13093 31297 13127 31331
rect 1409 31229 1443 31263
rect 10609 31229 10643 31263
rect 2881 31161 2915 31195
rect 3709 31161 3743 31195
rect 5365 31161 5399 31195
rect 8861 31161 8895 31195
rect 10241 31161 10275 31195
rect 11161 31161 11195 31195
rect 11897 31161 11931 31195
rect 13553 31229 13587 31263
rect 12909 31161 12943 31195
rect 3801 31093 3835 31127
rect 4813 31093 4847 31127
rect 5273 31093 5307 31127
rect 6009 31093 6043 31127
rect 6837 31093 6871 31127
rect 7205 31093 7239 31127
rect 7297 31093 7331 31127
rect 8769 31093 8803 31127
rect 9413 31093 9447 31127
rect 10793 31093 10827 31127
rect 11253 31093 11287 31127
rect 12449 31093 12483 31127
rect 13001 31093 13035 31127
rect 1685 30889 1719 30923
rect 2605 30889 2639 30923
rect 2881 30889 2915 30923
rect 3433 30889 3467 30923
rect 4077 30889 4111 30923
rect 5365 30889 5399 30923
rect 5641 30889 5675 30923
rect 6561 30889 6595 30923
rect 8033 30889 8067 30923
rect 8585 30889 8619 30923
rect 6193 30821 6227 30855
rect 12326 30821 12360 30855
rect 1961 30753 1995 30787
rect 4445 30753 4479 30787
rect 4537 30753 4571 30787
rect 6920 30753 6954 30787
rect 10885 30753 10919 30787
rect 12081 30753 12115 30787
rect 4721 30685 4755 30719
rect 6653 30685 6687 30719
rect 10057 30685 10091 30719
rect 10977 30685 11011 30719
rect 11069 30685 11103 30719
rect 2145 30617 2179 30651
rect 3893 30617 3927 30651
rect 10425 30617 10459 30651
rect 11529 30617 11563 30651
rect 11897 30617 11931 30651
rect 10517 30549 10551 30583
rect 13461 30549 13495 30583
rect 3801 30345 3835 30379
rect 12449 30345 12483 30379
rect 9321 30277 9355 30311
rect 9689 30277 9723 30311
rect 12173 30277 12207 30311
rect 13829 30277 13863 30311
rect 3341 30209 3375 30243
rect 4445 30209 4479 30243
rect 6193 30209 6227 30243
rect 7205 30209 7239 30243
rect 12909 30209 12943 30243
rect 13093 30209 13127 30243
rect 2053 30141 2087 30175
rect 4905 30141 4939 30175
rect 5549 30141 5583 30175
rect 7297 30141 7331 30175
rect 7564 30141 7598 30175
rect 9781 30141 9815 30175
rect 10048 30141 10082 30175
rect 12817 30141 12851 30175
rect 4261 30073 4295 30107
rect 3617 30005 3651 30039
rect 4169 30005 4203 30039
rect 5365 30005 5399 30039
rect 5825 30005 5859 30039
rect 6653 30005 6687 30039
rect 8677 30005 8711 30039
rect 11161 30005 11195 30039
rect 11897 30005 11931 30039
rect 13461 30005 13495 30039
rect 4353 29801 4387 29835
rect 6101 29801 6135 29835
rect 8033 29801 8067 29835
rect 9505 29801 9539 29835
rect 12173 29801 12207 29835
rect 3893 29733 3927 29767
rect 7389 29733 7423 29767
rect 12081 29733 12115 29767
rect 12633 29733 12667 29767
rect 4977 29665 5011 29699
rect 8401 29665 8435 29699
rect 9956 29665 9990 29699
rect 12541 29665 12575 29699
rect 4721 29597 4755 29631
rect 7941 29597 7975 29631
rect 8493 29597 8527 29631
rect 8585 29597 8619 29631
rect 9689 29597 9723 29631
rect 12817 29597 12851 29631
rect 11069 29529 11103 29563
rect 6929 29461 6963 29495
rect 13185 29461 13219 29495
rect 4261 29257 4295 29291
rect 4353 29257 4387 29291
rect 4537 29257 4571 29291
rect 6837 29257 6871 29291
rect 8677 29257 8711 29291
rect 10241 29257 10275 29291
rect 10609 29257 10643 29291
rect 12541 29257 12575 29291
rect 13553 29257 13587 29291
rect 4077 29121 4111 29155
rect 6653 29189 6687 29223
rect 9689 29189 9723 29223
rect 11805 29189 11839 29223
rect 12173 29189 12207 29223
rect 5089 29121 5123 29155
rect 5549 29121 5583 29155
rect 7297 29121 7331 29155
rect 7481 29121 7515 29155
rect 8493 29121 8527 29155
rect 9229 29121 9263 29155
rect 11253 29121 11287 29155
rect 13093 29121 13127 29155
rect 4905 29053 4939 29087
rect 10425 29053 10459 29087
rect 12909 29053 12943 29087
rect 4261 28985 4295 29019
rect 4997 28985 5031 29019
rect 6285 28985 6319 29019
rect 7205 28985 7239 29019
rect 8125 28985 8159 29019
rect 9137 28985 9171 29019
rect 10149 28985 10183 29019
rect 10977 28985 11011 29019
rect 9045 28917 9079 28951
rect 11069 28917 11103 28951
rect 13001 28917 13035 28951
rect 7297 28713 7331 28747
rect 8401 28713 8435 28747
rect 9137 28713 9171 28747
rect 9965 28713 9999 28747
rect 10333 28713 10367 28747
rect 11989 28713 12023 28747
rect 12909 28713 12943 28747
rect 13093 28713 13127 28747
rect 11897 28645 11931 28679
rect 6561 28577 6595 28611
rect 7205 28577 7239 28611
rect 7665 28577 7699 28611
rect 11069 28577 11103 28611
rect 7757 28509 7791 28543
rect 7849 28509 7883 28543
rect 12173 28509 12207 28543
rect 6929 28441 6963 28475
rect 11529 28441 11563 28475
rect 4537 28373 4571 28407
rect 4997 28373 5031 28407
rect 6101 28373 6135 28407
rect 7021 28373 7055 28407
rect 8677 28373 8711 28407
rect 10701 28373 10735 28407
rect 12541 28373 12575 28407
rect 6653 28169 6687 28203
rect 8217 28169 8251 28203
rect 8769 28169 8803 28203
rect 11161 28169 11195 28203
rect 11989 28169 12023 28203
rect 11621 28101 11655 28135
rect 9321 28033 9355 28067
rect 6837 27965 6871 27999
rect 5733 27897 5767 27931
rect 7104 27897 7138 27931
rect 5365 27829 5399 27863
rect 6285 27829 6319 27863
rect 9137 27625 9171 27659
rect 12817 27625 12851 27659
rect 1685 27557 1719 27591
rect 7665 27557 7699 27591
rect 11682 27557 11716 27591
rect 1409 27489 1443 27523
rect 5549 27489 5583 27523
rect 6009 27489 6043 27523
rect 9321 27489 9355 27523
rect 6101 27421 6135 27455
rect 6193 27421 6227 27455
rect 7757 27421 7791 27455
rect 7849 27421 7883 27455
rect 11437 27421 11471 27455
rect 5365 27353 5399 27387
rect 6837 27353 6871 27387
rect 7297 27353 7331 27387
rect 5181 27285 5215 27319
rect 5641 27285 5675 27319
rect 8769 27285 8803 27319
rect 4813 27081 4847 27115
rect 6101 27081 6135 27115
rect 9689 27081 9723 27115
rect 11437 27081 11471 27115
rect 5733 27013 5767 27047
rect 7389 26945 7423 26979
rect 9229 26945 9263 26979
rect 3433 26877 3467 26911
rect 7205 26877 7239 26911
rect 3678 26809 3712 26843
rect 6653 26809 6687 26843
rect 7297 26809 7331 26843
rect 9137 26809 9171 26843
rect 1685 26741 1719 26775
rect 3249 26741 3283 26775
rect 6837 26741 6871 26775
rect 7849 26741 7883 26775
rect 8493 26741 8527 26775
rect 8677 26741 8711 26775
rect 9045 26741 9079 26775
rect 11805 26741 11839 26775
rect 2421 26537 2455 26571
rect 3433 26537 3467 26571
rect 6929 26537 6963 26571
rect 7389 26537 7423 26571
rect 7757 26537 7791 26571
rect 2789 26469 2823 26503
rect 10302 26469 10336 26503
rect 2881 26401 2915 26435
rect 4905 26401 4939 26435
rect 5172 26401 5206 26435
rect 2973 26333 3007 26367
rect 10057 26333 10091 26367
rect 6285 26265 6319 26299
rect 11437 26265 11471 26299
rect 8677 26197 8711 26231
rect 9229 26197 9263 26231
rect 1777 25993 1811 26027
rect 5089 25993 5123 26027
rect 6101 25993 6135 26027
rect 8769 25993 8803 26027
rect 8861 25993 8895 26027
rect 4629 25857 4663 25891
rect 5549 25857 5583 25891
rect 5733 25857 5767 25891
rect 9137 25857 9171 25891
rect 2605 25789 2639 25823
rect 5457 25789 5491 25823
rect 9045 25789 9079 25823
rect 2850 25721 2884 25755
rect 9382 25721 9416 25755
rect 2145 25653 2179 25687
rect 2513 25653 2547 25687
rect 3985 25653 4019 25687
rect 4997 25653 5031 25687
rect 8125 25653 8159 25687
rect 10517 25653 10551 25687
rect 11161 25653 11195 25687
rect 4077 25449 4111 25483
rect 5181 25449 5215 25483
rect 5549 25449 5583 25483
rect 8493 25449 8527 25483
rect 9045 25449 9079 25483
rect 2697 25381 2731 25415
rect 7573 25381 7607 25415
rect 8401 25381 8435 25415
rect 3065 25313 3099 25347
rect 4445 25313 4479 25347
rect 5825 25313 5859 25347
rect 10600 25313 10634 25347
rect 4537 25245 4571 25279
rect 4721 25245 4755 25279
rect 7941 25245 7975 25279
rect 8677 25245 8711 25279
rect 10333 25245 10367 25279
rect 5641 25177 5675 25211
rect 8033 25177 8067 25211
rect 7205 25109 7239 25143
rect 10057 25109 10091 25143
rect 11713 25109 11747 25143
rect 4721 24905 4755 24939
rect 6101 24905 6135 24939
rect 8769 24905 8803 24939
rect 3893 24837 3927 24871
rect 1593 24769 1627 24803
rect 4261 24769 4295 24803
rect 5273 24769 5307 24803
rect 6653 24769 6687 24803
rect 7665 24769 7699 24803
rect 7757 24769 7791 24803
rect 8585 24769 8619 24803
rect 9229 24769 9263 24803
rect 9413 24769 9447 24803
rect 10149 24769 10183 24803
rect 10793 24769 10827 24803
rect 10885 24769 10919 24803
rect 11345 24769 11379 24803
rect 1409 24701 1443 24735
rect 3525 24701 3559 24735
rect 4629 24633 4663 24667
rect 5089 24633 5123 24667
rect 9873 24633 9907 24667
rect 10701 24633 10735 24667
rect 2237 24565 2271 24599
rect 5181 24565 5215 24599
rect 5733 24565 5767 24599
rect 7021 24565 7055 24599
rect 7205 24565 7239 24599
rect 7573 24565 7607 24599
rect 8309 24565 8343 24599
rect 9137 24565 9171 24599
rect 10333 24565 10367 24599
rect 4353 24361 4387 24395
rect 4721 24361 4755 24395
rect 9137 24361 9171 24395
rect 9689 24361 9723 24395
rect 10701 24361 10735 24395
rect 5089 24225 5123 24259
rect 7380 24225 7414 24259
rect 10057 24225 10091 24259
rect 10149 24225 10183 24259
rect 5181 24157 5215 24191
rect 5273 24157 5307 24191
rect 7113 24157 7147 24191
rect 10241 24157 10275 24191
rect 6929 24021 6963 24055
rect 8493 24021 8527 24055
rect 11161 24021 11195 24055
rect 3893 23817 3927 23851
rect 4261 23817 4295 23851
rect 4905 23817 4939 23851
rect 5089 23817 5123 23851
rect 6193 23817 6227 23851
rect 6653 23817 6687 23851
rect 10149 23817 10183 23851
rect 10793 23817 10827 23851
rect 4629 23749 4663 23783
rect 9321 23749 9355 23783
rect 5549 23681 5583 23715
rect 5641 23681 5675 23715
rect 6837 23681 6871 23715
rect 8861 23681 8895 23715
rect 9965 23681 9999 23715
rect 9229 23613 9263 23647
rect 9689 23613 9723 23647
rect 7104 23545 7138 23579
rect 5457 23477 5491 23511
rect 8217 23477 8251 23511
rect 9781 23477 9815 23511
rect 10149 23477 10183 23511
rect 10333 23477 10367 23511
rect 4813 23273 4847 23307
rect 6745 23273 6779 23307
rect 8309 23273 8343 23307
rect 9873 23273 9907 23307
rect 5181 23205 5215 23239
rect 5610 23205 5644 23239
rect 11406 23205 11440 23239
rect 7297 23137 7331 23171
rect 8217 23137 8251 23171
rect 11161 23137 11195 23171
rect 5365 23069 5399 23103
rect 8401 23069 8435 23103
rect 7849 22933 7883 22967
rect 9321 22933 9355 22967
rect 10241 22933 10275 22967
rect 12541 22933 12575 22967
rect 4997 22729 5031 22763
rect 6837 22729 6871 22763
rect 8309 22729 8343 22763
rect 5641 22661 5675 22695
rect 6193 22661 6227 22695
rect 2237 22593 2271 22627
rect 7389 22593 7423 22627
rect 9781 22593 9815 22627
rect 10425 22593 10459 22627
rect 13093 22593 13127 22627
rect 1409 22525 1443 22559
rect 3617 22525 3651 22559
rect 7205 22525 7239 22559
rect 10241 22525 10275 22559
rect 1685 22457 1719 22491
rect 3862 22457 3896 22491
rect 10333 22457 10367 22491
rect 12265 22457 12299 22491
rect 12909 22457 12943 22491
rect 3433 22389 3467 22423
rect 6653 22389 6687 22423
rect 7297 22389 7331 22423
rect 7849 22389 7883 22423
rect 8677 22389 8711 22423
rect 9413 22389 9447 22423
rect 9873 22389 9907 22423
rect 11253 22389 11287 22423
rect 11805 22389 11839 22423
rect 12449 22389 12483 22423
rect 12817 22389 12851 22423
rect 2421 22185 2455 22219
rect 5089 22185 5123 22219
rect 6929 22185 6963 22219
rect 8033 22185 8067 22219
rect 9689 22185 9723 22219
rect 11253 22185 11287 22219
rect 11621 22185 11655 22219
rect 13185 22185 13219 22219
rect 3709 22117 3743 22151
rect 5457 22117 5491 22151
rect 11713 22117 11747 22151
rect 12449 22117 12483 22151
rect 2329 22049 2363 22083
rect 2789 22049 2823 22083
rect 6193 22049 6227 22083
rect 7481 22049 7515 22083
rect 7941 22049 7975 22083
rect 9505 22049 9539 22083
rect 10057 22049 10091 22083
rect 2881 21981 2915 22015
rect 3065 21981 3099 22015
rect 5549 21981 5583 22015
rect 5733 21981 5767 22015
rect 8125 21981 8159 22015
rect 10149 21981 10183 22015
rect 10333 21981 10367 22015
rect 11805 21981 11839 22015
rect 13277 21981 13311 22015
rect 13461 21981 13495 22015
rect 7573 21913 7607 21947
rect 8585 21913 8619 21947
rect 12817 21913 12851 21947
rect 10701 21845 10735 21879
rect 11161 21845 11195 21879
rect 2421 21641 2455 21675
rect 3893 21641 3927 21675
rect 5825 21641 5859 21675
rect 7665 21641 7699 21675
rect 8493 21641 8527 21675
rect 10241 21641 10275 21675
rect 11253 21641 11287 21675
rect 11989 21641 12023 21675
rect 13001 21641 13035 21675
rect 13277 21641 13311 21675
rect 13645 21641 13679 21675
rect 7297 21573 7331 21607
rect 11713 21573 11747 21607
rect 2513 21505 2547 21539
rect 7941 21505 7975 21539
rect 9045 21505 9079 21539
rect 9781 21505 9815 21539
rect 10885 21505 10919 21539
rect 12449 21505 12483 21539
rect 8861 21437 8895 21471
rect 2053 21369 2087 21403
rect 2780 21369 2814 21403
rect 10149 21369 10183 21403
rect 10609 21369 10643 21403
rect 1685 21301 1719 21335
rect 5181 21301 5215 21335
rect 5549 21301 5583 21335
rect 8401 21301 8435 21335
rect 8953 21301 8987 21335
rect 10701 21301 10735 21335
rect 2421 21097 2455 21131
rect 8585 21097 8619 21131
rect 9505 21097 9539 21131
rect 10333 21097 10367 21131
rect 11897 21097 11931 21131
rect 12357 21097 12391 21131
rect 2789 21029 2823 21063
rect 4445 21029 4479 21063
rect 9965 21029 9999 21063
rect 2881 20961 2915 20995
rect 4537 20961 4571 20995
rect 6469 20961 6503 20995
rect 6725 20961 6759 20995
rect 10701 20961 10735 20995
rect 12265 20961 12299 20995
rect 2973 20893 3007 20927
rect 4629 20893 4663 20927
rect 10793 20893 10827 20927
rect 10885 20893 10919 20927
rect 12449 20893 12483 20927
rect 2329 20757 2363 20791
rect 4077 20757 4111 20791
rect 7849 20757 7883 20791
rect 1869 20553 1903 20587
rect 4997 20553 5031 20587
rect 5641 20553 5675 20587
rect 6561 20553 6595 20587
rect 11621 20553 11655 20587
rect 11989 20553 12023 20587
rect 2237 20485 2271 20519
rect 4077 20485 4111 20519
rect 4629 20485 4663 20519
rect 7021 20485 7055 20519
rect 12633 20485 12667 20519
rect 2697 20417 2731 20451
rect 10057 20417 10091 20451
rect 11161 20417 11195 20451
rect 8033 20349 8067 20383
rect 10885 20349 10919 20383
rect 2605 20281 2639 20315
rect 2942 20281 2976 20315
rect 7941 20281 7975 20315
rect 8278 20281 8312 20315
rect 10977 20281 11011 20315
rect 5181 20213 5215 20247
rect 9413 20213 9447 20247
rect 10333 20213 10367 20247
rect 10517 20213 10551 20247
rect 3341 20009 3375 20043
rect 4537 20009 4571 20043
rect 4905 20009 4939 20043
rect 6377 20009 6411 20043
rect 7665 20009 7699 20043
rect 10241 20009 10275 20043
rect 10977 20009 11011 20043
rect 12541 20009 12575 20043
rect 2973 19941 3007 19975
rect 4353 19941 4387 19975
rect 9505 19941 9539 19975
rect 11428 19941 11462 19975
rect 1409 19873 1443 19907
rect 6929 19873 6963 19907
rect 7021 19873 7055 19907
rect 1593 19805 1627 19839
rect 4997 19805 5031 19839
rect 5089 19805 5123 19839
rect 7205 19805 7239 19839
rect 10517 19805 10551 19839
rect 11161 19805 11195 19839
rect 6561 19737 6595 19771
rect 2513 19669 2547 19703
rect 8125 19669 8159 19703
rect 1593 19465 1627 19499
rect 2973 19465 3007 19499
rect 10701 19465 10735 19499
rect 11345 19465 11379 19499
rect 11621 19397 11655 19431
rect 3525 19329 3559 19363
rect 5181 19329 5215 19363
rect 6837 19329 6871 19363
rect 2881 19261 2915 19295
rect 3341 19261 3375 19295
rect 4997 19261 5031 19295
rect 6561 19261 6595 19295
rect 7104 19261 7138 19295
rect 9321 19261 9355 19295
rect 4537 19193 4571 19227
rect 6285 19193 6319 19227
rect 9566 19193 9600 19227
rect 3433 19125 3467 19159
rect 4169 19125 4203 19159
rect 4629 19125 4663 19159
rect 5089 19125 5123 19159
rect 5641 19125 5675 19159
rect 8217 19125 8251 19159
rect 9137 19125 9171 19159
rect 4997 18921 5031 18955
rect 5733 18921 5767 18955
rect 6653 18921 6687 18955
rect 9321 18921 9355 18955
rect 10425 18921 10459 18955
rect 10885 18921 10919 18955
rect 4721 18853 4755 18887
rect 5641 18785 5675 18819
rect 6837 18785 6871 18819
rect 10793 18785 10827 18819
rect 5917 18717 5951 18751
rect 11069 18717 11103 18751
rect 3065 18581 3099 18615
rect 5273 18581 5307 18615
rect 8125 18581 8159 18615
rect 3065 18377 3099 18411
rect 4721 18377 4755 18411
rect 6561 18377 6595 18411
rect 10517 18377 10551 18411
rect 11161 18377 11195 18411
rect 5089 18309 5123 18343
rect 3617 18241 3651 18275
rect 5641 18241 5675 18275
rect 5733 18241 5767 18275
rect 7481 18241 7515 18275
rect 2973 18173 3007 18207
rect 3433 18173 3467 18207
rect 7205 18173 7239 18207
rect 2605 18105 2639 18139
rect 5549 18105 5583 18139
rect 3525 18037 3559 18071
rect 4353 18037 4387 18071
rect 5181 18037 5215 18071
rect 6193 18037 6227 18071
rect 6837 18037 6871 18071
rect 7297 18037 7331 18071
rect 8125 18037 8159 18071
rect 9137 18037 9171 18071
rect 10885 18037 10919 18071
rect 3157 17833 3191 17867
rect 5457 17833 5491 17867
rect 6009 17833 6043 17867
rect 7297 17833 7331 17867
rect 7941 17833 7975 17867
rect 8493 17833 8527 17867
rect 9689 17833 9723 17867
rect 8401 17765 8435 17799
rect 3801 17697 3835 17731
rect 4344 17697 4378 17731
rect 10057 17697 10091 17731
rect 10149 17697 10183 17731
rect 4077 17629 4111 17663
rect 8585 17629 8619 17663
rect 10241 17629 10275 17663
rect 6929 17493 6963 17527
rect 8033 17493 8067 17527
rect 3709 17289 3743 17323
rect 5273 17289 5307 17323
rect 5641 17289 5675 17323
rect 8953 17289 8987 17323
rect 9965 17289 9999 17323
rect 3617 17153 3651 17187
rect 4169 17153 4203 17187
rect 4353 17153 4387 17187
rect 7297 17153 7331 17187
rect 7941 17153 7975 17187
rect 8493 17153 8527 17187
rect 9597 17153 9631 17187
rect 7757 17085 7791 17119
rect 9321 17085 9355 17119
rect 4077 17017 4111 17051
rect 6653 17017 6687 17051
rect 7849 17017 7883 17051
rect 3249 16949 3283 16983
rect 4813 16949 4847 16983
rect 7389 16949 7423 16983
rect 8861 16949 8895 16983
rect 9413 16949 9447 16983
rect 10425 16949 10459 16983
rect 3801 16745 3835 16779
rect 5181 16745 5215 16779
rect 7573 16745 7607 16779
rect 8585 16745 8619 16779
rect 9045 16745 9079 16779
rect 1685 16677 1719 16711
rect 2973 16677 3007 16711
rect 7113 16677 7147 16711
rect 1409 16609 1443 16643
rect 2686 16609 2720 16643
rect 5089 16609 5123 16643
rect 6745 16609 6779 16643
rect 7481 16609 7515 16643
rect 7941 16609 7975 16643
rect 8033 16609 8067 16643
rect 10241 16609 10275 16643
rect 11069 16609 11103 16643
rect 11336 16609 11370 16643
rect 5273 16541 5307 16575
rect 8217 16541 8251 16575
rect 4721 16473 4755 16507
rect 9965 16473 9999 16507
rect 4353 16405 4387 16439
rect 12449 16405 12483 16439
rect 1593 16201 1627 16235
rect 2789 16201 2823 16235
rect 6193 16201 6227 16235
rect 8493 16201 8527 16235
rect 9045 16201 9079 16235
rect 9505 16065 9539 16099
rect 3433 15997 3467 16031
rect 4261 15997 4295 16031
rect 7113 15997 7147 16031
rect 9597 15997 9631 16031
rect 9864 15997 9898 16031
rect 4528 15929 4562 15963
rect 7380 15929 7414 15963
rect 11621 15929 11655 15963
rect 3801 15861 3835 15895
rect 4169 15861 4203 15895
rect 5641 15861 5675 15895
rect 6653 15861 6687 15895
rect 10977 15861 11011 15895
rect 11897 15861 11931 15895
rect 5457 15657 5491 15691
rect 7573 15657 7607 15691
rect 7665 15657 7699 15691
rect 8125 15657 8159 15691
rect 9689 15657 9723 15691
rect 11437 15657 11471 15691
rect 8033 15589 8067 15623
rect 4333 15521 4367 15555
rect 7205 15521 7239 15555
rect 10057 15521 10091 15555
rect 11877 15521 11911 15555
rect 4077 15453 4111 15487
rect 6561 15453 6595 15487
rect 8217 15453 8251 15487
rect 10149 15453 10183 15487
rect 10333 15453 10367 15487
rect 11621 15453 11655 15487
rect 9137 15317 9171 15351
rect 13001 15317 13035 15351
rect 4169 15113 4203 15147
rect 5181 15113 5215 15147
rect 7849 15113 7883 15147
rect 8309 15113 8343 15147
rect 10517 15113 10551 15147
rect 11069 15113 11103 15147
rect 11529 15113 11563 15147
rect 12173 15113 12207 15147
rect 6837 15045 6871 15079
rect 5089 14977 5123 15011
rect 5825 14977 5859 15011
rect 7389 14977 7423 15011
rect 13001 14977 13035 15011
rect 4721 14909 4755 14943
rect 5549 14909 5583 14943
rect 6285 14909 6319 14943
rect 7205 14909 7239 14943
rect 9137 14909 9171 14943
rect 9045 14841 9079 14875
rect 9404 14841 9438 14875
rect 11897 14841 11931 14875
rect 12817 14841 12851 14875
rect 3801 14773 3835 14807
rect 5641 14773 5675 14807
rect 6561 14773 6595 14807
rect 7297 14773 7331 14807
rect 12449 14773 12483 14807
rect 12909 14773 12943 14807
rect 7297 14569 7331 14603
rect 7941 14569 7975 14603
rect 8861 14569 8895 14603
rect 9505 14569 9539 14603
rect 11621 14569 11655 14603
rect 12081 14569 12115 14603
rect 12725 14569 12759 14603
rect 13277 14569 13311 14603
rect 1685 14501 1719 14535
rect 1409 14433 1443 14467
rect 6184 14433 6218 14467
rect 10517 14433 10551 14467
rect 10609 14433 10643 14467
rect 5917 14365 5951 14399
rect 10701 14365 10735 14399
rect 12173 14365 12207 14399
rect 12265 14365 12299 14399
rect 9965 14297 9999 14331
rect 11713 14297 11747 14331
rect 5273 14229 5307 14263
rect 10149 14229 10183 14263
rect 11161 14229 11195 14263
rect 6837 14025 6871 14059
rect 8585 14025 8619 14059
rect 8769 14025 8803 14059
rect 10609 14025 10643 14059
rect 11805 14025 11839 14059
rect 12449 14025 12483 14059
rect 13461 14025 13495 14059
rect 1685 13957 1719 13991
rect 6561 13957 6595 13991
rect 10241 13957 10275 13991
rect 5917 13889 5951 13923
rect 6193 13889 6227 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 11161 13889 11195 13923
rect 13001 13889 13035 13923
rect 5549 13821 5583 13855
rect 9873 13821 9907 13855
rect 12909 13821 12943 13855
rect 7205 13753 7239 13787
rect 9137 13753 9171 13787
rect 10977 13753 11011 13787
rect 12817 13753 12851 13787
rect 11069 13685 11103 13719
rect 12265 13685 12299 13719
rect 6929 13481 6963 13515
rect 8861 13481 8895 13515
rect 10701 13481 10735 13515
rect 10885 13481 10919 13515
rect 11253 13481 11287 13515
rect 10241 13413 10275 13447
rect 11897 13413 11931 13447
rect 12541 13413 12575 13447
rect 11345 13277 11379 13311
rect 11529 13277 11563 13311
rect 7941 13141 7975 13175
rect 10241 12937 10275 12971
rect 10977 12937 11011 12971
rect 11621 12937 11655 12971
rect 7941 12733 7975 12767
rect 7849 12665 7883 12699
rect 8186 12665 8220 12699
rect 11345 12665 11379 12699
rect 9321 12597 9355 12631
rect 10057 12325 10091 12359
rect 4629 12257 4663 12291
rect 7941 12257 7975 12291
rect 8401 12257 8435 12291
rect 3893 12189 3927 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 9689 12189 9723 12223
rect 10609 12257 10643 12291
rect 10885 12257 10919 12291
rect 11417 12257 11451 12291
rect 11161 12189 11195 12223
rect 10057 12121 10091 12155
rect 10149 12121 10183 12155
rect 10701 12121 10735 12155
rect 4261 12053 4295 12087
rect 8033 12053 8067 12087
rect 12541 12053 12575 12087
rect 3801 11849 3835 11883
rect 10149 11849 10183 11883
rect 11253 11849 11287 11883
rect 12449 11849 12483 11883
rect 9965 11781 9999 11815
rect 1593 11713 1627 11747
rect 4169 11713 4203 11747
rect 7665 11713 7699 11747
rect 10701 11713 10735 11747
rect 12173 11713 12207 11747
rect 13001 11713 13035 11747
rect 1409 11645 1443 11679
rect 4261 11645 4295 11679
rect 4517 11645 4551 11679
rect 7573 11645 7607 11679
rect 7932 11645 7966 11679
rect 9689 11645 9723 11679
rect 2237 11577 2271 11611
rect 3433 11577 3467 11611
rect 7205 11577 7239 11611
rect 10609 11577 10643 11611
rect 12909 11577 12943 11611
rect 5641 11509 5675 11543
rect 9045 11509 9079 11543
rect 10517 11509 10551 11543
rect 11805 11509 11839 11543
rect 12817 11509 12851 11543
rect 4813 11305 4847 11339
rect 7757 11305 7791 11339
rect 8125 11305 8159 11339
rect 8769 11305 8803 11339
rect 11069 11305 11103 11339
rect 12541 11305 12575 11339
rect 3893 11237 3927 11271
rect 7113 11237 7147 11271
rect 7665 11237 7699 11271
rect 11621 11237 11655 11271
rect 4537 11169 4571 11203
rect 4997 11169 5031 11203
rect 5089 11169 5123 11203
rect 5356 11169 5390 11203
rect 9956 11169 9990 11203
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 9689 11101 9723 11135
rect 3065 10965 3099 10999
rect 6469 10965 6503 10999
rect 4537 10761 4571 10795
rect 5917 10761 5951 10795
rect 8769 10761 8803 10795
rect 9413 10761 9447 10795
rect 10609 10761 10643 10795
rect 6561 10693 6595 10727
rect 9689 10693 9723 10727
rect 10517 10693 10551 10727
rect 2881 10625 2915 10659
rect 3525 10625 3559 10659
rect 5089 10625 5123 10659
rect 11253 10625 11287 10659
rect 3433 10557 3467 10591
rect 6837 10557 6871 10591
rect 7093 10557 7127 10591
rect 11069 10557 11103 10591
rect 4997 10489 5031 10523
rect 2973 10421 3007 10455
rect 3341 10421 3375 10455
rect 3985 10421 4019 10455
rect 4445 10421 4479 10455
rect 4905 10421 4939 10455
rect 5641 10421 5675 10455
rect 8217 10421 8251 10455
rect 10149 10421 10183 10455
rect 10977 10421 11011 10455
rect 3065 10217 3099 10251
rect 5089 10217 5123 10251
rect 7573 10217 7607 10251
rect 7941 10217 7975 10251
rect 8309 10217 8343 10251
rect 8585 10217 8619 10251
rect 10057 10217 10091 10251
rect 10149 10217 10183 10251
rect 10793 10217 10827 10251
rect 7205 10149 7239 10183
rect 5457 10081 5491 10115
rect 8769 10081 8803 10115
rect 4629 10013 4663 10047
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 6653 10013 6687 10047
rect 10333 10013 10367 10047
rect 9689 9945 9723 9979
rect 4997 9877 5031 9911
rect 4353 9673 4387 9707
rect 6193 9673 6227 9707
rect 8585 9673 8619 9707
rect 10057 9673 10091 9707
rect 9781 9605 9815 9639
rect 5733 9537 5767 9571
rect 6653 9537 6687 9571
rect 7573 9537 7607 9571
rect 8493 9537 8527 9571
rect 9137 9537 9171 9571
rect 4721 9469 4755 9503
rect 5641 9469 5675 9503
rect 7389 9469 7423 9503
rect 5089 9401 5123 9435
rect 8033 9401 8067 9435
rect 9045 9401 9079 9435
rect 5181 9333 5215 9367
rect 5549 9333 5583 9367
rect 7021 9333 7055 9367
rect 7481 9333 7515 9367
rect 8953 9333 8987 9367
rect 10517 9333 10551 9367
rect 4353 9129 4387 9163
rect 5733 9129 5767 9163
rect 6193 9129 6227 9163
rect 6469 9129 6503 9163
rect 9045 9129 9079 9163
rect 5457 9061 5491 9095
rect 7012 9061 7046 9095
rect 4721 8993 4755 9027
rect 6101 8993 6135 9027
rect 6193 8993 6227 9027
rect 4813 8925 4847 8959
rect 4905 8925 4939 8959
rect 6745 8925 6779 8959
rect 5917 8789 5951 8823
rect 8125 8789 8159 8823
rect 8677 8789 8711 8823
rect 10057 8789 10091 8823
rect 4445 8585 4479 8619
rect 5181 8585 5215 8619
rect 9137 8585 9171 8619
rect 7941 8517 7975 8551
rect 5733 8449 5767 8483
rect 6193 8449 6227 8483
rect 7389 8449 7423 8483
rect 7573 8449 7607 8483
rect 9505 8449 9539 8483
rect 10609 8449 10643 8483
rect 2421 8381 2455 8415
rect 5549 8381 5583 8415
rect 5641 8381 5675 8415
rect 6653 8381 6687 8415
rect 7297 8381 7331 8415
rect 8493 8381 8527 8415
rect 9781 8381 9815 8415
rect 10333 8381 10367 8415
rect 2329 8313 2363 8347
rect 2666 8313 2700 8347
rect 5089 8313 5123 8347
rect 10425 8313 10459 8347
rect 3801 8245 3835 8279
rect 6929 8245 6963 8279
rect 8401 8245 8435 8279
rect 8677 8245 8711 8279
rect 9597 8245 9631 8279
rect 9965 8245 9999 8279
rect 4445 8041 4479 8075
rect 4813 8041 4847 8075
rect 6377 8041 6411 8075
rect 7021 8041 7055 8075
rect 7481 8041 7515 8075
rect 8033 8041 8067 8075
rect 9045 8041 9079 8075
rect 10057 8041 10091 8075
rect 11989 8041 12023 8075
rect 1685 7973 1719 8007
rect 7389 7973 7423 8007
rect 10333 7973 10367 8007
rect 1409 7905 1443 7939
rect 5264 7905 5298 7939
rect 7665 7905 7699 7939
rect 8401 7905 8435 7939
rect 10876 7905 10910 7939
rect 4997 7837 5031 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 10609 7837 10643 7871
rect 2513 7701 2547 7735
rect 3341 7701 3375 7735
rect 2421 7497 2455 7531
rect 3157 7497 3191 7531
rect 6285 7497 6319 7531
rect 11805 7497 11839 7531
rect 6561 7429 6595 7463
rect 7389 7429 7423 7463
rect 8953 7361 8987 7395
rect 9781 7361 9815 7395
rect 1409 7293 1443 7327
rect 3249 7293 3283 7327
rect 3516 7293 3550 7327
rect 6837 7293 6871 7327
rect 8677 7293 8711 7327
rect 9873 7293 9907 7327
rect 10140 7293 10174 7327
rect 5549 7225 5583 7259
rect 8769 7225 8803 7259
rect 12173 7225 12207 7259
rect 1593 7157 1627 7191
rect 2053 7157 2087 7191
rect 4629 7157 4663 7191
rect 5181 7157 5215 7191
rect 7021 7157 7055 7191
rect 7849 7157 7883 7191
rect 8125 7157 8159 7191
rect 8309 7157 8343 7191
rect 9413 7157 9447 7191
rect 11253 7157 11287 7191
rect 4629 6953 4663 6987
rect 4997 6953 5031 6987
rect 6469 6953 6503 6987
rect 8033 6953 8067 6987
rect 9505 6953 9539 6987
rect 12541 6953 12575 6987
rect 6929 6885 6963 6919
rect 8401 6885 8435 6919
rect 12633 6885 12667 6919
rect 1409 6817 1443 6851
rect 3617 6817 3651 6851
rect 3893 6817 3927 6851
rect 5089 6817 5123 6851
rect 6377 6817 6411 6851
rect 6837 6817 6871 6851
rect 9137 6817 9171 6851
rect 9956 6817 9990 6851
rect 4353 6749 4387 6783
rect 5181 6749 5215 6783
rect 7021 6749 7055 6783
rect 7849 6749 7883 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 9689 6749 9723 6783
rect 12725 6749 12759 6783
rect 12173 6681 12207 6715
rect 1593 6613 1627 6647
rect 1961 6613 1995 6647
rect 2421 6613 2455 6647
rect 3249 6613 3283 6647
rect 3709 6613 3743 6647
rect 7573 6613 7607 6647
rect 11069 6613 11103 6647
rect 11989 6613 12023 6647
rect 4261 6409 4295 6443
rect 5457 6409 5491 6443
rect 5917 6409 5951 6443
rect 8677 6409 8711 6443
rect 9781 6409 9815 6443
rect 10057 6409 10091 6443
rect 11805 6409 11839 6443
rect 13461 6409 13495 6443
rect 3341 6341 3375 6375
rect 6469 6341 6503 6375
rect 6561 6341 6595 6375
rect 8585 6341 8619 6375
rect 1593 6273 1627 6307
rect 4905 6273 4939 6307
rect 6285 6273 6319 6307
rect 7665 6273 7699 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 1409 6205 1443 6239
rect 2685 6205 2719 6239
rect 3893 6205 3927 6239
rect 4813 6205 4847 6239
rect 6469 6205 6503 6239
rect 7481 6205 7515 6239
rect 8125 6205 8159 6239
rect 10241 6205 10275 6239
rect 10793 6205 10827 6239
rect 12265 6205 12299 6239
rect 2237 6137 2271 6171
rect 4721 6137 4755 6171
rect 7573 6137 7607 6171
rect 9045 6137 9079 6171
rect 11161 6137 11195 6171
rect 13829 6137 13863 6171
rect 2513 6069 2547 6103
rect 2881 6069 2915 6103
rect 4353 6069 4387 6103
rect 7113 6069 7147 6103
rect 10425 6069 10459 6103
rect 11345 6069 11379 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 3341 5865 3375 5899
rect 4629 5865 4663 5899
rect 5181 5865 5215 5899
rect 6561 5865 6595 5899
rect 7205 5865 7239 5899
rect 8125 5865 8159 5899
rect 8953 5865 8987 5899
rect 12081 5865 12115 5899
rect 12817 5865 12851 5899
rect 3617 5797 3651 5831
rect 1409 5729 1443 5763
rect 2697 5729 2731 5763
rect 4077 5729 4111 5763
rect 5549 5729 5583 5763
rect 5641 5729 5675 5763
rect 7113 5729 7147 5763
rect 8309 5729 8343 5763
rect 9689 5729 9723 5763
rect 13277 5729 13311 5763
rect 1593 5661 1627 5695
rect 5733 5661 5767 5695
rect 7297 5661 7331 5695
rect 12173 5661 12207 5695
rect 12265 5661 12299 5695
rect 2513 5593 2547 5627
rect 9873 5593 9907 5627
rect 10333 5593 10367 5627
rect 11713 5593 11747 5627
rect 2881 5525 2915 5559
rect 4261 5525 4295 5559
rect 4997 5525 5031 5559
rect 6745 5525 6779 5559
rect 8493 5525 8527 5559
rect 10609 5525 10643 5559
rect 13461 5525 13495 5559
rect 1961 5321 1995 5355
rect 2973 5321 3007 5355
rect 4905 5321 4939 5355
rect 8401 5321 8435 5355
rect 9229 5321 9263 5355
rect 9689 5321 9723 5355
rect 11805 5321 11839 5355
rect 12173 5321 12207 5355
rect 13001 5321 13035 5355
rect 13369 5321 13403 5355
rect 1869 5253 1903 5287
rect 5917 5253 5951 5287
rect 2421 5185 2455 5219
rect 2605 5185 2639 5219
rect 3525 5185 3559 5219
rect 7573 5185 7607 5219
rect 10793 5185 10827 5219
rect 2329 5117 2363 5151
rect 5549 5117 5583 5151
rect 8585 5117 8619 5151
rect 12449 5117 12483 5151
rect 3433 5049 3467 5083
rect 3770 5049 3804 5083
rect 7389 5049 7423 5083
rect 10057 5049 10091 5083
rect 6285 4981 6319 5015
rect 6561 4981 6595 5015
rect 7021 4981 7055 5015
rect 7481 4981 7515 5015
rect 8769 4981 8803 5015
rect 10149 4981 10183 5015
rect 10517 4981 10551 5015
rect 10609 4981 10643 5015
rect 11345 4981 11379 5015
rect 12633 4981 12667 5015
rect 2421 4777 2455 4811
rect 4261 4777 4295 4811
rect 4445 4777 4479 4811
rect 6009 4777 6043 4811
rect 6469 4777 6503 4811
rect 7021 4777 7055 4811
rect 7481 4777 7515 4811
rect 10701 4777 10735 4811
rect 11069 4777 11103 4811
rect 2329 4709 2363 4743
rect 4905 4709 4939 4743
rect 5917 4709 5951 4743
rect 8033 4709 8067 4743
rect 2789 4641 2823 4675
rect 4813 4641 4847 4675
rect 6377 4641 6411 4675
rect 7941 4641 7975 4675
rect 9505 4641 9539 4675
rect 10057 4641 10091 4675
rect 11509 4641 11543 4675
rect 1961 4573 1995 4607
rect 2881 4573 2915 4607
rect 2973 4573 3007 4607
rect 5089 4573 5123 4607
rect 5457 4573 5491 4607
rect 6561 4573 6595 4607
rect 8125 4573 8159 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 11253 4573 11287 4607
rect 7573 4505 7607 4539
rect 8953 4505 8987 4539
rect 3525 4437 3559 4471
rect 3893 4437 3927 4471
rect 8585 4437 8619 4471
rect 9689 4437 9723 4471
rect 12633 4437 12667 4471
rect 2329 4233 2363 4267
rect 4353 4233 4387 4267
rect 5365 4233 5399 4267
rect 6101 4233 6135 4267
rect 7481 4233 7515 4267
rect 9781 4233 9815 4267
rect 11621 4233 11655 4267
rect 11989 4233 12023 4267
rect 2789 4165 2823 4199
rect 4261 4165 4295 4199
rect 3341 4097 3375 4131
rect 4813 4097 4847 4131
rect 4997 4097 5031 4131
rect 8033 4097 8067 4131
rect 8861 4097 8895 4131
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 13001 4097 13035 4131
rect 1409 4029 1443 4063
rect 4721 4029 4755 4063
rect 7389 4029 7423 4063
rect 7849 4029 7883 4063
rect 9045 4029 9079 4063
rect 10425 4029 10459 4063
rect 12449 4029 12483 4063
rect 1685 3961 1719 3995
rect 3157 3961 3191 3995
rect 3893 3961 3927 3995
rect 7941 3961 7975 3995
rect 8585 3961 8619 3995
rect 2697 3893 2731 3927
rect 3249 3893 3283 3927
rect 6561 3893 6595 3927
rect 10057 3893 10091 3927
rect 11345 3893 11379 3927
rect 12633 3893 12667 3927
rect 2421 3689 2455 3723
rect 4537 3689 4571 3723
rect 5089 3689 5123 3723
rect 5733 3689 5767 3723
rect 6101 3689 6135 3723
rect 7665 3689 7699 3723
rect 9505 3689 9539 3723
rect 10609 3689 10643 3723
rect 12449 3689 12483 3723
rect 1685 3621 1719 3655
rect 2789 3621 2823 3655
rect 6552 3621 6586 3655
rect 10333 3621 10367 3655
rect 4445 3553 4479 3587
rect 9689 3553 9723 3587
rect 11069 3553 11103 3587
rect 11325 3553 11359 3587
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 3433 3485 3467 3519
rect 3893 3485 3927 3519
rect 4629 3485 4663 3519
rect 6285 3485 6319 3519
rect 13553 3485 13587 3519
rect 8309 3417 8343 3451
rect 2329 3349 2363 3383
rect 4077 3349 4111 3383
rect 8585 3349 8619 3383
rect 8953 3349 8987 3383
rect 9873 3349 9907 3383
rect 2513 3145 2547 3179
rect 3525 3145 3559 3179
rect 5457 3145 5491 3179
rect 6377 3145 6411 3179
rect 7113 3145 7147 3179
rect 8585 3145 8619 3179
rect 9137 3145 9171 3179
rect 9597 3145 9631 3179
rect 11805 3145 11839 3179
rect 12449 3145 12483 3179
rect 3157 3077 3191 3111
rect 3893 3077 3927 3111
rect 11069 3077 11103 3111
rect 2789 3009 2823 3043
rect 13093 3009 13127 3043
rect 1434 2941 1468 2975
rect 2973 2941 3007 2975
rect 4077 2941 4111 2975
rect 7205 2941 7239 2975
rect 7461 2941 7495 2975
rect 9689 2941 9723 2975
rect 9945 2941 9979 2975
rect 12817 2941 12851 2975
rect 12909 2941 12943 2975
rect 4344 2873 4378 2907
rect 12265 2873 12299 2907
rect 1593 2805 1627 2839
rect 1961 2805 1995 2839
rect 13461 2805 13495 2839
rect 2881 2601 2915 2635
rect 3525 2601 3559 2635
rect 4445 2601 4479 2635
rect 5089 2601 5123 2635
rect 5457 2601 5491 2635
rect 7205 2601 7239 2635
rect 8493 2601 8527 2635
rect 10241 2601 10275 2635
rect 12449 2601 12483 2635
rect 12633 2601 12667 2635
rect 3893 2533 3927 2567
rect 4537 2533 4571 2567
rect 6561 2533 6595 2567
rect 13093 2533 13127 2567
rect 1757 2465 1791 2499
rect 5641 2465 5675 2499
rect 7481 2465 7515 2499
rect 8033 2465 8067 2499
rect 8585 2465 8619 2499
rect 9597 2465 9631 2499
rect 10609 2465 10643 2499
rect 11989 2465 12023 2499
rect 13001 2465 13035 2499
rect 1501 2397 1535 2431
rect 4721 2397 4755 2431
rect 9229 2397 9263 2431
rect 10149 2397 10183 2431
rect 10701 2397 10735 2431
rect 10885 2397 10919 2431
rect 11345 2397 11379 2431
rect 11713 2397 11747 2431
rect 13277 2397 13311 2431
rect 13645 2397 13679 2431
rect 4077 2329 4111 2363
rect 6285 2329 6319 2363
rect 5825 2261 5859 2295
rect 7665 2261 7699 2295
rect 8769 2261 8803 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 4433 36363 4491 36369
rect 4433 36329 4445 36363
rect 4479 36360 4491 36363
rect 4522 36360 4528 36372
rect 4479 36332 4528 36360
rect 4479 36329 4491 36332
rect 4433 36323 4491 36329
rect 4522 36320 4528 36332
rect 4580 36320 4586 36372
rect 5534 36360 5540 36372
rect 5495 36332 5540 36360
rect 5534 36320 5540 36332
rect 5592 36320 5598 36372
rect 4246 36224 4252 36236
rect 4207 36196 4252 36224
rect 4246 36184 4252 36196
rect 4304 36184 4310 36236
rect 5353 36227 5411 36233
rect 5353 36193 5365 36227
rect 5399 36224 5411 36227
rect 5442 36224 5448 36236
rect 5399 36196 5448 36224
rect 5399 36193 5411 36196
rect 5353 36187 5411 36193
rect 5442 36184 5448 36196
rect 5500 36184 5506 36236
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 566 35776 572 35828
rect 624 35816 630 35828
rect 1581 35819 1639 35825
rect 1581 35816 1593 35819
rect 624 35788 1593 35816
rect 624 35776 630 35788
rect 1581 35785 1593 35788
rect 1627 35785 1639 35819
rect 1581 35779 1639 35785
rect 2590 35776 2596 35828
rect 2648 35816 2654 35828
rect 2685 35819 2743 35825
rect 2685 35816 2697 35819
rect 2648 35788 2697 35816
rect 2648 35776 2654 35788
rect 2685 35785 2697 35788
rect 2731 35785 2743 35819
rect 2685 35779 2743 35785
rect 3970 35776 3976 35828
rect 4028 35816 4034 35828
rect 4433 35819 4491 35825
rect 4433 35816 4445 35819
rect 4028 35788 4445 35816
rect 4028 35776 4034 35788
rect 4433 35785 4445 35788
rect 4479 35785 4491 35819
rect 4433 35779 4491 35785
rect 5813 35819 5871 35825
rect 5813 35785 5825 35819
rect 5859 35816 5871 35819
rect 6178 35816 6184 35828
rect 5859 35788 6184 35816
rect 5859 35785 5871 35788
rect 5813 35779 5871 35785
rect 6178 35776 6184 35788
rect 6236 35776 6242 35828
rect 6914 35776 6920 35828
rect 6972 35816 6978 35828
rect 7009 35819 7067 35825
rect 7009 35816 7021 35819
rect 6972 35788 7021 35816
rect 6972 35776 6978 35788
rect 7009 35785 7021 35788
rect 7055 35785 7067 35819
rect 7009 35779 7067 35785
rect 8018 35708 8024 35760
rect 8076 35748 8082 35760
rect 8113 35751 8171 35757
rect 8113 35748 8125 35751
rect 8076 35720 8125 35748
rect 8076 35708 8082 35720
rect 8113 35717 8125 35720
rect 8159 35717 8171 35751
rect 8113 35711 8171 35717
rect 1397 35615 1455 35621
rect 1397 35581 1409 35615
rect 1443 35612 1455 35615
rect 2501 35615 2559 35621
rect 1443 35584 2084 35612
rect 1443 35581 1455 35584
rect 1397 35575 1455 35581
rect 2056 35485 2084 35584
rect 2501 35581 2513 35615
rect 2547 35612 2559 35615
rect 3053 35615 3111 35621
rect 3053 35612 3065 35615
rect 2547 35584 3065 35612
rect 2547 35581 2559 35584
rect 2501 35575 2559 35581
rect 3053 35581 3065 35584
rect 3099 35612 3111 35615
rect 3234 35612 3240 35624
rect 3099 35584 3240 35612
rect 3099 35581 3111 35584
rect 3053 35575 3111 35581
rect 3234 35572 3240 35584
rect 3292 35572 3298 35624
rect 4249 35615 4307 35621
rect 4249 35581 4261 35615
rect 4295 35612 4307 35615
rect 5629 35615 5687 35621
rect 4295 35584 4329 35612
rect 4295 35581 4307 35584
rect 4249 35575 4307 35581
rect 5629 35581 5641 35615
rect 5675 35612 5687 35615
rect 6825 35615 6883 35621
rect 5675 35584 6040 35612
rect 5675 35581 5687 35584
rect 5629 35575 5687 35581
rect 4157 35547 4215 35553
rect 4157 35513 4169 35547
rect 4203 35544 4215 35547
rect 4264 35544 4292 35575
rect 5534 35544 5540 35556
rect 4203 35516 5540 35544
rect 4203 35513 4215 35516
rect 4157 35507 4215 35513
rect 5534 35504 5540 35516
rect 5592 35504 5598 35556
rect 6012 35488 6040 35584
rect 6825 35581 6837 35615
rect 6871 35612 6883 35615
rect 7929 35615 7987 35621
rect 6871 35584 7512 35612
rect 6871 35581 6883 35584
rect 6825 35575 6883 35581
rect 7484 35488 7512 35584
rect 7929 35581 7941 35615
rect 7975 35612 7987 35615
rect 9033 35615 9091 35621
rect 7975 35584 8340 35612
rect 7975 35581 7987 35584
rect 7929 35575 7987 35581
rect 8312 35488 8340 35584
rect 9033 35581 9045 35615
rect 9079 35612 9091 35615
rect 9677 35615 9735 35621
rect 9677 35612 9689 35615
rect 9079 35584 9689 35612
rect 9079 35581 9091 35584
rect 9033 35575 9091 35581
rect 9677 35581 9689 35584
rect 9723 35612 9735 35615
rect 10318 35612 10324 35624
rect 9723 35584 10324 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 10318 35572 10324 35584
rect 10376 35572 10382 35624
rect 2041 35479 2099 35485
rect 2041 35445 2053 35479
rect 2087 35476 2099 35479
rect 2222 35476 2228 35488
rect 2087 35448 2228 35476
rect 2087 35445 2099 35448
rect 2041 35439 2099 35445
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 4246 35436 4252 35488
rect 4304 35476 4310 35488
rect 4801 35479 4859 35485
rect 4801 35476 4813 35479
rect 4304 35448 4813 35476
rect 4304 35436 4310 35448
rect 4801 35445 4813 35448
rect 4847 35445 4859 35479
rect 5442 35476 5448 35488
rect 5403 35448 5448 35476
rect 4801 35439 4859 35445
rect 5442 35436 5448 35448
rect 5500 35436 5506 35488
rect 5994 35436 6000 35488
rect 6052 35476 6058 35488
rect 6181 35479 6239 35485
rect 6181 35476 6193 35479
rect 6052 35448 6193 35476
rect 6052 35436 6058 35448
rect 6181 35445 6193 35448
rect 6227 35445 6239 35479
rect 7466 35476 7472 35488
rect 7427 35448 7472 35476
rect 6181 35439 6239 35445
rect 7466 35436 7472 35448
rect 7524 35436 7530 35488
rect 8294 35436 8300 35488
rect 8352 35476 8358 35488
rect 8481 35479 8539 35485
rect 8481 35476 8493 35479
rect 8352 35448 8493 35476
rect 8352 35436 8358 35448
rect 8481 35445 8493 35448
rect 8527 35445 8539 35479
rect 9214 35476 9220 35488
rect 9175 35448 9220 35476
rect 8481 35439 8539 35445
rect 9214 35436 9220 35448
rect 9272 35436 9278 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 198 35232 204 35284
rect 256 35272 262 35284
rect 1581 35275 1639 35281
rect 1581 35272 1593 35275
rect 256 35244 1593 35272
rect 256 35232 262 35244
rect 1581 35241 1593 35244
rect 1627 35241 1639 35275
rect 1581 35235 1639 35241
rect 2130 35232 2136 35284
rect 2188 35272 2194 35284
rect 2685 35275 2743 35281
rect 2685 35272 2697 35275
rect 2188 35244 2697 35272
rect 2188 35232 2194 35244
rect 2685 35241 2697 35244
rect 2731 35241 2743 35275
rect 2685 35235 2743 35241
rect 4154 35232 4160 35284
rect 4212 35272 4218 35284
rect 4249 35275 4307 35281
rect 4249 35272 4261 35275
rect 4212 35244 4261 35272
rect 4212 35232 4218 35244
rect 4249 35241 4261 35244
rect 4295 35241 4307 35275
rect 4249 35235 4307 35241
rect 5997 35275 6055 35281
rect 5997 35241 6009 35275
rect 6043 35272 6055 35275
rect 6638 35272 6644 35284
rect 6043 35244 6644 35272
rect 6043 35241 6055 35244
rect 5997 35235 6055 35241
rect 6638 35232 6644 35244
rect 6696 35232 6702 35284
rect 7101 35275 7159 35281
rect 7101 35241 7113 35275
rect 7147 35272 7159 35275
rect 7742 35272 7748 35284
rect 7147 35244 7748 35272
rect 7147 35241 7159 35244
rect 7101 35235 7159 35241
rect 7742 35232 7748 35244
rect 7800 35232 7806 35284
rect 10134 35232 10140 35284
rect 10192 35272 10198 35284
rect 10597 35275 10655 35281
rect 10597 35272 10609 35275
rect 10192 35244 10609 35272
rect 10192 35232 10198 35244
rect 10597 35241 10609 35244
rect 10643 35272 10655 35275
rect 15378 35272 15384 35284
rect 10643 35244 15384 35272
rect 10643 35241 10655 35244
rect 10597 35235 10655 35241
rect 15378 35232 15384 35244
rect 15436 35232 15442 35284
rect 1397 35139 1455 35145
rect 1397 35105 1409 35139
rect 1443 35136 1455 35139
rect 1854 35136 1860 35148
rect 1443 35108 1860 35136
rect 1443 35105 1455 35108
rect 1397 35099 1455 35105
rect 1854 35096 1860 35108
rect 1912 35096 1918 35148
rect 2498 35136 2504 35148
rect 2459 35108 2504 35136
rect 2498 35096 2504 35108
rect 2556 35096 2562 35148
rect 4062 35136 4068 35148
rect 4023 35108 4068 35136
rect 4062 35096 4068 35108
rect 4120 35096 4126 35148
rect 5813 35139 5871 35145
rect 5813 35105 5825 35139
rect 5859 35136 5871 35139
rect 6178 35136 6184 35148
rect 5859 35108 6184 35136
rect 5859 35105 5871 35108
rect 5813 35099 5871 35105
rect 6178 35096 6184 35108
rect 6236 35096 6242 35148
rect 6914 35136 6920 35148
rect 6875 35108 6920 35136
rect 6914 35096 6920 35108
rect 6972 35096 6978 35148
rect 7561 35139 7619 35145
rect 7561 35105 7573 35139
rect 7607 35136 7619 35139
rect 8386 35136 8392 35148
rect 7607 35108 8392 35136
rect 7607 35105 7619 35108
rect 7561 35099 7619 35105
rect 8386 35096 8392 35108
rect 8444 35096 8450 35148
rect 10505 35139 10563 35145
rect 10505 35105 10517 35139
rect 10551 35136 10563 35139
rect 10962 35136 10968 35148
rect 10551 35108 10968 35136
rect 10551 35105 10563 35108
rect 10505 35099 10563 35105
rect 10962 35096 10968 35108
rect 11020 35096 11026 35148
rect 8481 35071 8539 35077
rect 8481 35037 8493 35071
rect 8527 35037 8539 35071
rect 8662 35068 8668 35080
rect 8623 35040 8668 35068
rect 8481 35031 8539 35037
rect 7926 35000 7932 35012
rect 7887 34972 7932 35000
rect 7926 34960 7932 34972
rect 7984 35000 7990 35012
rect 8496 35000 8524 35031
rect 8662 35028 8668 35040
rect 8720 35028 8726 35080
rect 10778 35068 10784 35080
rect 10739 35040 10784 35068
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 7984 34972 8524 35000
rect 7984 34960 7990 34972
rect 2038 34932 2044 34944
rect 1999 34904 2044 34932
rect 2038 34892 2044 34904
rect 2096 34892 2102 34944
rect 3510 34932 3516 34944
rect 3471 34904 3516 34932
rect 3510 34892 3516 34904
rect 3568 34892 3574 34944
rect 8018 34932 8024 34944
rect 7979 34904 8024 34932
rect 8018 34892 8024 34904
rect 8076 34892 8082 34944
rect 8846 34892 8852 34944
rect 8904 34932 8910 34944
rect 9033 34935 9091 34941
rect 9033 34932 9045 34935
rect 8904 34904 9045 34932
rect 8904 34892 8910 34904
rect 9033 34901 9045 34904
rect 9079 34901 9091 34935
rect 9033 34895 9091 34901
rect 10045 34935 10103 34941
rect 10045 34901 10057 34935
rect 10091 34932 10103 34935
rect 10137 34935 10195 34941
rect 10137 34932 10149 34935
rect 10091 34904 10149 34932
rect 10091 34901 10103 34904
rect 10045 34895 10103 34901
rect 10137 34901 10149 34904
rect 10183 34932 10195 34935
rect 10410 34932 10416 34944
rect 10183 34904 10416 34932
rect 10183 34901 10195 34904
rect 10137 34895 10195 34901
rect 10410 34892 10416 34904
rect 10468 34892 10474 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 3329 34731 3387 34737
rect 3329 34697 3341 34731
rect 3375 34728 3387 34731
rect 4062 34728 4068 34740
rect 3375 34700 4068 34728
rect 3375 34697 3387 34700
rect 3329 34691 3387 34697
rect 4062 34688 4068 34700
rect 4120 34688 4126 34740
rect 7374 34688 7380 34740
rect 7432 34728 7438 34740
rect 7561 34731 7619 34737
rect 7561 34728 7573 34731
rect 7432 34700 7573 34728
rect 7432 34688 7438 34700
rect 7561 34697 7573 34700
rect 7607 34697 7619 34731
rect 7561 34691 7619 34697
rect 9585 34731 9643 34737
rect 9585 34697 9597 34731
rect 9631 34728 9643 34731
rect 10962 34728 10968 34740
rect 9631 34700 10968 34728
rect 9631 34697 9643 34700
rect 9585 34691 9643 34697
rect 10962 34688 10968 34700
rect 11020 34688 11026 34740
rect 1854 34620 1860 34672
rect 1912 34660 1918 34672
rect 2225 34663 2283 34669
rect 2225 34660 2237 34663
rect 1912 34632 2237 34660
rect 1912 34620 1918 34632
rect 2225 34629 2237 34632
rect 2271 34660 2283 34663
rect 2590 34660 2596 34672
rect 2271 34632 2596 34660
rect 2271 34629 2283 34632
rect 2225 34623 2283 34629
rect 2590 34620 2596 34632
rect 2648 34620 2654 34672
rect 8478 34660 8484 34672
rect 8439 34632 8484 34660
rect 8478 34620 8484 34632
rect 8536 34620 8542 34672
rect 8846 34620 8852 34672
rect 8904 34660 8910 34672
rect 10045 34663 10103 34669
rect 10045 34660 10057 34663
rect 8904 34632 10057 34660
rect 8904 34620 8910 34632
rect 10045 34629 10057 34632
rect 10091 34629 10103 34663
rect 10045 34623 10103 34629
rect 10778 34620 10784 34672
rect 10836 34660 10842 34672
rect 11057 34663 11115 34669
rect 11057 34660 11069 34663
rect 10836 34632 11069 34660
rect 10836 34620 10842 34632
rect 11057 34629 11069 34632
rect 11103 34629 11115 34663
rect 11057 34623 11115 34629
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 8018 34552 8024 34604
rect 8076 34592 8082 34604
rect 8938 34592 8944 34604
rect 8076 34564 8944 34592
rect 8076 34552 8082 34564
rect 8938 34552 8944 34564
rect 8996 34552 9002 34604
rect 9033 34595 9091 34601
rect 9033 34561 9045 34595
rect 9079 34561 9091 34595
rect 9033 34555 9091 34561
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2038 34524 2044 34536
rect 1443 34496 2044 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2498 34524 2504 34536
rect 2459 34496 2504 34524
rect 2498 34484 2504 34496
rect 2556 34484 2562 34536
rect 3421 34527 3479 34533
rect 3421 34493 3433 34527
rect 3467 34524 3479 34527
rect 3510 34524 3516 34536
rect 3467 34496 3516 34524
rect 3467 34493 3479 34496
rect 3421 34487 3479 34493
rect 3510 34484 3516 34496
rect 3568 34524 3574 34536
rect 4062 34524 4068 34536
rect 3568 34496 4068 34524
rect 3568 34484 3574 34496
rect 4062 34484 4068 34496
rect 4120 34484 4126 34536
rect 5905 34527 5963 34533
rect 5905 34493 5917 34527
rect 5951 34524 5963 34527
rect 6178 34524 6184 34536
rect 5951 34496 6184 34524
rect 5951 34493 5963 34496
rect 5905 34487 5963 34493
rect 6178 34484 6184 34496
rect 6236 34484 6242 34536
rect 7377 34527 7435 34533
rect 7377 34493 7389 34527
rect 7423 34524 7435 34527
rect 7929 34527 7987 34533
rect 7929 34524 7941 34527
rect 7423 34496 7941 34524
rect 7423 34493 7435 34496
rect 7377 34487 7435 34493
rect 7929 34493 7941 34496
rect 7975 34524 7987 34527
rect 8202 34524 8208 34536
rect 7975 34496 8208 34524
rect 7975 34493 7987 34496
rect 7929 34487 7987 34493
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 8389 34527 8447 34533
rect 8389 34493 8401 34527
rect 8435 34524 8447 34527
rect 8846 34524 8852 34536
rect 8435 34496 8708 34524
rect 8807 34496 8852 34524
rect 8435 34493 8447 34496
rect 8389 34487 8447 34493
rect 3694 34465 3700 34468
rect 3688 34456 3700 34465
rect 3655 34428 3700 34456
rect 3688 34419 3700 34428
rect 3694 34416 3700 34419
rect 3752 34416 3758 34468
rect 8680 34456 8708 34496
rect 8846 34484 8852 34496
rect 8904 34484 8910 34536
rect 9048 34524 9076 34555
rect 9122 34552 9128 34604
rect 9180 34592 9186 34604
rect 10689 34595 10747 34601
rect 10689 34592 10701 34595
rect 9180 34564 10701 34592
rect 9180 34552 9186 34564
rect 10689 34561 10701 34564
rect 10735 34592 10747 34595
rect 11422 34592 11428 34604
rect 10735 34564 11428 34592
rect 10735 34561 10747 34564
rect 10689 34555 10747 34561
rect 11422 34552 11428 34564
rect 11480 34552 11486 34604
rect 9861 34527 9919 34533
rect 8956 34496 9628 34524
rect 8956 34456 8984 34496
rect 8680 34428 8984 34456
rect 9600 34456 9628 34496
rect 9861 34493 9873 34527
rect 9907 34524 9919 34527
rect 10134 34524 10140 34536
rect 9907 34496 10140 34524
rect 9907 34493 9919 34496
rect 9861 34487 9919 34493
rect 10134 34484 10140 34496
rect 10192 34484 10198 34536
rect 10410 34524 10416 34536
rect 10371 34496 10416 34524
rect 10410 34484 10416 34496
rect 10468 34484 10474 34536
rect 10502 34484 10508 34536
rect 10560 34524 10566 34536
rect 11793 34527 11851 34533
rect 11793 34524 11805 34527
rect 10560 34496 11805 34524
rect 10560 34484 10566 34496
rect 11793 34493 11805 34496
rect 11839 34493 11851 34527
rect 11793 34487 11851 34493
rect 9950 34456 9956 34468
rect 9600 34428 9956 34456
rect 9950 34416 9956 34428
rect 10008 34416 10014 34468
rect 4614 34348 4620 34400
rect 4672 34388 4678 34400
rect 4801 34391 4859 34397
rect 4801 34388 4813 34391
rect 4672 34360 4813 34388
rect 4672 34348 4678 34360
rect 4801 34357 4813 34360
rect 4847 34357 4859 34391
rect 4801 34351 4859 34357
rect 6914 34348 6920 34400
rect 6972 34388 6978 34400
rect 7101 34391 7159 34397
rect 7101 34388 7113 34391
rect 6972 34360 7113 34388
rect 6972 34348 6978 34360
rect 7101 34357 7113 34360
rect 7147 34388 7159 34391
rect 7650 34388 7656 34400
rect 7147 34360 7656 34388
rect 7147 34357 7159 34360
rect 7101 34351 7159 34357
rect 7650 34348 7656 34360
rect 7708 34348 7714 34400
rect 11422 34388 11428 34400
rect 11383 34360 11428 34388
rect 11422 34348 11428 34360
rect 11480 34348 11486 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1762 34144 1768 34196
rect 1820 34184 1826 34196
rect 2869 34187 2927 34193
rect 2869 34184 2881 34187
rect 1820 34156 2881 34184
rect 1820 34144 1826 34156
rect 2869 34153 2881 34156
rect 2915 34153 2927 34187
rect 2869 34147 2927 34153
rect 5537 34187 5595 34193
rect 5537 34153 5549 34187
rect 5583 34153 5595 34187
rect 8938 34184 8944 34196
rect 8899 34156 8944 34184
rect 5537 34147 5595 34153
rect 1670 34116 1676 34128
rect 1631 34088 1676 34116
rect 1670 34076 1676 34088
rect 1728 34076 1734 34128
rect 4424 34119 4482 34125
rect 4424 34085 4436 34119
rect 4470 34116 4482 34119
rect 4614 34116 4620 34128
rect 4470 34088 4620 34116
rect 4470 34085 4482 34088
rect 4424 34079 4482 34085
rect 4614 34076 4620 34088
rect 4672 34076 4678 34128
rect 5552 34116 5580 34147
rect 8938 34144 8944 34156
rect 8996 34144 9002 34196
rect 11241 34187 11299 34193
rect 11241 34153 11253 34187
rect 11287 34184 11299 34187
rect 11422 34184 11428 34196
rect 11287 34156 11428 34184
rect 11287 34153 11299 34156
rect 11241 34147 11299 34153
rect 11422 34144 11428 34156
rect 11480 34144 11486 34196
rect 6730 34116 6736 34128
rect 5552 34088 6736 34116
rect 6730 34076 6736 34088
rect 6788 34116 6794 34128
rect 6886 34119 6944 34125
rect 6886 34116 6898 34119
rect 6788 34088 6898 34116
rect 6788 34076 6794 34088
rect 6886 34085 6898 34088
rect 6932 34085 6944 34119
rect 8662 34116 8668 34128
rect 8575 34088 8668 34116
rect 6886 34079 6944 34085
rect 8662 34076 8668 34088
rect 8720 34116 8726 34128
rect 9122 34116 9128 34128
rect 8720 34088 9128 34116
rect 8720 34076 8726 34088
rect 9122 34076 9128 34088
rect 9180 34076 9186 34128
rect 10134 34125 10140 34128
rect 10128 34116 10140 34125
rect 10047 34088 10140 34116
rect 10128 34079 10140 34088
rect 10192 34116 10198 34128
rect 10778 34116 10784 34128
rect 10192 34088 10784 34116
rect 10134 34076 10140 34079
rect 10192 34076 10198 34088
rect 10778 34076 10784 34088
rect 10836 34076 10842 34128
rect 1397 34051 1455 34057
rect 1397 34017 1409 34051
rect 1443 34048 1455 34051
rect 1486 34048 1492 34060
rect 1443 34020 1492 34048
rect 1443 34017 1455 34020
rect 1397 34011 1455 34017
rect 1486 34008 1492 34020
rect 1544 34008 1550 34060
rect 2685 34051 2743 34057
rect 2685 34017 2697 34051
rect 2731 34048 2743 34051
rect 2958 34048 2964 34060
rect 2731 34020 2964 34048
rect 2731 34017 2743 34020
rect 2685 34011 2743 34017
rect 2958 34008 2964 34020
rect 3016 34008 3022 34060
rect 4062 34008 4068 34060
rect 4120 34048 4126 34060
rect 4157 34051 4215 34057
rect 4157 34048 4169 34051
rect 4120 34020 4169 34048
rect 4120 34008 4126 34020
rect 4157 34017 4169 34020
rect 4203 34048 4215 34051
rect 5810 34048 5816 34060
rect 4203 34020 5816 34048
rect 4203 34017 4215 34020
rect 4157 34011 4215 34017
rect 5810 34008 5816 34020
rect 5868 34008 5874 34060
rect 6641 33983 6699 33989
rect 6641 33980 6653 33983
rect 6472 33952 6653 33980
rect 3694 33872 3700 33924
rect 3752 33872 3758 33924
rect 3513 33847 3571 33853
rect 3513 33813 3525 33847
rect 3559 33844 3571 33847
rect 3712 33844 3740 33872
rect 4338 33844 4344 33856
rect 3559 33816 4344 33844
rect 3559 33813 3571 33816
rect 3513 33807 3571 33813
rect 4338 33804 4344 33816
rect 4396 33804 4402 33856
rect 5810 33804 5816 33856
rect 5868 33844 5874 33856
rect 6472 33853 6500 33952
rect 6641 33949 6653 33952
rect 6687 33949 6699 33983
rect 6641 33943 6699 33949
rect 9306 33940 9312 33992
rect 9364 33980 9370 33992
rect 9861 33983 9919 33989
rect 9861 33980 9873 33983
rect 9364 33952 9873 33980
rect 9364 33940 9370 33952
rect 9861 33949 9873 33952
rect 9907 33949 9919 33983
rect 9861 33943 9919 33949
rect 6457 33847 6515 33853
rect 6457 33844 6469 33847
rect 5868 33816 6469 33844
rect 5868 33804 5874 33816
rect 6457 33813 6469 33816
rect 6503 33813 6515 33847
rect 8018 33844 8024 33856
rect 7979 33816 8024 33844
rect 6457 33807 6515 33813
rect 8018 33804 8024 33816
rect 8076 33804 8082 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1394 33600 1400 33652
rect 1452 33640 1458 33652
rect 1949 33643 2007 33649
rect 1949 33640 1961 33643
rect 1452 33612 1961 33640
rect 1452 33600 1458 33612
rect 1949 33609 1961 33612
rect 1995 33609 2007 33643
rect 1949 33603 2007 33609
rect 5629 33643 5687 33649
rect 5629 33609 5641 33643
rect 5675 33640 5687 33643
rect 5718 33640 5724 33652
rect 5675 33612 5724 33640
rect 5675 33609 5687 33612
rect 5629 33603 5687 33609
rect 5718 33600 5724 33612
rect 5776 33600 5782 33652
rect 8662 33640 8668 33652
rect 8623 33612 8668 33640
rect 8662 33600 8668 33612
rect 8720 33600 8726 33652
rect 9766 33600 9772 33652
rect 9824 33640 9830 33652
rect 9950 33640 9956 33652
rect 9824 33612 9956 33640
rect 9824 33600 9830 33612
rect 9950 33600 9956 33612
rect 10008 33640 10014 33652
rect 10229 33643 10287 33649
rect 10229 33640 10241 33643
rect 10008 33612 10241 33640
rect 10008 33600 10014 33612
rect 10229 33609 10241 33612
rect 10275 33609 10287 33643
rect 10229 33603 10287 33609
rect 1486 33532 1492 33584
rect 1544 33572 1550 33584
rect 1581 33575 1639 33581
rect 1581 33572 1593 33575
rect 1544 33544 1593 33572
rect 1544 33532 1550 33544
rect 1581 33541 1593 33544
rect 1627 33541 1639 33575
rect 1581 33535 1639 33541
rect 7653 33575 7711 33581
rect 7653 33541 7665 33575
rect 7699 33572 7711 33575
rect 7929 33575 7987 33581
rect 7929 33572 7941 33575
rect 7699 33544 7941 33572
rect 7699 33541 7711 33544
rect 7653 33535 7711 33541
rect 7929 33541 7941 33544
rect 7975 33572 7987 33575
rect 8570 33572 8576 33584
rect 7975 33544 8576 33572
rect 7975 33541 7987 33544
rect 7929 33535 7987 33541
rect 8570 33532 8576 33544
rect 8628 33532 8634 33584
rect 2406 33504 2412 33516
rect 1780 33476 2412 33504
rect 1780 33445 1808 33476
rect 2406 33464 2412 33476
rect 2464 33464 2470 33516
rect 6730 33464 6736 33516
rect 6788 33504 6794 33516
rect 7377 33507 7435 33513
rect 7377 33504 7389 33507
rect 6788 33476 7389 33504
rect 6788 33464 6794 33476
rect 7377 33473 7389 33476
rect 7423 33504 7435 33507
rect 8205 33507 8263 33513
rect 8205 33504 8217 33507
rect 7423 33476 8217 33504
rect 7423 33473 7435 33476
rect 7377 33467 7435 33473
rect 8205 33473 8217 33476
rect 8251 33473 8263 33507
rect 8680 33504 8708 33600
rect 8680 33476 8984 33504
rect 8205 33467 8263 33473
rect 1765 33439 1823 33445
rect 1765 33405 1777 33439
rect 1811 33405 1823 33439
rect 1765 33399 1823 33405
rect 2961 33439 3019 33445
rect 2961 33405 2973 33439
rect 3007 33436 3019 33439
rect 4062 33436 4068 33448
rect 3007 33408 4068 33436
rect 3007 33405 3019 33408
rect 2961 33399 3019 33405
rect 4062 33396 4068 33408
rect 4120 33396 4126 33448
rect 4798 33396 4804 33448
rect 4856 33436 4862 33448
rect 5445 33439 5503 33445
rect 5445 33436 5457 33439
rect 4856 33408 5457 33436
rect 4856 33396 4862 33408
rect 5445 33405 5457 33408
rect 5491 33436 5503 33439
rect 5997 33439 6055 33445
rect 5997 33436 6009 33439
rect 5491 33408 6009 33436
rect 5491 33405 5503 33408
rect 5445 33399 5503 33405
rect 5997 33405 6009 33408
rect 6043 33405 6055 33439
rect 5997 33399 6055 33405
rect 7193 33439 7251 33445
rect 7193 33405 7205 33439
rect 7239 33436 7251 33439
rect 7653 33439 7711 33445
rect 7653 33436 7665 33439
rect 7239 33408 7665 33436
rect 7239 33405 7251 33408
rect 7193 33399 7251 33405
rect 7653 33405 7665 33408
rect 7699 33405 7711 33439
rect 7653 33399 7711 33405
rect 8849 33439 8907 33445
rect 8849 33405 8861 33439
rect 8895 33405 8907 33439
rect 8956 33436 8984 33476
rect 11054 33464 11060 33516
rect 11112 33504 11118 33516
rect 11333 33507 11391 33513
rect 11333 33504 11345 33507
rect 11112 33476 11345 33504
rect 11112 33464 11118 33476
rect 11333 33473 11345 33476
rect 11379 33473 11391 33507
rect 11333 33467 11391 33473
rect 9105 33439 9163 33445
rect 9105 33436 9117 33439
rect 8956 33408 9117 33436
rect 8849 33399 8907 33405
rect 9105 33405 9117 33408
rect 9151 33405 9163 33439
rect 9105 33399 9163 33405
rect 3050 33328 3056 33380
rect 3108 33368 3114 33380
rect 3206 33371 3264 33377
rect 3206 33368 3218 33371
rect 3108 33340 3218 33368
rect 3108 33328 3114 33340
rect 3206 33337 3218 33340
rect 3252 33337 3264 33371
rect 7285 33371 7343 33377
rect 7285 33368 7297 33371
rect 3206 33331 3264 33337
rect 6564 33340 7297 33368
rect 2777 33303 2835 33309
rect 2777 33269 2789 33303
rect 2823 33300 2835 33303
rect 2958 33300 2964 33312
rect 2823 33272 2964 33300
rect 2823 33269 2835 33272
rect 2777 33263 2835 33269
rect 2958 33260 2964 33272
rect 3016 33260 3022 33312
rect 4338 33300 4344 33312
rect 4299 33272 4344 33300
rect 4338 33260 4344 33272
rect 4396 33260 4402 33312
rect 4614 33260 4620 33312
rect 4672 33300 4678 33312
rect 4893 33303 4951 33309
rect 4893 33300 4905 33303
rect 4672 33272 4905 33300
rect 4672 33260 4678 33272
rect 4893 33269 4905 33272
rect 4939 33269 4951 33303
rect 4893 33263 4951 33269
rect 5353 33303 5411 33309
rect 5353 33269 5365 33303
rect 5399 33300 5411 33303
rect 5810 33300 5816 33312
rect 5399 33272 5816 33300
rect 5399 33269 5411 33272
rect 5353 33263 5411 33269
rect 5810 33260 5816 33272
rect 5868 33260 5874 33312
rect 6086 33260 6092 33312
rect 6144 33300 6150 33312
rect 6564 33309 6592 33340
rect 7285 33337 7297 33340
rect 7331 33368 7343 33371
rect 8202 33368 8208 33380
rect 7331 33340 8208 33368
rect 7331 33337 7343 33340
rect 7285 33331 7343 33337
rect 8202 33328 8208 33340
rect 8260 33328 8266 33380
rect 8864 33368 8892 33399
rect 9306 33368 9312 33380
rect 8864 33340 9312 33368
rect 9306 33328 9312 33340
rect 9364 33368 9370 33380
rect 10781 33371 10839 33377
rect 10781 33368 10793 33371
rect 9364 33340 10793 33368
rect 9364 33328 9370 33340
rect 10781 33337 10793 33340
rect 10827 33337 10839 33371
rect 10781 33331 10839 33337
rect 6549 33303 6607 33309
rect 6549 33300 6561 33303
rect 6144 33272 6561 33300
rect 6144 33260 6150 33272
rect 6549 33269 6561 33272
rect 6595 33269 6607 33303
rect 6549 33263 6607 33269
rect 6638 33260 6644 33312
rect 6696 33300 6702 33312
rect 6825 33303 6883 33309
rect 6825 33300 6837 33303
rect 6696 33272 6837 33300
rect 6696 33260 6702 33272
rect 6825 33269 6837 33272
rect 6871 33269 6883 33303
rect 6825 33263 6883 33269
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 3789 33099 3847 33105
rect 3789 33065 3801 33099
rect 3835 33096 3847 33099
rect 4062 33096 4068 33108
rect 3835 33068 4068 33096
rect 3835 33065 3847 33068
rect 3789 33059 3847 33065
rect 4062 33056 4068 33068
rect 4120 33056 4126 33108
rect 4801 33099 4859 33105
rect 4801 33065 4813 33099
rect 4847 33096 4859 33099
rect 4982 33096 4988 33108
rect 4847 33068 4988 33096
rect 4847 33065 4859 33068
rect 4801 33059 4859 33065
rect 4982 33056 4988 33068
rect 5040 33056 5046 33108
rect 6730 33096 6736 33108
rect 6691 33068 6736 33096
rect 6730 33056 6736 33068
rect 6788 33056 6794 33108
rect 7282 33096 7288 33108
rect 7243 33068 7288 33096
rect 7282 33056 7288 33068
rect 7340 33056 7346 33108
rect 10137 33099 10195 33105
rect 10137 33065 10149 33099
rect 10183 33096 10195 33099
rect 10502 33096 10508 33108
rect 10183 33068 10508 33096
rect 10183 33065 10195 33068
rect 10137 33059 10195 33065
rect 10502 33056 10508 33068
rect 10560 33056 10566 33108
rect 10597 33031 10655 33037
rect 10597 32997 10609 33031
rect 10643 33028 10655 33031
rect 10778 33028 10784 33040
rect 10643 33000 10784 33028
rect 10643 32997 10655 33000
rect 10597 32991 10655 32997
rect 10778 32988 10784 33000
rect 10836 32988 10842 33040
rect 4430 32920 4436 32972
rect 4488 32960 4494 32972
rect 4617 32963 4675 32969
rect 4617 32960 4629 32963
rect 4488 32932 4629 32960
rect 4488 32920 4494 32932
rect 4617 32929 4629 32932
rect 4663 32929 4675 32963
rect 4617 32923 4675 32929
rect 8941 32963 8999 32969
rect 8941 32929 8953 32963
rect 8987 32960 8999 32963
rect 9490 32960 9496 32972
rect 8987 32932 9496 32960
rect 8987 32929 8999 32932
rect 8941 32923 8999 32929
rect 9490 32920 9496 32932
rect 9548 32960 9554 32972
rect 9953 32963 10011 32969
rect 9953 32960 9965 32963
rect 9548 32932 9965 32960
rect 9548 32920 9554 32932
rect 9953 32929 9965 32932
rect 9999 32960 10011 32963
rect 10134 32960 10140 32972
rect 9999 32932 10140 32960
rect 9999 32929 10011 32932
rect 9953 32923 10011 32929
rect 10134 32920 10140 32932
rect 10192 32920 10198 32972
rect 10226 32920 10232 32972
rect 10284 32960 10290 32972
rect 10505 32963 10563 32969
rect 10505 32960 10517 32963
rect 10284 32932 10517 32960
rect 10284 32920 10290 32932
rect 10505 32929 10517 32932
rect 10551 32929 10563 32963
rect 10505 32923 10563 32929
rect 6638 32852 6644 32904
rect 6696 32892 6702 32904
rect 7377 32895 7435 32901
rect 7377 32892 7389 32895
rect 6696 32864 7389 32892
rect 6696 32852 6702 32864
rect 7377 32861 7389 32864
rect 7423 32861 7435 32895
rect 7377 32855 7435 32861
rect 7561 32895 7619 32901
rect 7561 32861 7573 32895
rect 7607 32892 7619 32895
rect 8018 32892 8024 32904
rect 7607 32864 8024 32892
rect 7607 32861 7619 32864
rect 7561 32855 7619 32861
rect 6270 32784 6276 32836
rect 6328 32824 6334 32836
rect 7576 32824 7604 32855
rect 8018 32852 8024 32864
rect 8076 32852 8082 32904
rect 10152 32892 10180 32920
rect 10689 32895 10747 32901
rect 10689 32892 10701 32895
rect 10152 32864 10701 32892
rect 10689 32861 10701 32864
rect 10735 32892 10747 32895
rect 10870 32892 10876 32904
rect 10735 32864 10876 32892
rect 10735 32861 10747 32864
rect 10689 32855 10747 32861
rect 10870 32852 10876 32864
rect 10928 32852 10934 32904
rect 6328 32796 7604 32824
rect 6328 32784 6334 32796
rect 3050 32756 3056 32768
rect 3011 32728 3056 32756
rect 3050 32716 3056 32728
rect 3108 32716 3114 32768
rect 3418 32756 3424 32768
rect 3379 32728 3424 32756
rect 3418 32716 3424 32728
rect 3476 32716 3482 32768
rect 4522 32756 4528 32768
rect 4483 32728 4528 32756
rect 4522 32716 4528 32728
rect 4580 32716 4586 32768
rect 5258 32756 5264 32768
rect 5219 32728 5264 32756
rect 5258 32716 5264 32728
rect 5316 32716 5322 32768
rect 5350 32716 5356 32768
rect 5408 32756 5414 32768
rect 5537 32759 5595 32765
rect 5537 32756 5549 32759
rect 5408 32728 5549 32756
rect 5408 32716 5414 32728
rect 5537 32725 5549 32728
rect 5583 32725 5595 32759
rect 6914 32756 6920 32768
rect 6875 32728 6920 32756
rect 5537 32719 5595 32725
rect 6914 32716 6920 32728
rect 6972 32716 6978 32768
rect 9306 32756 9312 32768
rect 9267 32728 9312 32756
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 12526 32756 12532 32768
rect 12487 32728 12532 32756
rect 12526 32716 12532 32728
rect 12584 32716 12590 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 6270 32552 6276 32564
rect 6231 32524 6276 32552
rect 6270 32512 6276 32524
rect 6328 32512 6334 32564
rect 7101 32555 7159 32561
rect 7101 32521 7113 32555
rect 7147 32552 7159 32555
rect 7282 32552 7288 32564
rect 7147 32524 7288 32552
rect 7147 32521 7159 32524
rect 7101 32515 7159 32521
rect 7282 32512 7288 32524
rect 7340 32552 7346 32564
rect 7466 32552 7472 32564
rect 7340 32524 7472 32552
rect 7340 32512 7346 32524
rect 7466 32512 7472 32524
rect 7524 32512 7530 32564
rect 8386 32512 8392 32564
rect 8444 32552 8450 32564
rect 8849 32555 8907 32561
rect 8849 32552 8861 32555
rect 8444 32524 8861 32552
rect 8444 32512 8450 32524
rect 8849 32521 8861 32524
rect 8895 32521 8907 32555
rect 10870 32552 10876 32564
rect 10831 32524 10876 32552
rect 8849 32515 8907 32521
rect 10870 32512 10876 32524
rect 10928 32512 10934 32564
rect 3237 32487 3295 32493
rect 3237 32453 3249 32487
rect 3283 32484 3295 32487
rect 4338 32484 4344 32496
rect 3283 32456 4344 32484
rect 3283 32453 3295 32456
rect 3237 32447 3295 32453
rect 1578 32416 1584 32428
rect 1539 32388 1584 32416
rect 1578 32376 1584 32388
rect 1636 32376 1642 32428
rect 3418 32376 3424 32428
rect 3476 32416 3482 32428
rect 3988 32425 4016 32456
rect 4338 32444 4344 32456
rect 4396 32484 4402 32496
rect 5258 32484 5264 32496
rect 4396 32456 5264 32484
rect 4396 32444 4402 32456
rect 5258 32444 5264 32456
rect 5316 32484 5322 32496
rect 5316 32456 5488 32484
rect 5316 32444 5322 32456
rect 3789 32419 3847 32425
rect 3789 32416 3801 32419
rect 3476 32388 3801 32416
rect 3476 32376 3482 32388
rect 3789 32385 3801 32388
rect 3835 32385 3847 32419
rect 3789 32379 3847 32385
rect 3973 32419 4031 32425
rect 3973 32385 3985 32419
rect 4019 32385 4031 32419
rect 5350 32416 5356 32428
rect 5311 32388 5356 32416
rect 3973 32379 4031 32385
rect 5350 32376 5356 32388
rect 5408 32376 5414 32428
rect 5460 32425 5488 32456
rect 7558 32444 7564 32496
rect 7616 32484 7622 32496
rect 8665 32487 8723 32493
rect 8665 32484 8677 32487
rect 7616 32456 8677 32484
rect 7616 32444 7622 32456
rect 8665 32453 8677 32456
rect 8711 32453 8723 32487
rect 10226 32484 10232 32496
rect 10187 32456 10232 32484
rect 8665 32447 8723 32453
rect 5445 32419 5503 32425
rect 5445 32385 5457 32419
rect 5491 32385 5503 32419
rect 5445 32379 5503 32385
rect 5534 32376 5540 32428
rect 5592 32416 5598 32428
rect 6641 32419 6699 32425
rect 6641 32416 6653 32419
rect 5592 32388 6653 32416
rect 5592 32376 5598 32388
rect 6641 32385 6653 32388
rect 6687 32416 6699 32419
rect 7929 32419 7987 32425
rect 6687 32388 7696 32416
rect 6687 32385 6699 32388
rect 6641 32379 6699 32385
rect 1397 32351 1455 32357
rect 1397 32317 1409 32351
rect 1443 32317 1455 32351
rect 1397 32311 1455 32317
rect 1412 32212 1440 32311
rect 4522 32308 4528 32360
rect 4580 32348 4586 32360
rect 5261 32351 5319 32357
rect 5261 32348 5273 32351
rect 4580 32320 5273 32348
rect 4580 32308 4586 32320
rect 5261 32317 5273 32320
rect 5307 32348 5319 32351
rect 6822 32348 6828 32360
rect 5307 32320 6828 32348
rect 5307 32317 5319 32320
rect 5261 32311 5319 32317
rect 6822 32308 6828 32320
rect 6880 32308 6886 32360
rect 2869 32283 2927 32289
rect 2869 32249 2881 32283
rect 2915 32280 2927 32283
rect 3697 32283 3755 32289
rect 3697 32280 3709 32283
rect 2915 32252 3709 32280
rect 2915 32249 2927 32252
rect 2869 32243 2927 32249
rect 3697 32249 3709 32252
rect 3743 32280 3755 32283
rect 4154 32280 4160 32292
rect 3743 32252 4160 32280
rect 3743 32249 3755 32252
rect 3697 32243 3755 32249
rect 4154 32240 4160 32252
rect 4212 32240 4218 32292
rect 2222 32212 2228 32224
rect 1412 32184 2228 32212
rect 2222 32172 2228 32184
rect 2280 32172 2286 32224
rect 3326 32212 3332 32224
rect 3287 32184 3332 32212
rect 3326 32172 3332 32184
rect 3384 32172 3390 32224
rect 4430 32172 4436 32224
rect 4488 32212 4494 32224
rect 4617 32215 4675 32221
rect 4617 32212 4629 32215
rect 4488 32184 4629 32212
rect 4488 32172 4494 32184
rect 4617 32181 4629 32184
rect 4663 32181 4675 32215
rect 4890 32212 4896 32224
rect 4851 32184 4896 32212
rect 4617 32175 4675 32181
rect 4890 32172 4896 32184
rect 4948 32172 4954 32224
rect 7282 32212 7288 32224
rect 7243 32184 7288 32212
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 7668 32221 7696 32388
rect 7929 32385 7941 32419
rect 7975 32416 7987 32419
rect 8018 32416 8024 32428
rect 7975 32388 8024 32416
rect 7975 32385 7987 32388
rect 7929 32379 7987 32385
rect 8018 32376 8024 32388
rect 8076 32376 8082 32428
rect 8680 32348 8708 32447
rect 10226 32444 10232 32456
rect 10284 32444 10290 32496
rect 10597 32487 10655 32493
rect 10597 32453 10609 32487
rect 10643 32484 10655 32487
rect 10778 32484 10784 32496
rect 10643 32456 10784 32484
rect 10643 32453 10655 32456
rect 10597 32447 10655 32453
rect 9490 32416 9496 32428
rect 9451 32388 9496 32416
rect 9490 32376 9496 32388
rect 9548 32376 9554 32428
rect 10134 32376 10140 32428
rect 10192 32416 10198 32428
rect 10612 32416 10640 32447
rect 10778 32444 10784 32456
rect 10836 32444 10842 32496
rect 10192 32388 10640 32416
rect 10192 32376 10198 32388
rect 12526 32376 12532 32428
rect 12584 32416 12590 32428
rect 12894 32416 12900 32428
rect 12584 32388 12900 32416
rect 12584 32376 12590 32388
rect 12894 32376 12900 32388
rect 12952 32376 12958 32428
rect 13078 32416 13084 32428
rect 13039 32388 13084 32416
rect 13078 32376 13084 32388
rect 13136 32376 13142 32428
rect 9217 32351 9275 32357
rect 9217 32348 9229 32351
rect 8680 32320 9229 32348
rect 9217 32317 9229 32320
rect 9263 32317 9275 32351
rect 9217 32311 9275 32317
rect 12158 32308 12164 32360
rect 12216 32348 12222 32360
rect 12253 32351 12311 32357
rect 12253 32348 12265 32351
rect 12216 32320 12265 32348
rect 12216 32308 12222 32320
rect 12253 32317 12265 32320
rect 12299 32348 12311 32351
rect 13096 32348 13124 32376
rect 12299 32320 13124 32348
rect 12299 32317 12311 32320
rect 12253 32311 12311 32317
rect 7745 32283 7803 32289
rect 7745 32249 7757 32283
rect 7791 32280 7803 32283
rect 7834 32280 7840 32292
rect 7791 32252 7840 32280
rect 7791 32249 7803 32252
rect 7745 32243 7803 32249
rect 7834 32240 7840 32252
rect 7892 32280 7898 32292
rect 8389 32283 8447 32289
rect 8389 32280 8401 32283
rect 7892 32252 8401 32280
rect 7892 32240 7898 32252
rect 8389 32249 8401 32252
rect 8435 32280 8447 32283
rect 9398 32280 9404 32292
rect 8435 32252 9404 32280
rect 8435 32249 8447 32252
rect 8389 32243 8447 32249
rect 9398 32240 9404 32252
rect 9456 32240 9462 32292
rect 11885 32283 11943 32289
rect 11885 32249 11897 32283
rect 11931 32280 11943 32283
rect 12526 32280 12532 32292
rect 11931 32252 12532 32280
rect 11931 32249 11943 32252
rect 11885 32243 11943 32249
rect 12526 32240 12532 32252
rect 12584 32280 12590 32292
rect 12805 32283 12863 32289
rect 12805 32280 12817 32283
rect 12584 32252 12817 32280
rect 12584 32240 12590 32252
rect 12805 32249 12817 32252
rect 12851 32249 12863 32283
rect 12805 32243 12863 32249
rect 7653 32215 7711 32221
rect 7653 32181 7665 32215
rect 7699 32212 7711 32215
rect 8662 32212 8668 32224
rect 7699 32184 8668 32212
rect 7699 32181 7711 32184
rect 7653 32175 7711 32181
rect 8662 32172 8668 32184
rect 8720 32172 8726 32224
rect 8846 32172 8852 32224
rect 8904 32212 8910 32224
rect 9309 32215 9367 32221
rect 9309 32212 9321 32215
rect 8904 32184 9321 32212
rect 8904 32172 8910 32184
rect 9309 32181 9321 32184
rect 9355 32181 9367 32215
rect 9309 32175 9367 32181
rect 12434 32172 12440 32224
rect 12492 32212 12498 32224
rect 12492 32184 12537 32212
rect 12492 32172 12498 32184
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 2774 31968 2780 32020
rect 2832 32008 2838 32020
rect 2869 32011 2927 32017
rect 2869 32008 2881 32011
rect 2832 31980 2881 32008
rect 2832 31968 2838 31980
rect 2869 31977 2881 31980
rect 2915 32008 2927 32011
rect 3326 32008 3332 32020
rect 2915 31980 3332 32008
rect 2915 31977 2927 31980
rect 2869 31971 2927 31977
rect 3326 31968 3332 31980
rect 3384 31968 3390 32020
rect 5261 32011 5319 32017
rect 5261 31977 5273 32011
rect 5307 32008 5319 32011
rect 5350 32008 5356 32020
rect 5307 31980 5356 32008
rect 5307 31977 5319 31980
rect 5261 31971 5319 31977
rect 5350 31968 5356 31980
rect 5408 31968 5414 32020
rect 6365 32011 6423 32017
rect 6365 31977 6377 32011
rect 6411 32008 6423 32011
rect 6638 32008 6644 32020
rect 6411 31980 6644 32008
rect 6411 31977 6423 31980
rect 6365 31971 6423 31977
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 6822 32008 6828 32020
rect 6783 31980 6828 32008
rect 6822 31968 6828 31980
rect 6880 31968 6886 32020
rect 8570 31968 8576 32020
rect 8628 32008 8634 32020
rect 9398 32008 9404 32020
rect 8628 31980 9404 32008
rect 8628 31968 8634 31980
rect 9398 31968 9404 31980
rect 9456 31968 9462 32020
rect 10502 32008 10508 32020
rect 10463 31980 10508 32008
rect 10502 31968 10508 31980
rect 10560 31968 10566 32020
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 13449 32011 13507 32017
rect 13449 32008 13461 32011
rect 13136 31980 13461 32008
rect 13136 31968 13142 31980
rect 13449 31977 13461 31980
rect 13495 32008 13507 32011
rect 13814 32008 13820 32020
rect 13495 31980 13820 32008
rect 13495 31977 13507 31980
rect 13449 31971 13507 31977
rect 13814 31968 13820 31980
rect 13872 31968 13878 32020
rect 6730 31900 6736 31952
rect 6788 31940 6794 31952
rect 7285 31943 7343 31949
rect 7285 31940 7297 31943
rect 6788 31912 7297 31940
rect 6788 31900 6794 31912
rect 7285 31909 7297 31912
rect 7331 31940 7343 31943
rect 8478 31940 8484 31952
rect 7331 31912 8484 31940
rect 7331 31909 7343 31912
rect 7285 31903 7343 31909
rect 8478 31900 8484 31912
rect 8536 31900 8542 31952
rect 8846 31940 8852 31952
rect 8807 31912 8852 31940
rect 8846 31900 8852 31912
rect 8904 31900 8910 31952
rect 2777 31875 2835 31881
rect 2777 31841 2789 31875
rect 2823 31872 2835 31875
rect 2866 31872 2872 31884
rect 2823 31844 2872 31872
rect 2823 31841 2835 31844
rect 2777 31835 2835 31841
rect 2866 31832 2872 31844
rect 2924 31872 2930 31884
rect 4890 31872 4896 31884
rect 2924 31844 4896 31872
rect 2924 31832 2930 31844
rect 4890 31832 4896 31844
rect 4948 31832 4954 31884
rect 5629 31875 5687 31881
rect 5629 31841 5641 31875
rect 5675 31872 5687 31875
rect 6178 31872 6184 31884
rect 5675 31844 6184 31872
rect 5675 31841 5687 31844
rect 5629 31835 5687 31841
rect 6178 31832 6184 31844
rect 6236 31832 6242 31884
rect 6546 31832 6552 31884
rect 6604 31872 6610 31884
rect 7193 31875 7251 31881
rect 7193 31872 7205 31875
rect 6604 31844 7205 31872
rect 6604 31832 6610 31844
rect 7193 31841 7205 31844
rect 7239 31841 7251 31875
rect 7193 31835 7251 31841
rect 8202 31832 8208 31884
rect 8260 31872 8266 31884
rect 9490 31872 9496 31884
rect 8260 31844 9496 31872
rect 8260 31832 8266 31844
rect 9490 31832 9496 31844
rect 9548 31832 9554 31884
rect 10413 31875 10471 31881
rect 10413 31841 10425 31875
rect 10459 31872 10471 31875
rect 10870 31872 10876 31884
rect 10459 31844 10876 31872
rect 10459 31841 10471 31844
rect 10413 31835 10471 31841
rect 10870 31832 10876 31844
rect 10928 31832 10934 31884
rect 12342 31881 12348 31884
rect 12336 31872 12348 31881
rect 12303 31844 12348 31872
rect 12336 31835 12348 31844
rect 12342 31832 12348 31835
rect 12400 31832 12406 31884
rect 2961 31807 3019 31813
rect 2961 31773 2973 31807
rect 3007 31804 3019 31807
rect 5718 31804 5724 31816
rect 3007 31776 3041 31804
rect 5679 31776 5724 31804
rect 3007 31773 3019 31776
rect 2961 31767 3019 31773
rect 2682 31696 2688 31748
rect 2740 31736 2746 31748
rect 2976 31736 3004 31767
rect 5718 31764 5724 31776
rect 5776 31764 5782 31816
rect 5905 31807 5963 31813
rect 5905 31773 5917 31807
rect 5951 31804 5963 31807
rect 5951 31776 5985 31804
rect 5951 31773 5963 31776
rect 5905 31767 5963 31773
rect 4614 31736 4620 31748
rect 2740 31708 4620 31736
rect 2740 31696 2746 31708
rect 4614 31696 4620 31708
rect 4672 31696 4678 31748
rect 4985 31739 5043 31745
rect 4985 31705 4997 31739
rect 5031 31736 5043 31739
rect 5534 31736 5540 31748
rect 5031 31708 5540 31736
rect 5031 31705 5043 31708
rect 4985 31699 5043 31705
rect 5534 31696 5540 31708
rect 5592 31736 5598 31748
rect 5920 31736 5948 31767
rect 6822 31764 6828 31816
rect 6880 31804 6886 31816
rect 7282 31804 7288 31816
rect 6880 31776 7288 31804
rect 6880 31764 6886 31776
rect 7282 31764 7288 31776
rect 7340 31764 7346 31816
rect 7469 31807 7527 31813
rect 7469 31773 7481 31807
rect 7515 31804 7527 31807
rect 7515 31776 7549 31804
rect 7515 31773 7527 31776
rect 7469 31767 7527 31773
rect 7484 31736 7512 31767
rect 10318 31764 10324 31816
rect 10376 31804 10382 31816
rect 10376 31776 10456 31804
rect 10376 31764 10382 31776
rect 8202 31736 8208 31748
rect 5592 31708 8208 31736
rect 5592 31696 5598 31708
rect 8202 31696 8208 31708
rect 8260 31696 8266 31748
rect 10428 31680 10456 31776
rect 10594 31764 10600 31816
rect 10652 31764 10658 31816
rect 10778 31764 10784 31816
rect 10836 31804 10842 31816
rect 10965 31807 11023 31813
rect 10965 31804 10977 31807
rect 10836 31776 10977 31804
rect 10836 31764 10842 31776
rect 10965 31773 10977 31776
rect 11011 31773 11023 31807
rect 10965 31767 11023 31773
rect 11057 31807 11115 31813
rect 11057 31773 11069 31807
rect 11103 31804 11115 31807
rect 11977 31807 12035 31813
rect 11103 31776 11137 31804
rect 11103 31773 11115 31776
rect 11057 31767 11115 31773
rect 11977 31773 11989 31807
rect 12023 31804 12035 31807
rect 12066 31804 12072 31816
rect 12023 31776 12072 31804
rect 12023 31773 12035 31776
rect 11977 31767 12035 31773
rect 10502 31696 10508 31748
rect 10560 31736 10566 31748
rect 10612 31736 10640 31764
rect 10560 31708 10640 31736
rect 11072 31736 11100 31767
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 11146 31736 11152 31748
rect 11072 31708 11152 31736
rect 10560 31696 10566 31708
rect 11146 31696 11152 31708
rect 11204 31696 11210 31748
rect 2406 31668 2412 31680
rect 2367 31640 2412 31668
rect 2406 31628 2412 31640
rect 2464 31628 2470 31680
rect 4522 31668 4528 31680
rect 4483 31640 4528 31668
rect 4522 31628 4528 31640
rect 4580 31628 4586 31680
rect 6733 31671 6791 31677
rect 6733 31637 6745 31671
rect 6779 31668 6791 31671
rect 7374 31668 7380 31680
rect 6779 31640 7380 31668
rect 6779 31637 6791 31640
rect 6733 31631 6791 31637
rect 7374 31628 7380 31640
rect 7432 31628 7438 31680
rect 7742 31628 7748 31680
rect 7800 31668 7806 31680
rect 7837 31671 7895 31677
rect 7837 31668 7849 31671
rect 7800 31640 7849 31668
rect 7800 31628 7806 31640
rect 7837 31637 7849 31640
rect 7883 31668 7895 31671
rect 8018 31668 8024 31680
rect 7883 31640 8024 31668
rect 7883 31637 7895 31640
rect 7837 31631 7895 31637
rect 8018 31628 8024 31640
rect 8076 31628 8082 31680
rect 8478 31668 8484 31680
rect 8439 31640 8484 31668
rect 8478 31628 8484 31640
rect 8536 31628 8542 31680
rect 9858 31628 9864 31680
rect 9916 31668 9922 31680
rect 10042 31668 10048 31680
rect 9916 31640 10048 31668
rect 9916 31628 9922 31640
rect 10042 31628 10048 31640
rect 10100 31628 10106 31680
rect 10410 31628 10416 31680
rect 10468 31628 10474 31680
rect 11514 31668 11520 31680
rect 11475 31640 11520 31668
rect 11514 31628 11520 31640
rect 11572 31628 11578 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 2501 31467 2559 31473
rect 2501 31433 2513 31467
rect 2547 31464 2559 31467
rect 2682 31464 2688 31476
rect 2547 31436 2688 31464
rect 2547 31433 2559 31436
rect 2501 31427 2559 31433
rect 2682 31424 2688 31436
rect 2740 31424 2746 31476
rect 3329 31467 3387 31473
rect 3329 31433 3341 31467
rect 3375 31464 3387 31467
rect 3418 31464 3424 31476
rect 3375 31436 3424 31464
rect 3375 31433 3387 31436
rect 3329 31427 3387 31433
rect 3418 31424 3424 31436
rect 3476 31424 3482 31476
rect 4154 31424 4160 31476
rect 4212 31464 4218 31476
rect 4893 31467 4951 31473
rect 4893 31464 4905 31467
rect 4212 31436 4905 31464
rect 4212 31424 4218 31436
rect 4893 31433 4905 31436
rect 4939 31433 4951 31467
rect 4893 31427 4951 31433
rect 6086 31424 6092 31476
rect 6144 31464 6150 31476
rect 6641 31467 6699 31473
rect 6641 31464 6653 31467
rect 6144 31436 6653 31464
rect 6144 31424 6150 31436
rect 6641 31433 6653 31436
rect 6687 31464 6699 31467
rect 6730 31464 6736 31476
rect 6687 31436 6736 31464
rect 6687 31433 6699 31436
rect 6641 31427 6699 31433
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 7098 31424 7104 31476
rect 7156 31464 7162 31476
rect 7742 31464 7748 31476
rect 7156 31436 7748 31464
rect 7156 31424 7162 31436
rect 7742 31424 7748 31436
rect 7800 31424 7806 31476
rect 8202 31464 8208 31476
rect 8163 31436 8208 31464
rect 8202 31424 8208 31436
rect 8260 31424 8266 31476
rect 8386 31464 8392 31476
rect 8347 31436 8392 31464
rect 8386 31424 8392 31436
rect 8444 31424 8450 31476
rect 9490 31424 9496 31476
rect 9548 31464 9554 31476
rect 9858 31464 9864 31476
rect 9548 31436 9864 31464
rect 9548 31424 9554 31436
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 12526 31464 12532 31476
rect 12487 31436 12532 31464
rect 12526 31424 12532 31436
rect 12584 31424 12590 31476
rect 5626 31356 5632 31408
rect 5684 31396 5690 31408
rect 6546 31396 6552 31408
rect 5684 31368 6552 31396
rect 5684 31356 5690 31368
rect 6546 31356 6552 31368
rect 6604 31396 6610 31408
rect 7837 31399 7895 31405
rect 7837 31396 7849 31399
rect 6604 31368 7849 31396
rect 6604 31356 6610 31368
rect 7837 31365 7849 31368
rect 7883 31365 7895 31399
rect 7837 31359 7895 31365
rect 1578 31328 1584 31340
rect 1539 31300 1584 31328
rect 1578 31288 1584 31300
rect 1636 31288 1642 31340
rect 3050 31288 3056 31340
rect 3108 31328 3114 31340
rect 3237 31331 3295 31337
rect 3237 31328 3249 31331
rect 3108 31300 3249 31328
rect 3108 31288 3114 31300
rect 3237 31297 3249 31300
rect 3283 31328 3295 31331
rect 3973 31331 4031 31337
rect 3973 31328 3985 31331
rect 3283 31300 3985 31328
rect 3283 31297 3295 31300
rect 3237 31291 3295 31297
rect 3973 31297 3985 31300
rect 4019 31328 4031 31331
rect 4433 31331 4491 31337
rect 4433 31328 4445 31331
rect 4019 31300 4445 31328
rect 4019 31297 4031 31300
rect 3973 31291 4031 31297
rect 4433 31297 4445 31300
rect 4479 31328 4491 31331
rect 5534 31328 5540 31340
rect 4479 31300 5540 31328
rect 4479 31297 4491 31300
rect 4433 31291 4491 31297
rect 5534 31288 5540 31300
rect 5592 31288 5598 31340
rect 7374 31328 7380 31340
rect 7335 31300 7380 31328
rect 7374 31288 7380 31300
rect 7432 31288 7438 31340
rect 8478 31288 8484 31340
rect 8536 31328 8542 31340
rect 8941 31331 8999 31337
rect 8941 31328 8953 31331
rect 8536 31300 8953 31328
rect 8536 31288 8542 31300
rect 8941 31297 8953 31300
rect 8987 31297 8999 31331
rect 8941 31291 8999 31297
rect 9861 31331 9919 31337
rect 9861 31297 9873 31331
rect 9907 31328 9919 31331
rect 10778 31328 10784 31340
rect 9907 31300 10784 31328
rect 9907 31297 9919 31300
rect 9861 31291 9919 31297
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 11425 31331 11483 31337
rect 11425 31297 11437 31331
rect 11471 31297 11483 31331
rect 11425 31291 11483 31297
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31328 12311 31331
rect 12437 31331 12495 31337
rect 12437 31328 12449 31331
rect 12299 31300 12449 31328
rect 12299 31297 12311 31300
rect 12253 31291 12311 31297
rect 12437 31297 12449 31300
rect 12483 31297 12495 31331
rect 12437 31291 12495 31297
rect 13081 31331 13139 31337
rect 13081 31297 13093 31331
rect 13127 31297 13139 31331
rect 13081 31291 13139 31297
rect 1397 31263 1455 31269
rect 1397 31229 1409 31263
rect 1443 31260 1455 31263
rect 1670 31260 1676 31272
rect 1443 31232 1676 31260
rect 1443 31229 1455 31232
rect 1397 31223 1455 31229
rect 1670 31220 1676 31232
rect 1728 31260 1734 31272
rect 2406 31260 2412 31272
rect 1728 31232 2412 31260
rect 1728 31220 1734 31232
rect 2406 31220 2412 31232
rect 2464 31220 2470 31272
rect 6822 31220 6828 31272
rect 6880 31260 6886 31272
rect 10597 31263 10655 31269
rect 6880 31232 6951 31260
rect 6880 31220 6886 31232
rect 2869 31195 2927 31201
rect 2869 31161 2881 31195
rect 2915 31192 2927 31195
rect 3697 31195 3755 31201
rect 3697 31192 3709 31195
rect 2915 31164 3709 31192
rect 2915 31161 2927 31164
rect 2869 31155 2927 31161
rect 3697 31161 3709 31164
rect 3743 31192 3755 31195
rect 3970 31192 3976 31204
rect 3743 31164 3976 31192
rect 3743 31161 3755 31164
rect 3697 31155 3755 31161
rect 3970 31152 3976 31164
rect 4028 31152 4034 31204
rect 4522 31152 4528 31204
rect 4580 31192 4586 31204
rect 5353 31195 5411 31201
rect 5353 31192 5365 31195
rect 4580 31164 5365 31192
rect 4580 31152 4586 31164
rect 5353 31161 5365 31164
rect 5399 31161 5411 31195
rect 5353 31155 5411 31161
rect 3786 31084 3792 31136
rect 3844 31124 3850 31136
rect 3844 31096 3889 31124
rect 3844 31084 3850 31096
rect 4430 31084 4436 31136
rect 4488 31124 4494 31136
rect 4801 31127 4859 31133
rect 4801 31124 4813 31127
rect 4488 31096 4813 31124
rect 4488 31084 4494 31096
rect 4801 31093 4813 31096
rect 4847 31124 4859 31127
rect 5074 31124 5080 31136
rect 4847 31096 5080 31124
rect 4847 31093 4859 31096
rect 4801 31087 4859 31093
rect 5074 31084 5080 31096
rect 5132 31124 5138 31136
rect 5261 31127 5319 31133
rect 5261 31124 5273 31127
rect 5132 31096 5273 31124
rect 5132 31084 5138 31096
rect 5261 31093 5273 31096
rect 5307 31093 5319 31127
rect 5261 31087 5319 31093
rect 5997 31127 6055 31133
rect 5997 31093 6009 31127
rect 6043 31124 6055 31127
rect 6178 31124 6184 31136
rect 6043 31096 6184 31124
rect 6043 31093 6055 31096
rect 5997 31087 6055 31093
rect 6178 31084 6184 31096
rect 6236 31084 6242 31136
rect 6822 31124 6828 31136
rect 6783 31096 6828 31124
rect 6822 31084 6828 31096
rect 6880 31084 6886 31136
rect 6923 31124 6951 31232
rect 10597 31229 10609 31263
rect 10643 31260 10655 31263
rect 10962 31260 10968 31272
rect 10643 31232 10968 31260
rect 10643 31229 10655 31232
rect 10597 31223 10655 31229
rect 10962 31220 10968 31232
rect 11020 31220 11026 31272
rect 11440 31260 11468 31291
rect 12342 31260 12348 31272
rect 11440 31232 12348 31260
rect 12342 31220 12348 31232
rect 12400 31260 12406 31272
rect 12802 31260 12808 31272
rect 12400 31232 12808 31260
rect 12400 31220 12406 31232
rect 12802 31220 12808 31232
rect 12860 31260 12866 31272
rect 13096 31260 13124 31291
rect 13541 31263 13599 31269
rect 13541 31260 13553 31263
rect 12860 31232 13553 31260
rect 12860 31220 12866 31232
rect 13541 31229 13553 31232
rect 13587 31229 13599 31263
rect 13541 31223 13599 31229
rect 8570 31152 8576 31204
rect 8628 31192 8634 31204
rect 8849 31195 8907 31201
rect 8849 31192 8861 31195
rect 8628 31164 8861 31192
rect 8628 31152 8634 31164
rect 8849 31161 8861 31164
rect 8895 31161 8907 31195
rect 8849 31155 8907 31161
rect 10229 31195 10287 31201
rect 10229 31161 10241 31195
rect 10275 31192 10287 31195
rect 10318 31192 10324 31204
rect 10275 31164 10324 31192
rect 10275 31161 10287 31164
rect 10229 31155 10287 31161
rect 10318 31152 10324 31164
rect 10376 31192 10382 31204
rect 11149 31195 11207 31201
rect 11149 31192 11161 31195
rect 10376 31164 11161 31192
rect 10376 31152 10382 31164
rect 11149 31161 11161 31164
rect 11195 31192 11207 31195
rect 11422 31192 11428 31204
rect 11195 31164 11428 31192
rect 11195 31161 11207 31164
rect 11149 31155 11207 31161
rect 11422 31152 11428 31164
rect 11480 31152 11486 31204
rect 11885 31195 11943 31201
rect 11885 31161 11897 31195
rect 11931 31192 11943 31195
rect 12897 31195 12955 31201
rect 12897 31192 12909 31195
rect 11931 31164 12909 31192
rect 11931 31161 11943 31164
rect 11885 31155 11943 31161
rect 12897 31161 12909 31164
rect 12943 31192 12955 31195
rect 13078 31192 13084 31204
rect 12943 31164 13084 31192
rect 12943 31161 12955 31164
rect 12897 31155 12955 31161
rect 13078 31152 13084 31164
rect 13136 31152 13142 31204
rect 7193 31127 7251 31133
rect 7193 31124 7205 31127
rect 6923 31096 7205 31124
rect 7193 31093 7205 31096
rect 7239 31093 7251 31127
rect 7193 31087 7251 31093
rect 7282 31084 7288 31136
rect 7340 31124 7346 31136
rect 8754 31124 8760 31136
rect 7340 31096 7385 31124
rect 8715 31096 8760 31124
rect 7340 31084 7346 31096
rect 8754 31084 8760 31096
rect 8812 31124 8818 31136
rect 9401 31127 9459 31133
rect 9401 31124 9413 31127
rect 8812 31096 9413 31124
rect 8812 31084 8818 31096
rect 9401 31093 9413 31096
rect 9447 31093 9459 31127
rect 9401 31087 9459 31093
rect 10781 31127 10839 31133
rect 10781 31093 10793 31127
rect 10827 31124 10839 31127
rect 11054 31124 11060 31136
rect 10827 31096 11060 31124
rect 10827 31093 10839 31096
rect 10781 31087 10839 31093
rect 11054 31084 11060 31096
rect 11112 31084 11118 31136
rect 11241 31127 11299 31133
rect 11241 31093 11253 31127
rect 11287 31124 11299 31127
rect 11514 31124 11520 31136
rect 11287 31096 11520 31124
rect 11287 31093 11299 31096
rect 11241 31087 11299 31093
rect 11514 31084 11520 31096
rect 11572 31124 11578 31136
rect 12342 31124 12348 31136
rect 11572 31096 12348 31124
rect 11572 31084 11578 31096
rect 12342 31084 12348 31096
rect 12400 31084 12406 31136
rect 12437 31127 12495 31133
rect 12437 31093 12449 31127
rect 12483 31124 12495 31127
rect 12989 31127 13047 31133
rect 12989 31124 13001 31127
rect 12483 31096 13001 31124
rect 12483 31093 12495 31096
rect 12437 31087 12495 31093
rect 12989 31093 13001 31096
rect 13035 31124 13047 31127
rect 13262 31124 13268 31136
rect 13035 31096 13268 31124
rect 13035 31093 13047 31096
rect 12989 31087 13047 31093
rect 13262 31084 13268 31096
rect 13320 31084 13326 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 1670 30920 1676 30932
rect 1631 30892 1676 30920
rect 1670 30880 1676 30892
rect 1728 30880 1734 30932
rect 2593 30923 2651 30929
rect 2593 30889 2605 30923
rect 2639 30920 2651 30923
rect 2682 30920 2688 30932
rect 2639 30892 2688 30920
rect 2639 30889 2651 30892
rect 2593 30883 2651 30889
rect 2682 30880 2688 30892
rect 2740 30880 2746 30932
rect 2866 30920 2872 30932
rect 2827 30892 2872 30920
rect 2866 30880 2872 30892
rect 2924 30880 2930 30932
rect 3421 30923 3479 30929
rect 3421 30889 3433 30923
rect 3467 30920 3479 30923
rect 3510 30920 3516 30932
rect 3467 30892 3516 30920
rect 3467 30889 3479 30892
rect 3421 30883 3479 30889
rect 3510 30880 3516 30892
rect 3568 30920 3574 30932
rect 3786 30920 3792 30932
rect 3568 30892 3792 30920
rect 3568 30880 3574 30892
rect 3786 30880 3792 30892
rect 3844 30880 3850 30932
rect 3970 30880 3976 30932
rect 4028 30920 4034 30932
rect 4065 30923 4123 30929
rect 4065 30920 4077 30923
rect 4028 30892 4077 30920
rect 4028 30880 4034 30892
rect 4065 30889 4077 30892
rect 4111 30889 4123 30923
rect 5350 30920 5356 30932
rect 5311 30892 5356 30920
rect 4065 30883 4123 30889
rect 5350 30880 5356 30892
rect 5408 30880 5414 30932
rect 5626 30920 5632 30932
rect 5587 30892 5632 30920
rect 5626 30880 5632 30892
rect 5684 30880 5690 30932
rect 6549 30923 6607 30929
rect 6549 30889 6561 30923
rect 6595 30920 6607 30923
rect 6914 30920 6920 30932
rect 6595 30892 6920 30920
rect 6595 30889 6607 30892
rect 6549 30883 6607 30889
rect 6914 30880 6920 30892
rect 6972 30920 6978 30932
rect 7282 30920 7288 30932
rect 6972 30892 7288 30920
rect 6972 30880 6978 30892
rect 7282 30880 7288 30892
rect 7340 30880 7346 30932
rect 8018 30920 8024 30932
rect 7931 30892 8024 30920
rect 8018 30880 8024 30892
rect 8076 30920 8082 30932
rect 8386 30920 8392 30932
rect 8076 30892 8392 30920
rect 8076 30880 8082 30892
rect 8386 30880 8392 30892
rect 8444 30880 8450 30932
rect 8570 30920 8576 30932
rect 8531 30892 8576 30920
rect 8570 30880 8576 30892
rect 8628 30880 8634 30932
rect 6181 30855 6239 30861
rect 6181 30821 6193 30855
rect 6227 30852 6239 30855
rect 6730 30852 6736 30864
rect 6227 30824 6736 30852
rect 6227 30821 6239 30824
rect 6181 30815 6239 30821
rect 6730 30812 6736 30824
rect 6788 30812 6794 30864
rect 12158 30812 12164 30864
rect 12216 30852 12222 30864
rect 12314 30855 12372 30861
rect 12314 30852 12326 30855
rect 12216 30824 12326 30852
rect 12216 30812 12222 30824
rect 12314 30821 12326 30824
rect 12360 30821 12372 30855
rect 12314 30815 12372 30821
rect 1949 30787 2007 30793
rect 1949 30753 1961 30787
rect 1995 30784 2007 30787
rect 2038 30784 2044 30796
rect 1995 30756 2044 30784
rect 1995 30753 2007 30756
rect 1949 30747 2007 30753
rect 2038 30744 2044 30756
rect 2096 30744 2102 30796
rect 4430 30784 4436 30796
rect 4391 30756 4436 30784
rect 4430 30744 4436 30756
rect 4488 30744 4494 30796
rect 4525 30787 4583 30793
rect 4525 30753 4537 30787
rect 4571 30784 4583 30787
rect 4982 30784 4988 30796
rect 4571 30756 4988 30784
rect 4571 30753 4583 30756
rect 4525 30747 4583 30753
rect 4982 30744 4988 30756
rect 5040 30744 5046 30796
rect 6914 30793 6920 30796
rect 6908 30784 6920 30793
rect 6875 30756 6920 30784
rect 6908 30747 6920 30756
rect 6972 30784 6978 30796
rect 7374 30784 7380 30796
rect 6972 30756 7380 30784
rect 6914 30744 6920 30747
rect 6972 30744 6978 30756
rect 7374 30744 7380 30756
rect 7432 30744 7438 30796
rect 10870 30784 10876 30796
rect 10831 30756 10876 30784
rect 10870 30744 10876 30756
rect 10928 30744 10934 30796
rect 12066 30784 12072 30796
rect 12027 30756 12072 30784
rect 12066 30744 12072 30756
rect 12124 30744 12130 30796
rect 4709 30719 4767 30725
rect 4709 30685 4721 30719
rect 4755 30716 4767 30719
rect 4798 30716 4804 30728
rect 4755 30688 4804 30716
rect 4755 30685 4767 30688
rect 4709 30679 4767 30685
rect 934 30608 940 30660
rect 992 30648 998 30660
rect 2133 30651 2191 30657
rect 2133 30648 2145 30651
rect 992 30620 2145 30648
rect 992 30608 998 30620
rect 2133 30617 2145 30620
rect 2179 30617 2191 30651
rect 2133 30611 2191 30617
rect 3881 30651 3939 30657
rect 3881 30617 3893 30651
rect 3927 30648 3939 30651
rect 4724 30648 4752 30679
rect 4798 30676 4804 30688
rect 4856 30676 4862 30728
rect 6546 30676 6552 30728
rect 6604 30716 6610 30728
rect 6641 30719 6699 30725
rect 6641 30716 6653 30719
rect 6604 30688 6653 30716
rect 6604 30676 6610 30688
rect 6641 30685 6653 30688
rect 6687 30685 6699 30719
rect 6641 30679 6699 30685
rect 10045 30719 10103 30725
rect 10045 30685 10057 30719
rect 10091 30716 10103 30719
rect 10594 30716 10600 30728
rect 10091 30688 10600 30716
rect 10091 30685 10103 30688
rect 10045 30679 10103 30685
rect 10594 30676 10600 30688
rect 10652 30716 10658 30728
rect 10965 30719 11023 30725
rect 10965 30716 10977 30719
rect 10652 30688 10977 30716
rect 10652 30676 10658 30688
rect 10965 30685 10977 30688
rect 11011 30685 11023 30719
rect 10965 30679 11023 30685
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30685 11115 30719
rect 11057 30679 11115 30685
rect 3927 30620 4752 30648
rect 10413 30651 10471 30657
rect 3927 30617 3939 30620
rect 3881 30611 3939 30617
rect 10413 30617 10425 30651
rect 10459 30648 10471 30651
rect 11072 30648 11100 30679
rect 11517 30651 11575 30657
rect 11517 30648 11529 30651
rect 10459 30620 11529 30648
rect 10459 30617 10471 30620
rect 10413 30611 10471 30617
rect 11517 30617 11529 30620
rect 11563 30648 11575 30651
rect 11885 30651 11943 30657
rect 11885 30648 11897 30651
rect 11563 30620 11897 30648
rect 11563 30617 11575 30620
rect 11517 30611 11575 30617
rect 11885 30617 11897 30620
rect 11931 30617 11943 30651
rect 11885 30611 11943 30617
rect 10505 30583 10563 30589
rect 10505 30549 10517 30583
rect 10551 30580 10563 30583
rect 10962 30580 10968 30592
rect 10551 30552 10968 30580
rect 10551 30549 10563 30552
rect 10505 30543 10563 30549
rect 10962 30540 10968 30552
rect 11020 30540 11026 30592
rect 11900 30580 11928 30611
rect 12802 30580 12808 30592
rect 11900 30552 12808 30580
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 13446 30580 13452 30592
rect 13407 30552 13452 30580
rect 13446 30540 13452 30552
rect 13504 30540 13510 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 3510 30336 3516 30388
rect 3568 30376 3574 30388
rect 3789 30379 3847 30385
rect 3789 30376 3801 30379
rect 3568 30348 3801 30376
rect 3568 30336 3574 30348
rect 3789 30345 3801 30348
rect 3835 30345 3847 30379
rect 3789 30339 3847 30345
rect 6178 30336 6184 30388
rect 6236 30376 6242 30388
rect 6730 30376 6736 30388
rect 6236 30348 6736 30376
rect 6236 30336 6242 30348
rect 6730 30336 6736 30348
rect 6788 30336 6794 30388
rect 10870 30376 10876 30388
rect 9600 30348 10876 30376
rect 9309 30311 9367 30317
rect 9309 30277 9321 30311
rect 9355 30308 9367 30311
rect 9600 30308 9628 30348
rect 10870 30336 10876 30348
rect 10928 30336 10934 30388
rect 12434 30336 12440 30388
rect 12492 30376 12498 30388
rect 12492 30348 12537 30376
rect 12492 30336 12498 30348
rect 9355 30280 9628 30308
rect 9355 30277 9367 30280
rect 9309 30271 9367 30277
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 9732 30280 9777 30308
rect 9732 30268 9738 30280
rect 11514 30268 11520 30320
rect 11572 30308 11578 30320
rect 11974 30308 11980 30320
rect 11572 30280 11980 30308
rect 11572 30268 11578 30280
rect 11974 30268 11980 30280
rect 12032 30308 12038 30320
rect 12161 30311 12219 30317
rect 12161 30308 12173 30311
rect 12032 30280 12173 30308
rect 12032 30268 12038 30280
rect 12161 30277 12173 30280
rect 12207 30277 12219 30311
rect 13814 30308 13820 30320
rect 13775 30280 13820 30308
rect 12161 30271 12219 30277
rect 3329 30243 3387 30249
rect 3329 30209 3341 30243
rect 3375 30240 3387 30243
rect 4433 30243 4491 30249
rect 4433 30240 4445 30243
rect 3375 30212 4445 30240
rect 3375 30209 3387 30212
rect 3329 30203 3387 30209
rect 4433 30209 4445 30212
rect 4479 30240 4491 30243
rect 4798 30240 4804 30252
rect 4479 30212 4804 30240
rect 4479 30209 4491 30212
rect 4433 30203 4491 30209
rect 4798 30200 4804 30212
rect 4856 30200 4862 30252
rect 5810 30240 5816 30252
rect 5368 30212 5816 30240
rect 2038 30172 2044 30184
rect 1999 30144 2044 30172
rect 2038 30132 2044 30144
rect 2096 30132 2102 30184
rect 4893 30175 4951 30181
rect 4893 30141 4905 30175
rect 4939 30172 4951 30175
rect 4982 30172 4988 30184
rect 4939 30144 4988 30172
rect 4939 30141 4951 30144
rect 4893 30135 4951 30141
rect 4982 30132 4988 30144
rect 5040 30132 5046 30184
rect 4249 30107 4307 30113
rect 4249 30104 4261 30107
rect 3620 30076 4261 30104
rect 2590 29996 2596 30048
rect 2648 30036 2654 30048
rect 3620 30045 3648 30076
rect 4249 30073 4261 30076
rect 4295 30104 4307 30107
rect 5258 30104 5264 30116
rect 4295 30076 5264 30104
rect 4295 30073 4307 30076
rect 4249 30067 4307 30073
rect 5258 30064 5264 30076
rect 5316 30064 5322 30116
rect 3605 30039 3663 30045
rect 3605 30036 3617 30039
rect 2648 30008 3617 30036
rect 2648 29996 2654 30008
rect 3605 30005 3617 30008
rect 3651 30005 3663 30039
rect 4154 30036 4160 30048
rect 4115 30008 4160 30036
rect 3605 29999 3663 30005
rect 4154 29996 4160 30008
rect 4212 29996 4218 30048
rect 4982 29996 4988 30048
rect 5040 30036 5046 30048
rect 5368 30045 5396 30212
rect 5810 30200 5816 30212
rect 5868 30240 5874 30252
rect 6181 30243 6239 30249
rect 6181 30240 6193 30243
rect 5868 30212 6193 30240
rect 5868 30200 5874 30212
rect 6181 30209 6193 30212
rect 6227 30240 6239 30243
rect 6546 30240 6552 30252
rect 6227 30212 6552 30240
rect 6227 30209 6239 30212
rect 6181 30203 6239 30209
rect 6546 30200 6552 30212
rect 6604 30200 6610 30252
rect 7193 30243 7251 30249
rect 7193 30209 7205 30243
rect 7239 30240 7251 30243
rect 12176 30240 12204 30271
rect 13814 30268 13820 30280
rect 13872 30268 13878 30320
rect 12897 30243 12955 30249
rect 12897 30240 12909 30243
rect 7239 30212 7420 30240
rect 12176 30212 12909 30240
rect 7239 30209 7251 30212
rect 7193 30203 7251 30209
rect 5537 30175 5595 30181
rect 5537 30141 5549 30175
rect 5583 30172 5595 30175
rect 7282 30172 7288 30184
rect 5583 30144 5764 30172
rect 7243 30144 7288 30172
rect 5583 30141 5595 30144
rect 5537 30135 5595 30141
rect 5736 30048 5764 30144
rect 7282 30132 7288 30144
rect 7340 30132 7346 30184
rect 7392 30172 7420 30212
rect 12897 30209 12909 30212
rect 12943 30209 12955 30243
rect 12897 30203 12955 30209
rect 13081 30243 13139 30249
rect 13081 30209 13093 30243
rect 13127 30240 13139 30243
rect 13446 30240 13452 30252
rect 13127 30212 13452 30240
rect 13127 30209 13139 30212
rect 13081 30203 13139 30209
rect 13446 30200 13452 30212
rect 13504 30200 13510 30252
rect 7552 30175 7610 30181
rect 7552 30172 7564 30175
rect 7392 30144 7564 30172
rect 7552 30141 7564 30144
rect 7598 30172 7610 30175
rect 8018 30172 8024 30184
rect 7598 30144 8024 30172
rect 7598 30141 7610 30144
rect 7552 30135 7610 30141
rect 8018 30132 8024 30144
rect 8076 30132 8082 30184
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 9674 30172 9680 30184
rect 9364 30144 9680 30172
rect 9364 30132 9370 30144
rect 9674 30132 9680 30144
rect 9732 30172 9738 30184
rect 9769 30175 9827 30181
rect 9769 30172 9781 30175
rect 9732 30144 9781 30172
rect 9732 30132 9738 30144
rect 9769 30141 9781 30144
rect 9815 30141 9827 30175
rect 9769 30135 9827 30141
rect 10036 30175 10094 30181
rect 10036 30141 10048 30175
rect 10082 30172 10094 30175
rect 10318 30172 10324 30184
rect 10082 30144 10324 30172
rect 10082 30141 10094 30144
rect 10036 30135 10094 30141
rect 10318 30132 10324 30144
rect 10376 30132 10382 30184
rect 12342 30132 12348 30184
rect 12400 30172 12406 30184
rect 12805 30175 12863 30181
rect 12805 30172 12817 30175
rect 12400 30144 12817 30172
rect 12400 30132 12406 30144
rect 12805 30141 12817 30144
rect 12851 30141 12863 30175
rect 12805 30135 12863 30141
rect 5353 30039 5411 30045
rect 5353 30036 5365 30039
rect 5040 30008 5365 30036
rect 5040 29996 5046 30008
rect 5353 30005 5365 30008
rect 5399 30005 5411 30039
rect 5353 29999 5411 30005
rect 5718 29996 5724 30048
rect 5776 30036 5782 30048
rect 5813 30039 5871 30045
rect 5813 30036 5825 30039
rect 5776 30008 5825 30036
rect 5776 29996 5782 30008
rect 5813 30005 5825 30008
rect 5859 30005 5871 30039
rect 6638 30036 6644 30048
rect 6599 30008 6644 30036
rect 5813 29999 5871 30005
rect 6638 29996 6644 30008
rect 6696 30036 6702 30048
rect 6914 30036 6920 30048
rect 6696 30008 6920 30036
rect 6696 29996 6702 30008
rect 6914 29996 6920 30008
rect 6972 29996 6978 30048
rect 8662 30036 8668 30048
rect 8623 30008 8668 30036
rect 8662 29996 8668 30008
rect 8720 29996 8726 30048
rect 11149 30039 11207 30045
rect 11149 30005 11161 30039
rect 11195 30036 11207 30039
rect 11238 30036 11244 30048
rect 11195 30008 11244 30036
rect 11195 30005 11207 30008
rect 11149 29999 11207 30005
rect 11238 29996 11244 30008
rect 11296 29996 11302 30048
rect 11885 30039 11943 30045
rect 11885 30005 11897 30039
rect 11931 30036 11943 30039
rect 12250 30036 12256 30048
rect 11931 30008 12256 30036
rect 11931 30005 11943 30008
rect 11885 29999 11943 30005
rect 12250 29996 12256 30008
rect 12308 29996 12314 30048
rect 13446 30036 13452 30048
rect 13407 30008 13452 30036
rect 13446 29996 13452 30008
rect 13504 29996 13510 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 4341 29835 4399 29841
rect 4341 29801 4353 29835
rect 4387 29832 4399 29835
rect 4430 29832 4436 29844
rect 4387 29804 4436 29832
rect 4387 29801 4399 29804
rect 4341 29795 4399 29801
rect 4430 29792 4436 29804
rect 4488 29792 4494 29844
rect 5534 29792 5540 29844
rect 5592 29832 5598 29844
rect 6089 29835 6147 29841
rect 6089 29832 6101 29835
rect 5592 29804 6101 29832
rect 5592 29792 5598 29804
rect 6089 29801 6101 29804
rect 6135 29801 6147 29835
rect 6089 29795 6147 29801
rect 7926 29792 7932 29844
rect 7984 29832 7990 29844
rect 8021 29835 8079 29841
rect 8021 29832 8033 29835
rect 7984 29804 8033 29832
rect 7984 29792 7990 29804
rect 8021 29801 8033 29804
rect 8067 29801 8079 29835
rect 8021 29795 8079 29801
rect 9493 29835 9551 29841
rect 9493 29801 9505 29835
rect 9539 29832 9551 29835
rect 9539 29804 9720 29832
rect 9539 29801 9551 29804
rect 9493 29795 9551 29801
rect 3881 29767 3939 29773
rect 3881 29733 3893 29767
rect 3927 29764 3939 29767
rect 4154 29764 4160 29776
rect 3927 29736 4160 29764
rect 3927 29733 3939 29736
rect 3881 29727 3939 29733
rect 4154 29724 4160 29736
rect 4212 29764 4218 29776
rect 4212 29736 5120 29764
rect 4212 29724 4218 29736
rect 4798 29656 4804 29708
rect 4856 29696 4862 29708
rect 4965 29699 5023 29705
rect 4965 29696 4977 29699
rect 4856 29668 4977 29696
rect 4856 29656 4862 29668
rect 4965 29665 4977 29668
rect 5011 29665 5023 29699
rect 5092 29696 5120 29736
rect 7282 29724 7288 29776
rect 7340 29764 7346 29776
rect 7377 29767 7435 29773
rect 7377 29764 7389 29767
rect 7340 29736 7389 29764
rect 7340 29724 7346 29736
rect 7377 29733 7389 29736
rect 7423 29764 7435 29767
rect 9692 29764 9720 29804
rect 10870 29792 10876 29844
rect 10928 29832 10934 29844
rect 12161 29835 12219 29841
rect 12161 29832 12173 29835
rect 10928 29804 12173 29832
rect 10928 29792 10934 29804
rect 12161 29801 12173 29804
rect 12207 29801 12219 29835
rect 12161 29795 12219 29801
rect 9766 29764 9772 29776
rect 7423 29736 9772 29764
rect 7423 29733 7435 29736
rect 7377 29727 7435 29733
rect 8110 29696 8116 29708
rect 5092 29668 8116 29696
rect 4965 29659 5023 29665
rect 8110 29656 8116 29668
rect 8168 29656 8174 29708
rect 8386 29696 8392 29708
rect 8347 29668 8392 29696
rect 8386 29656 8392 29668
rect 8444 29656 8450 29708
rect 4709 29631 4767 29637
rect 4709 29597 4721 29631
rect 4755 29597 4767 29631
rect 4709 29591 4767 29597
rect 7929 29631 7987 29637
rect 7929 29597 7941 29631
rect 7975 29628 7987 29631
rect 8478 29628 8484 29640
rect 7975 29600 8484 29628
rect 7975 29597 7987 29600
rect 7929 29591 7987 29597
rect 4724 29492 4752 29591
rect 8478 29588 8484 29600
rect 8536 29588 8542 29640
rect 8570 29588 8576 29640
rect 8628 29628 8634 29640
rect 9692 29637 9720 29736
rect 9766 29724 9772 29736
rect 9824 29764 9830 29776
rect 11146 29764 11152 29776
rect 9824 29736 11152 29764
rect 9824 29724 9830 29736
rect 11146 29724 11152 29736
rect 11204 29764 11210 29776
rect 12066 29764 12072 29776
rect 11204 29736 12072 29764
rect 11204 29724 11210 29736
rect 12066 29724 12072 29736
rect 12124 29724 12130 29776
rect 12250 29724 12256 29776
rect 12308 29764 12314 29776
rect 12621 29767 12679 29773
rect 12621 29764 12633 29767
rect 12308 29736 12633 29764
rect 12308 29724 12314 29736
rect 12621 29733 12633 29736
rect 12667 29733 12679 29767
rect 12621 29727 12679 29733
rect 9944 29699 10002 29705
rect 9944 29665 9956 29699
rect 9990 29696 10002 29699
rect 10318 29696 10324 29708
rect 9990 29668 10324 29696
rect 9990 29665 10002 29668
rect 9944 29659 10002 29665
rect 10318 29656 10324 29668
rect 10376 29656 10382 29708
rect 12526 29696 12532 29708
rect 12487 29668 12532 29696
rect 12526 29656 12532 29668
rect 12584 29656 12590 29708
rect 9677 29631 9735 29637
rect 8628 29600 8673 29628
rect 8628 29588 8634 29600
rect 9677 29597 9689 29631
rect 9723 29597 9735 29631
rect 9677 29591 9735 29597
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29628 12863 29631
rect 13446 29628 13452 29640
rect 12851 29600 13452 29628
rect 12851 29597 12863 29600
rect 12805 29591 12863 29597
rect 11057 29563 11115 29569
rect 11057 29529 11069 29563
rect 11103 29560 11115 29563
rect 11146 29560 11152 29572
rect 11103 29532 11152 29560
rect 11103 29529 11115 29532
rect 11057 29523 11115 29529
rect 11146 29520 11152 29532
rect 11204 29520 11210 29572
rect 11238 29520 11244 29572
rect 11296 29560 11302 29572
rect 12820 29560 12848 29591
rect 13446 29588 13452 29600
rect 13504 29588 13510 29640
rect 11296 29532 12848 29560
rect 11296 29520 11302 29532
rect 4982 29492 4988 29504
rect 4724 29464 4988 29492
rect 4982 29452 4988 29464
rect 5040 29452 5046 29504
rect 6914 29492 6920 29504
rect 6875 29464 6920 29492
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 12802 29452 12808 29504
rect 12860 29492 12866 29504
rect 13173 29495 13231 29501
rect 13173 29492 13185 29495
rect 12860 29464 13185 29492
rect 12860 29452 12866 29464
rect 13173 29461 13185 29464
rect 13219 29461 13231 29495
rect 13173 29455 13231 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 3234 29248 3240 29300
rect 3292 29288 3298 29300
rect 4249 29291 4307 29297
rect 4249 29288 4261 29291
rect 3292 29260 4261 29288
rect 3292 29248 3298 29260
rect 3344 28960 3372 29260
rect 4249 29257 4261 29260
rect 4295 29288 4307 29291
rect 4341 29291 4399 29297
rect 4341 29288 4353 29291
rect 4295 29260 4353 29288
rect 4295 29257 4307 29260
rect 4249 29251 4307 29257
rect 4341 29257 4353 29260
rect 4387 29257 4399 29291
rect 4522 29288 4528 29300
rect 4483 29260 4528 29288
rect 4341 29251 4399 29257
rect 4522 29248 4528 29260
rect 4580 29248 4586 29300
rect 6822 29288 6828 29300
rect 6783 29260 6828 29288
rect 6822 29248 6828 29260
rect 6880 29248 6886 29300
rect 8478 29248 8484 29300
rect 8536 29288 8542 29300
rect 8665 29291 8723 29297
rect 8665 29288 8677 29291
rect 8536 29260 8677 29288
rect 8536 29248 8542 29260
rect 8665 29257 8677 29260
rect 8711 29257 8723 29291
rect 8665 29251 8723 29257
rect 9766 29248 9772 29300
rect 9824 29288 9830 29300
rect 10042 29288 10048 29300
rect 9824 29260 10048 29288
rect 9824 29248 9830 29260
rect 10042 29248 10048 29260
rect 10100 29288 10106 29300
rect 10229 29291 10287 29297
rect 10229 29288 10241 29291
rect 10100 29260 10241 29288
rect 10100 29248 10106 29260
rect 10229 29257 10241 29260
rect 10275 29257 10287 29291
rect 10594 29288 10600 29300
rect 10555 29260 10600 29288
rect 10229 29251 10287 29257
rect 10594 29248 10600 29260
rect 10652 29248 10658 29300
rect 12529 29291 12587 29297
rect 12529 29257 12541 29291
rect 12575 29288 12587 29291
rect 12894 29288 12900 29300
rect 12575 29260 12900 29288
rect 12575 29257 12587 29260
rect 12529 29251 12587 29257
rect 12894 29248 12900 29260
rect 12952 29248 12958 29300
rect 13446 29248 13452 29300
rect 13504 29288 13510 29300
rect 13541 29291 13599 29297
rect 13541 29288 13553 29291
rect 13504 29260 13553 29288
rect 13504 29248 13510 29260
rect 13541 29257 13553 29260
rect 13587 29257 13599 29291
rect 13541 29251 13599 29257
rect 6638 29220 6644 29232
rect 6551 29192 6644 29220
rect 6638 29180 6644 29192
rect 6696 29220 6702 29232
rect 9677 29223 9735 29229
rect 6696 29192 7512 29220
rect 6696 29180 6702 29192
rect 4065 29155 4123 29161
rect 4065 29121 4077 29155
rect 4111 29152 4123 29155
rect 4798 29152 4804 29164
rect 4111 29124 4804 29152
rect 4111 29121 4123 29124
rect 4065 29115 4123 29121
rect 4798 29112 4804 29124
rect 4856 29152 4862 29164
rect 5077 29155 5135 29161
rect 5077 29152 5089 29155
rect 4856 29124 5089 29152
rect 4856 29112 4862 29124
rect 5077 29121 5089 29124
rect 5123 29152 5135 29155
rect 5537 29155 5595 29161
rect 5537 29152 5549 29155
rect 5123 29124 5549 29152
rect 5123 29121 5135 29124
rect 5077 29115 5135 29121
rect 5537 29121 5549 29124
rect 5583 29121 5595 29155
rect 5537 29115 5595 29121
rect 6914 29112 6920 29164
rect 6972 29152 6978 29164
rect 7282 29152 7288 29164
rect 6972 29124 7288 29152
rect 6972 29112 6978 29124
rect 7282 29112 7288 29124
rect 7340 29112 7346 29164
rect 7484 29161 7512 29192
rect 9677 29189 9689 29223
rect 9723 29220 9735 29223
rect 10318 29220 10324 29232
rect 9723 29192 10324 29220
rect 9723 29189 9735 29192
rect 9677 29183 9735 29189
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29152 7527 29155
rect 8202 29152 8208 29164
rect 7515 29124 8208 29152
rect 7515 29121 7527 29124
rect 7469 29115 7527 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 8478 29152 8484 29164
rect 8439 29124 8484 29152
rect 8478 29112 8484 29124
rect 8536 29112 8542 29164
rect 8662 29112 8668 29164
rect 8720 29152 8726 29164
rect 9122 29152 9128 29164
rect 8720 29124 9128 29152
rect 8720 29112 8726 29124
rect 9122 29112 9128 29124
rect 9180 29152 9186 29164
rect 9217 29155 9275 29161
rect 9217 29152 9229 29155
rect 9180 29124 9229 29152
rect 9180 29112 9186 29124
rect 9217 29121 9229 29124
rect 9263 29152 9275 29155
rect 9692 29152 9720 29183
rect 10318 29180 10324 29192
rect 10376 29180 10382 29232
rect 10502 29180 10508 29232
rect 10560 29220 10566 29232
rect 11793 29223 11851 29229
rect 11793 29220 11805 29223
rect 10560 29192 11805 29220
rect 10560 29180 10566 29192
rect 11793 29189 11805 29192
rect 11839 29189 11851 29223
rect 11793 29183 11851 29189
rect 9263 29124 9720 29152
rect 9263 29121 9275 29124
rect 9217 29115 9275 29121
rect 9858 29112 9864 29164
rect 9916 29152 9922 29164
rect 10594 29152 10600 29164
rect 9916 29124 10600 29152
rect 9916 29112 9922 29124
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 11238 29152 11244 29164
rect 11199 29124 11244 29152
rect 11238 29112 11244 29124
rect 11296 29112 11302 29164
rect 11808 29152 11836 29183
rect 11974 29180 11980 29232
rect 12032 29220 12038 29232
rect 12161 29223 12219 29229
rect 12161 29220 12173 29223
rect 12032 29192 12173 29220
rect 12032 29180 12038 29192
rect 12161 29189 12173 29192
rect 12207 29189 12219 29223
rect 12161 29183 12219 29189
rect 12250 29152 12256 29164
rect 11808 29124 12256 29152
rect 12250 29112 12256 29124
rect 12308 29112 12314 29164
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 12860 29124 13093 29152
rect 12860 29112 12866 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 4893 29087 4951 29093
rect 4893 29053 4905 29087
rect 4939 29084 4951 29087
rect 5166 29084 5172 29096
rect 4939 29056 5172 29084
rect 4939 29053 4951 29056
rect 4893 29047 4951 29053
rect 5166 29044 5172 29056
rect 5224 29044 5230 29096
rect 6086 29044 6092 29096
rect 6144 29084 6150 29096
rect 6638 29084 6644 29096
rect 6144 29056 6644 29084
rect 6144 29044 6150 29056
rect 6638 29044 6644 29056
rect 6696 29044 6702 29096
rect 4249 29019 4307 29025
rect 4249 28985 4261 29019
rect 4295 29016 4307 29019
rect 4985 29019 5043 29025
rect 4985 29016 4997 29019
rect 4295 28988 4997 29016
rect 4295 28985 4307 28988
rect 4249 28979 4307 28985
rect 4985 28985 4997 28988
rect 5031 28985 5043 29019
rect 4985 28979 5043 28985
rect 6273 29019 6331 29025
rect 6273 28985 6285 29019
rect 6319 29016 6331 29019
rect 7190 29016 7196 29028
rect 6319 28988 7196 29016
rect 6319 28985 6331 28988
rect 6273 28979 6331 28985
rect 7190 28976 7196 28988
rect 7248 28976 7254 29028
rect 8113 29019 8171 29025
rect 8113 28985 8125 29019
rect 8159 29016 8171 29019
rect 8386 29016 8392 29028
rect 8159 28988 8392 29016
rect 8159 28985 8171 28988
rect 8113 28979 8171 28985
rect 8386 28976 8392 28988
rect 8444 28976 8450 29028
rect 8496 29016 8524 29112
rect 10318 29044 10324 29096
rect 10376 29084 10382 29096
rect 10413 29087 10471 29093
rect 10413 29084 10425 29087
rect 10376 29056 10425 29084
rect 10376 29044 10382 29056
rect 10413 29053 10425 29056
rect 10459 29053 10471 29087
rect 12894 29084 12900 29096
rect 12855 29056 12900 29084
rect 10413 29047 10471 29053
rect 12894 29044 12900 29056
rect 12952 29044 12958 29096
rect 9125 29019 9183 29025
rect 9125 29016 9137 29019
rect 8496 28988 9137 29016
rect 9125 28985 9137 28988
rect 9171 28985 9183 29019
rect 9125 28979 9183 28985
rect 9398 28976 9404 29028
rect 9456 29016 9462 29028
rect 10137 29019 10195 29025
rect 10137 29016 10149 29019
rect 9456 28988 10149 29016
rect 9456 28976 9462 28988
rect 10137 28985 10149 28988
rect 10183 29016 10195 29019
rect 10870 29016 10876 29028
rect 10183 28988 10876 29016
rect 10183 28985 10195 28988
rect 10137 28979 10195 28985
rect 10870 28976 10876 28988
rect 10928 29016 10934 29028
rect 10965 29019 11023 29025
rect 10965 29016 10977 29019
rect 10928 28988 10977 29016
rect 10928 28976 10934 28988
rect 10965 28985 10977 28988
rect 11011 28985 11023 29019
rect 12912 29016 12940 29044
rect 13446 29016 13452 29028
rect 12912 28988 13452 29016
rect 10965 28979 11023 28985
rect 13446 28976 13452 28988
rect 13504 28976 13510 29028
rect 14182 29016 14188 29028
rect 13740 28988 14188 29016
rect 3326 28908 3332 28960
rect 3384 28908 3390 28960
rect 8662 28908 8668 28960
rect 8720 28948 8726 28960
rect 9033 28951 9091 28957
rect 9033 28948 9045 28951
rect 8720 28920 9045 28948
rect 8720 28908 8726 28920
rect 9033 28917 9045 28920
rect 9079 28917 9091 28951
rect 9033 28911 9091 28917
rect 10410 28908 10416 28960
rect 10468 28948 10474 28960
rect 10502 28948 10508 28960
rect 10468 28920 10508 28948
rect 10468 28908 10474 28920
rect 10502 28908 10508 28920
rect 10560 28908 10566 28960
rect 10594 28908 10600 28960
rect 10652 28948 10658 28960
rect 11057 28951 11115 28957
rect 11057 28948 11069 28951
rect 10652 28920 11069 28948
rect 10652 28908 10658 28920
rect 11057 28917 11069 28920
rect 11103 28917 11115 28951
rect 11057 28911 11115 28917
rect 12894 28908 12900 28960
rect 12952 28948 12958 28960
rect 12989 28951 13047 28957
rect 12989 28948 13001 28951
rect 12952 28920 13001 28948
rect 12952 28908 12958 28920
rect 12989 28917 13001 28920
rect 13035 28948 13047 28951
rect 13740 28948 13768 28988
rect 14182 28976 14188 28988
rect 14240 28976 14246 29028
rect 13035 28920 13768 28948
rect 13035 28917 13047 28920
rect 12989 28911 13047 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 2958 28704 2964 28756
rect 3016 28744 3022 28756
rect 4062 28744 4068 28756
rect 3016 28716 4068 28744
rect 3016 28704 3022 28716
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 7190 28704 7196 28756
rect 7248 28744 7254 28756
rect 7285 28747 7343 28753
rect 7285 28744 7297 28747
rect 7248 28716 7297 28744
rect 7248 28704 7254 28716
rect 7285 28713 7297 28716
rect 7331 28713 7343 28747
rect 7285 28707 7343 28713
rect 8389 28747 8447 28753
rect 8389 28713 8401 28747
rect 8435 28744 8447 28747
rect 8570 28744 8576 28756
rect 8435 28716 8576 28744
rect 8435 28713 8447 28716
rect 8389 28707 8447 28713
rect 8570 28704 8576 28716
rect 8628 28704 8634 28756
rect 9122 28744 9128 28756
rect 9083 28716 9128 28744
rect 9122 28704 9128 28716
rect 9180 28704 9186 28756
rect 9953 28747 10011 28753
rect 9953 28713 9965 28747
rect 9999 28744 10011 28747
rect 10042 28744 10048 28756
rect 9999 28716 10048 28744
rect 9999 28713 10011 28716
rect 9953 28707 10011 28713
rect 10042 28704 10048 28716
rect 10100 28704 10106 28756
rect 10318 28744 10324 28756
rect 10279 28716 10324 28744
rect 10318 28704 10324 28716
rect 10376 28704 10382 28756
rect 10962 28704 10968 28756
rect 11020 28744 11026 28756
rect 11974 28744 11980 28756
rect 11020 28716 11980 28744
rect 11020 28704 11026 28716
rect 11974 28704 11980 28716
rect 12032 28704 12038 28756
rect 12526 28704 12532 28756
rect 12584 28744 12590 28756
rect 12897 28747 12955 28753
rect 12897 28744 12909 28747
rect 12584 28716 12909 28744
rect 12584 28704 12590 28716
rect 12897 28713 12909 28716
rect 12943 28713 12955 28747
rect 13078 28744 13084 28756
rect 13039 28716 13084 28744
rect 12897 28707 12955 28713
rect 13078 28704 13084 28716
rect 13136 28704 13142 28756
rect 7926 28676 7932 28688
rect 7208 28648 7932 28676
rect 7208 28617 7236 28648
rect 7926 28636 7932 28648
rect 7984 28636 7990 28688
rect 11146 28636 11152 28688
rect 11204 28676 11210 28688
rect 11885 28679 11943 28685
rect 11885 28676 11897 28679
rect 11204 28648 11897 28676
rect 11204 28636 11210 28648
rect 11885 28645 11897 28648
rect 11931 28645 11943 28679
rect 11885 28639 11943 28645
rect 6549 28611 6607 28617
rect 6549 28577 6561 28611
rect 6595 28608 6607 28611
rect 7193 28611 7251 28617
rect 7193 28608 7205 28611
rect 6595 28580 7205 28608
rect 6595 28577 6607 28580
rect 6549 28571 6607 28577
rect 7193 28577 7205 28580
rect 7239 28577 7251 28611
rect 7193 28571 7251 28577
rect 7653 28611 7711 28617
rect 7653 28577 7665 28611
rect 7699 28608 7711 28611
rect 8754 28608 8760 28620
rect 7699 28580 8760 28608
rect 7699 28577 7711 28580
rect 7653 28571 7711 28577
rect 8754 28568 8760 28580
rect 8812 28568 8818 28620
rect 11057 28611 11115 28617
rect 11057 28577 11069 28611
rect 11103 28608 11115 28611
rect 11238 28608 11244 28620
rect 11103 28580 11244 28608
rect 11103 28577 11115 28580
rect 11057 28571 11115 28577
rect 11238 28568 11244 28580
rect 11296 28568 11302 28620
rect 7742 28540 7748 28552
rect 7703 28512 7748 28540
rect 7742 28500 7748 28512
rect 7800 28500 7806 28552
rect 7834 28500 7840 28552
rect 7892 28540 7898 28552
rect 12158 28540 12164 28552
rect 7892 28512 7937 28540
rect 12119 28512 12164 28540
rect 7892 28500 7898 28512
rect 12158 28500 12164 28512
rect 12216 28500 12222 28552
rect 5166 28472 5172 28484
rect 4540 28444 5172 28472
rect 4338 28364 4344 28416
rect 4396 28404 4402 28416
rect 4540 28413 4568 28444
rect 5166 28432 5172 28444
rect 5224 28432 5230 28484
rect 6917 28475 6975 28481
rect 6917 28441 6929 28475
rect 6963 28472 6975 28475
rect 7098 28472 7104 28484
rect 6963 28444 7104 28472
rect 6963 28441 6975 28444
rect 6917 28435 6975 28441
rect 7098 28432 7104 28444
rect 7156 28472 7162 28484
rect 7852 28472 7880 28500
rect 7156 28444 7880 28472
rect 7156 28432 7162 28444
rect 10778 28432 10784 28484
rect 10836 28472 10842 28484
rect 11517 28475 11575 28481
rect 11517 28472 11529 28475
rect 10836 28444 11529 28472
rect 10836 28432 10842 28444
rect 11517 28441 11529 28444
rect 11563 28441 11575 28475
rect 11517 28435 11575 28441
rect 4525 28407 4583 28413
rect 4525 28404 4537 28407
rect 4396 28376 4537 28404
rect 4396 28364 4402 28376
rect 4525 28373 4537 28376
rect 4571 28373 4583 28407
rect 4982 28404 4988 28416
rect 4943 28376 4988 28404
rect 4525 28367 4583 28373
rect 4982 28364 4988 28376
rect 5040 28404 5046 28416
rect 6089 28407 6147 28413
rect 6089 28404 6101 28407
rect 5040 28376 6101 28404
rect 5040 28364 5046 28376
rect 6089 28373 6101 28376
rect 6135 28404 6147 28407
rect 6822 28404 6828 28416
rect 6135 28376 6828 28404
rect 6135 28373 6147 28376
rect 6089 28367 6147 28373
rect 6822 28364 6828 28376
rect 6880 28364 6886 28416
rect 7009 28407 7067 28413
rect 7009 28373 7021 28407
rect 7055 28404 7067 28407
rect 8110 28404 8116 28416
rect 7055 28376 8116 28404
rect 7055 28373 7067 28376
rect 7009 28367 7067 28373
rect 8110 28364 8116 28376
rect 8168 28364 8174 28416
rect 8570 28364 8576 28416
rect 8628 28404 8634 28416
rect 8665 28407 8723 28413
rect 8665 28404 8677 28407
rect 8628 28376 8677 28404
rect 8628 28364 8634 28376
rect 8665 28373 8677 28376
rect 8711 28373 8723 28407
rect 8665 28367 8723 28373
rect 10594 28364 10600 28416
rect 10652 28404 10658 28416
rect 10689 28407 10747 28413
rect 10689 28404 10701 28407
rect 10652 28376 10701 28404
rect 10652 28364 10658 28376
rect 10689 28373 10701 28376
rect 10735 28404 10747 28407
rect 10962 28404 10968 28416
rect 10735 28376 10968 28404
rect 10735 28373 10747 28376
rect 10689 28367 10747 28373
rect 10962 28364 10968 28376
rect 11020 28364 11026 28416
rect 12526 28404 12532 28416
rect 12487 28376 12532 28404
rect 12526 28364 12532 28376
rect 12584 28404 12590 28416
rect 12894 28404 12900 28416
rect 12584 28376 12900 28404
rect 12584 28364 12590 28376
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 6641 28203 6699 28209
rect 6641 28169 6653 28203
rect 6687 28200 6699 28203
rect 7742 28200 7748 28212
rect 6687 28172 7748 28200
rect 6687 28169 6699 28172
rect 6641 28163 6699 28169
rect 7742 28160 7748 28172
rect 7800 28160 7806 28212
rect 8202 28200 8208 28212
rect 8163 28172 8208 28200
rect 8202 28160 8208 28172
rect 8260 28160 8266 28212
rect 8754 28200 8760 28212
rect 8715 28172 8760 28200
rect 8754 28160 8760 28172
rect 8812 28160 8818 28212
rect 11146 28200 11152 28212
rect 11107 28172 11152 28200
rect 11146 28160 11152 28172
rect 11204 28160 11210 28212
rect 11974 28200 11980 28212
rect 11935 28172 11980 28200
rect 11974 28160 11980 28172
rect 12032 28160 12038 28212
rect 8772 28064 8800 28160
rect 11609 28135 11667 28141
rect 11609 28101 11621 28135
rect 11655 28132 11667 28135
rect 12158 28132 12164 28144
rect 11655 28104 12164 28132
rect 11655 28101 11667 28104
rect 11609 28095 11667 28101
rect 12158 28092 12164 28104
rect 12216 28092 12222 28144
rect 9309 28067 9367 28073
rect 9309 28064 9321 28067
rect 8772 28036 9321 28064
rect 9309 28033 9321 28036
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 11146 28024 11152 28076
rect 11204 28064 11210 28076
rect 11422 28064 11428 28076
rect 11204 28036 11428 28064
rect 11204 28024 11210 28036
rect 11422 28024 11428 28036
rect 11480 28024 11486 28076
rect 6822 27996 6828 28008
rect 6783 27968 6828 27996
rect 6822 27956 6828 27968
rect 6880 27956 6886 28008
rect 5721 27931 5779 27937
rect 5721 27897 5733 27931
rect 5767 27928 5779 27931
rect 6914 27928 6920 27940
rect 5767 27900 6920 27928
rect 5767 27897 5779 27900
rect 5721 27891 5779 27897
rect 6914 27888 6920 27900
rect 6972 27888 6978 27940
rect 7092 27931 7150 27937
rect 7092 27897 7104 27931
rect 7138 27928 7150 27931
rect 7834 27928 7840 27940
rect 7138 27900 7840 27928
rect 7138 27897 7150 27900
rect 7092 27891 7150 27897
rect 5350 27860 5356 27872
rect 5311 27832 5356 27860
rect 5350 27820 5356 27832
rect 5408 27820 5414 27872
rect 6273 27863 6331 27869
rect 6273 27829 6285 27863
rect 6319 27860 6331 27863
rect 7107 27860 7135 27891
rect 7834 27888 7840 27900
rect 7892 27888 7898 27940
rect 6319 27832 7135 27860
rect 6319 27829 6331 27832
rect 6273 27823 6331 27829
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 5350 27616 5356 27668
rect 5408 27656 5414 27668
rect 8110 27656 8116 27668
rect 5408 27628 5488 27656
rect 5408 27616 5414 27628
rect 1670 27588 1676 27600
rect 1631 27560 1676 27588
rect 1670 27548 1676 27560
rect 1728 27548 1734 27600
rect 5460 27588 5488 27628
rect 6840 27628 8116 27656
rect 6840 27588 6868 27628
rect 8110 27616 8116 27628
rect 8168 27616 8174 27668
rect 9125 27659 9183 27665
rect 9125 27625 9137 27659
rect 9171 27656 9183 27659
rect 10318 27656 10324 27668
rect 9171 27628 10324 27656
rect 9171 27625 9183 27628
rect 9125 27619 9183 27625
rect 5460 27560 6868 27588
rect 7653 27591 7711 27597
rect 5552 27529 5580 27560
rect 7653 27557 7665 27591
rect 7699 27588 7711 27591
rect 7742 27588 7748 27600
rect 7699 27560 7748 27588
rect 7699 27557 7711 27560
rect 7653 27551 7711 27557
rect 7742 27548 7748 27560
rect 7800 27548 7806 27600
rect 8846 27548 8852 27600
rect 8904 27588 8910 27600
rect 9140 27588 9168 27619
rect 10318 27616 10324 27628
rect 10376 27616 10382 27668
rect 12802 27656 12808 27668
rect 12763 27628 12808 27656
rect 12802 27616 12808 27628
rect 12860 27616 12866 27668
rect 8904 27560 9168 27588
rect 8904 27548 8910 27560
rect 11238 27548 11244 27600
rect 11296 27588 11302 27600
rect 11670 27591 11728 27597
rect 11670 27588 11682 27591
rect 11296 27560 11682 27588
rect 11296 27548 11302 27560
rect 11670 27557 11682 27560
rect 11716 27557 11728 27591
rect 11670 27551 11728 27557
rect 1397 27523 1455 27529
rect 1397 27489 1409 27523
rect 1443 27489 1455 27523
rect 1397 27483 1455 27489
rect 5537 27523 5595 27529
rect 5537 27489 5549 27523
rect 5583 27489 5595 27523
rect 5994 27520 6000 27532
rect 5955 27492 6000 27520
rect 5537 27483 5595 27489
rect 1412 27452 1440 27483
rect 5994 27480 6000 27492
rect 6052 27480 6058 27532
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 9309 27523 9367 27529
rect 9309 27520 9321 27523
rect 8168 27492 9321 27520
rect 8168 27480 8174 27492
rect 9309 27489 9321 27492
rect 9355 27520 9367 27523
rect 9674 27520 9680 27532
rect 9355 27492 9680 27520
rect 9355 27489 9367 27492
rect 9309 27483 9367 27489
rect 9674 27480 9680 27492
rect 9732 27480 9738 27532
rect 1670 27452 1676 27464
rect 1412 27424 1676 27452
rect 1670 27412 1676 27424
rect 1728 27412 1734 27464
rect 6086 27452 6092 27464
rect 5184 27424 5856 27452
rect 6047 27424 6092 27452
rect 5184 27328 5212 27424
rect 5353 27387 5411 27393
rect 5353 27353 5365 27387
rect 5399 27384 5411 27387
rect 5718 27384 5724 27396
rect 5399 27356 5724 27384
rect 5399 27353 5411 27356
rect 5353 27347 5411 27353
rect 5718 27344 5724 27356
rect 5776 27344 5782 27396
rect 5828 27384 5856 27424
rect 6086 27412 6092 27424
rect 6144 27412 6150 27464
rect 6181 27455 6239 27461
rect 6181 27421 6193 27455
rect 6227 27452 6239 27455
rect 6227 27424 6261 27452
rect 6227 27421 6239 27424
rect 6181 27415 6239 27421
rect 6196 27384 6224 27415
rect 7374 27412 7380 27464
rect 7432 27452 7438 27464
rect 7745 27455 7803 27461
rect 7745 27452 7757 27455
rect 7432 27424 7757 27452
rect 7432 27412 7438 27424
rect 7745 27421 7757 27424
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 7834 27412 7840 27464
rect 7892 27452 7898 27464
rect 11422 27452 11428 27464
rect 7892 27424 7937 27452
rect 11383 27424 11428 27452
rect 7892 27412 7898 27424
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 6822 27384 6828 27396
rect 5828 27356 6828 27384
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 7282 27384 7288 27396
rect 7243 27356 7288 27384
rect 7282 27344 7288 27356
rect 7340 27344 7346 27396
rect 5166 27316 5172 27328
rect 5127 27288 5172 27316
rect 5166 27276 5172 27288
rect 5224 27276 5230 27328
rect 5534 27276 5540 27328
rect 5592 27316 5598 27328
rect 5629 27319 5687 27325
rect 5629 27316 5641 27319
rect 5592 27288 5641 27316
rect 5592 27276 5598 27288
rect 5629 27285 5641 27288
rect 5675 27285 5687 27319
rect 8754 27316 8760 27328
rect 8715 27288 8760 27316
rect 5629 27279 5687 27285
rect 8754 27276 8760 27288
rect 8812 27276 8818 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 4798 27112 4804 27124
rect 4759 27084 4804 27112
rect 4798 27072 4804 27084
rect 4856 27072 4862 27124
rect 6086 27112 6092 27124
rect 6047 27084 6092 27112
rect 6086 27072 6092 27084
rect 6144 27072 6150 27124
rect 9674 27112 9680 27124
rect 9635 27084 9680 27112
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 11238 27072 11244 27124
rect 11296 27112 11302 27124
rect 11425 27115 11483 27121
rect 11425 27112 11437 27115
rect 11296 27084 11437 27112
rect 11296 27072 11302 27084
rect 11425 27081 11437 27084
rect 11471 27081 11483 27115
rect 11425 27075 11483 27081
rect 5721 27047 5779 27053
rect 5721 27013 5733 27047
rect 5767 27044 5779 27047
rect 5994 27044 6000 27056
rect 5767 27016 6000 27044
rect 5767 27013 5779 27016
rect 5721 27007 5779 27013
rect 5994 27004 6000 27016
rect 6052 27004 6058 27056
rect 10502 27004 10508 27056
rect 10560 27044 10566 27056
rect 12066 27044 12072 27056
rect 10560 27016 12072 27044
rect 10560 27004 10566 27016
rect 12066 27004 12072 27016
rect 12124 27004 12130 27056
rect 6822 26936 6828 26988
rect 6880 26976 6886 26988
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 6880 26948 7389 26976
rect 6880 26936 6886 26948
rect 7377 26945 7389 26948
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 8754 26936 8760 26988
rect 8812 26976 8818 26988
rect 9217 26979 9275 26985
rect 9217 26976 9229 26979
rect 8812 26948 9229 26976
rect 8812 26936 8818 26948
rect 9217 26945 9229 26948
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 3418 26908 3424 26920
rect 3379 26880 3424 26908
rect 3418 26868 3424 26880
rect 3476 26868 3482 26920
rect 6914 26868 6920 26920
rect 6972 26908 6978 26920
rect 7193 26911 7251 26917
rect 7193 26908 7205 26911
rect 6972 26880 7205 26908
rect 6972 26868 6978 26880
rect 7193 26877 7205 26880
rect 7239 26877 7251 26911
rect 7193 26871 7251 26877
rect 8662 26868 8668 26920
rect 8720 26908 8726 26920
rect 9030 26908 9036 26920
rect 8720 26880 9036 26908
rect 8720 26868 8726 26880
rect 9030 26868 9036 26880
rect 9088 26868 9094 26920
rect 3666 26843 3724 26849
rect 3666 26840 3678 26843
rect 3252 26812 3678 26840
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 2958 26732 2964 26784
rect 3016 26772 3022 26784
rect 3252 26781 3280 26812
rect 3666 26809 3678 26812
rect 3712 26809 3724 26843
rect 3666 26803 3724 26809
rect 6641 26843 6699 26849
rect 6641 26809 6653 26843
rect 6687 26840 6699 26843
rect 7282 26840 7288 26852
rect 6687 26812 7288 26840
rect 6687 26809 6699 26812
rect 6641 26803 6699 26809
rect 7282 26800 7288 26812
rect 7340 26800 7346 26852
rect 9125 26843 9183 26849
rect 9125 26840 9137 26843
rect 8496 26812 9137 26840
rect 3237 26775 3295 26781
rect 3237 26772 3249 26775
rect 3016 26744 3249 26772
rect 3016 26732 3022 26744
rect 3237 26741 3249 26744
rect 3283 26741 3295 26775
rect 6822 26772 6828 26784
rect 6783 26744 6828 26772
rect 3237 26735 3295 26741
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 7742 26732 7748 26784
rect 7800 26772 7806 26784
rect 7837 26775 7895 26781
rect 7837 26772 7849 26775
rect 7800 26744 7849 26772
rect 7800 26732 7806 26744
rect 7837 26741 7849 26744
rect 7883 26741 7895 26775
rect 7837 26735 7895 26741
rect 8202 26732 8208 26784
rect 8260 26772 8266 26784
rect 8386 26772 8392 26784
rect 8260 26744 8392 26772
rect 8260 26732 8266 26744
rect 8386 26732 8392 26744
rect 8444 26772 8450 26784
rect 8496 26781 8524 26812
rect 9125 26809 9137 26812
rect 9171 26809 9183 26843
rect 9125 26803 9183 26809
rect 8481 26775 8539 26781
rect 8481 26772 8493 26775
rect 8444 26744 8493 26772
rect 8444 26732 8450 26744
rect 8481 26741 8493 26744
rect 8527 26741 8539 26775
rect 8662 26772 8668 26784
rect 8623 26744 8668 26772
rect 8481 26735 8539 26741
rect 8662 26732 8668 26744
rect 8720 26732 8726 26784
rect 9030 26772 9036 26784
rect 8991 26744 9036 26772
rect 9030 26732 9036 26744
rect 9088 26732 9094 26784
rect 9766 26732 9772 26784
rect 9824 26772 9830 26784
rect 10686 26772 10692 26784
rect 9824 26744 10692 26772
rect 9824 26732 9830 26744
rect 10686 26732 10692 26744
rect 10744 26732 10750 26784
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 11422 26772 11428 26784
rect 11296 26744 11428 26772
rect 11296 26732 11302 26744
rect 11422 26732 11428 26744
rect 11480 26772 11486 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 11480 26744 11805 26772
rect 11480 26732 11486 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 11793 26735 11851 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 1670 26528 1676 26580
rect 1728 26568 1734 26580
rect 2409 26571 2467 26577
rect 2409 26568 2421 26571
rect 1728 26540 2421 26568
rect 1728 26528 1734 26540
rect 2409 26537 2421 26540
rect 2455 26537 2467 26571
rect 3418 26568 3424 26580
rect 3379 26540 3424 26568
rect 2409 26531 2467 26537
rect 3418 26528 3424 26540
rect 3476 26528 3482 26580
rect 6914 26568 6920 26580
rect 6875 26540 6920 26568
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 7374 26568 7380 26580
rect 7335 26540 7380 26568
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 7745 26571 7803 26577
rect 7745 26537 7757 26571
rect 7791 26568 7803 26571
rect 7834 26568 7840 26580
rect 7791 26540 7840 26568
rect 7791 26537 7803 26540
rect 7745 26531 7803 26537
rect 7834 26528 7840 26540
rect 7892 26528 7898 26580
rect 2774 26460 2780 26512
rect 2832 26500 2838 26512
rect 3970 26500 3976 26512
rect 2832 26472 3976 26500
rect 2832 26460 2838 26472
rect 3970 26460 3976 26472
rect 4028 26460 4034 26512
rect 4982 26500 4988 26512
rect 4895 26472 4988 26500
rect 2866 26392 2872 26444
rect 2924 26432 2930 26444
rect 4908 26441 4936 26472
rect 4982 26460 4988 26472
rect 5040 26500 5046 26512
rect 5626 26500 5632 26512
rect 5040 26472 5632 26500
rect 5040 26460 5046 26472
rect 5626 26460 5632 26472
rect 5684 26460 5690 26512
rect 10042 26460 10048 26512
rect 10100 26500 10106 26512
rect 10290 26503 10348 26509
rect 10290 26500 10302 26503
rect 10100 26472 10302 26500
rect 10100 26460 10106 26472
rect 10290 26469 10302 26472
rect 10336 26469 10348 26503
rect 10290 26463 10348 26469
rect 5166 26441 5172 26444
rect 4893 26435 4951 26441
rect 2924 26404 2969 26432
rect 2924 26392 2930 26404
rect 4893 26401 4905 26435
rect 4939 26401 4951 26435
rect 5160 26432 5172 26441
rect 5127 26404 5172 26432
rect 4893 26395 4951 26401
rect 5160 26395 5172 26404
rect 5166 26392 5172 26395
rect 5224 26392 5230 26444
rect 2958 26364 2964 26376
rect 2919 26336 2964 26364
rect 2958 26324 2964 26336
rect 3016 26324 3022 26376
rect 10045 26367 10103 26373
rect 10045 26333 10057 26367
rect 10091 26333 10103 26367
rect 10045 26327 10103 26333
rect 5902 26256 5908 26308
rect 5960 26296 5966 26308
rect 6273 26299 6331 26305
rect 6273 26296 6285 26299
rect 5960 26268 6285 26296
rect 5960 26256 5966 26268
rect 6273 26265 6285 26268
rect 6319 26265 6331 26299
rect 9030 26296 9036 26308
rect 6273 26259 6331 26265
rect 8680 26268 9036 26296
rect 8386 26188 8392 26240
rect 8444 26228 8450 26240
rect 8680 26237 8708 26268
rect 9030 26256 9036 26268
rect 9088 26256 9094 26308
rect 8665 26231 8723 26237
rect 8665 26228 8677 26231
rect 8444 26200 8677 26228
rect 8444 26188 8450 26200
rect 8665 26197 8677 26200
rect 8711 26197 8723 26231
rect 8665 26191 8723 26197
rect 9217 26231 9275 26237
rect 9217 26197 9229 26231
rect 9263 26228 9275 26231
rect 9306 26228 9312 26240
rect 9263 26200 9312 26228
rect 9263 26197 9275 26200
rect 9217 26191 9275 26197
rect 9306 26188 9312 26200
rect 9364 26228 9370 26240
rect 10060 26228 10088 26327
rect 11422 26296 11428 26308
rect 11383 26268 11428 26296
rect 11422 26256 11428 26268
rect 11480 26256 11486 26308
rect 10318 26228 10324 26240
rect 9364 26200 10324 26228
rect 9364 26188 9370 26200
rect 10318 26188 10324 26200
rect 10376 26188 10382 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 1765 26027 1823 26033
rect 1765 25993 1777 26027
rect 1811 26024 1823 26027
rect 2590 26024 2596 26036
rect 1811 25996 2596 26024
rect 1811 25993 1823 25996
rect 1765 25987 1823 25993
rect 2590 25984 2596 25996
rect 2648 25984 2654 26036
rect 3970 25984 3976 26036
rect 4028 26024 4034 26036
rect 5077 26027 5135 26033
rect 5077 26024 5089 26027
rect 4028 25996 5089 26024
rect 4028 25984 4034 25996
rect 5077 25993 5089 25996
rect 5123 25993 5135 26027
rect 5077 25987 5135 25993
rect 5626 25984 5632 26036
rect 5684 26024 5690 26036
rect 6089 26027 6147 26033
rect 6089 26024 6101 26027
rect 5684 25996 6101 26024
rect 5684 25984 5690 25996
rect 6089 25993 6101 25996
rect 6135 25993 6147 26027
rect 8754 26024 8760 26036
rect 8715 25996 8760 26024
rect 6089 25987 6147 25993
rect 8754 25984 8760 25996
rect 8812 25984 8818 26036
rect 8849 26027 8907 26033
rect 8849 25993 8861 26027
rect 8895 26024 8907 26027
rect 9306 26024 9312 26036
rect 8895 25996 9312 26024
rect 8895 25993 8907 25996
rect 8849 25987 8907 25993
rect 5166 25916 5172 25968
rect 5224 25956 5230 25968
rect 5224 25928 5764 25956
rect 5224 25916 5230 25928
rect 4617 25891 4675 25897
rect 4617 25857 4629 25891
rect 4663 25888 4675 25891
rect 5534 25888 5540 25900
rect 4663 25860 5540 25888
rect 4663 25857 4675 25860
rect 4617 25851 4675 25857
rect 5534 25848 5540 25860
rect 5592 25848 5598 25900
rect 5736 25897 5764 25928
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25888 5779 25891
rect 5902 25888 5908 25900
rect 5767 25860 5908 25888
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 5902 25848 5908 25860
rect 5960 25848 5966 25900
rect 9140 25897 9168 25996
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 9125 25891 9183 25897
rect 9125 25857 9137 25891
rect 9171 25857 9183 25891
rect 9125 25851 9183 25857
rect 2593 25823 2651 25829
rect 2593 25789 2605 25823
rect 2639 25820 2651 25823
rect 3418 25820 3424 25832
rect 2639 25792 3424 25820
rect 2639 25789 2651 25792
rect 2593 25783 2651 25789
rect 3418 25780 3424 25792
rect 3476 25780 3482 25832
rect 5445 25823 5503 25829
rect 5445 25789 5457 25823
rect 5491 25820 5503 25823
rect 6822 25820 6828 25832
rect 5491 25792 6828 25820
rect 5491 25789 5503 25792
rect 5445 25783 5503 25789
rect 5552 25764 5580 25792
rect 6822 25780 6828 25792
rect 6880 25780 6886 25832
rect 8846 25780 8852 25832
rect 8904 25820 8910 25832
rect 9033 25823 9091 25829
rect 9033 25820 9045 25823
rect 8904 25792 9045 25820
rect 8904 25780 8910 25792
rect 9033 25789 9045 25792
rect 9079 25789 9091 25823
rect 9033 25783 9091 25789
rect 2774 25712 2780 25764
rect 2832 25761 2838 25764
rect 2832 25755 2896 25761
rect 2832 25721 2850 25755
rect 2884 25721 2896 25755
rect 2832 25715 2896 25721
rect 2832 25712 2838 25715
rect 5534 25712 5540 25764
rect 5592 25712 5598 25764
rect 8754 25712 8760 25764
rect 8812 25752 8818 25764
rect 9398 25761 9404 25764
rect 9370 25755 9404 25761
rect 9370 25752 9382 25755
rect 8812 25724 9382 25752
rect 8812 25712 8818 25724
rect 9370 25721 9382 25724
rect 9456 25752 9462 25764
rect 9456 25724 9518 25752
rect 9370 25715 9404 25721
rect 9398 25712 9404 25715
rect 9456 25712 9462 25724
rect 2130 25684 2136 25696
rect 2091 25656 2136 25684
rect 2130 25644 2136 25656
rect 2188 25644 2194 25696
rect 2501 25687 2559 25693
rect 2501 25653 2513 25687
rect 2547 25684 2559 25687
rect 2958 25684 2964 25696
rect 2547 25656 2964 25684
rect 2547 25653 2559 25656
rect 2501 25647 2559 25653
rect 2958 25644 2964 25656
rect 3016 25684 3022 25696
rect 3973 25687 4031 25693
rect 3973 25684 3985 25687
rect 3016 25656 3985 25684
rect 3016 25644 3022 25656
rect 3973 25653 3985 25656
rect 4019 25653 4031 25687
rect 3973 25647 4031 25653
rect 4985 25687 5043 25693
rect 4985 25653 4997 25687
rect 5031 25684 5043 25687
rect 5258 25684 5264 25696
rect 5031 25656 5264 25684
rect 5031 25653 5043 25656
rect 4985 25647 5043 25653
rect 5258 25644 5264 25656
rect 5316 25644 5322 25696
rect 8113 25687 8171 25693
rect 8113 25653 8125 25687
rect 8159 25684 8171 25687
rect 8478 25684 8484 25696
rect 8159 25656 8484 25684
rect 8159 25653 8171 25656
rect 8113 25647 8171 25653
rect 8478 25644 8484 25656
rect 8536 25644 8542 25696
rect 10505 25687 10563 25693
rect 10505 25653 10517 25687
rect 10551 25684 10563 25687
rect 10778 25684 10784 25696
rect 10551 25656 10784 25684
rect 10551 25653 10563 25656
rect 10505 25647 10563 25653
rect 10778 25644 10784 25656
rect 10836 25644 10842 25696
rect 11149 25687 11207 25693
rect 11149 25653 11161 25687
rect 11195 25684 11207 25687
rect 11238 25684 11244 25696
rect 11195 25656 11244 25684
rect 11195 25653 11207 25656
rect 11149 25647 11207 25653
rect 11238 25644 11244 25656
rect 11296 25644 11302 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 2130 25440 2136 25492
rect 2188 25480 2194 25492
rect 2866 25480 2872 25492
rect 2188 25452 2872 25480
rect 2188 25440 2194 25452
rect 2866 25440 2872 25452
rect 2924 25480 2930 25492
rect 4065 25483 4123 25489
rect 4065 25480 4077 25483
rect 2924 25452 4077 25480
rect 2924 25440 2930 25452
rect 4065 25449 4077 25452
rect 4111 25449 4123 25483
rect 5166 25480 5172 25492
rect 5127 25452 5172 25480
rect 4065 25443 4123 25449
rect 5166 25440 5172 25452
rect 5224 25440 5230 25492
rect 5534 25480 5540 25492
rect 5495 25452 5540 25480
rect 5534 25440 5540 25452
rect 5592 25440 5598 25492
rect 8478 25480 8484 25492
rect 8439 25452 8484 25480
rect 8478 25440 8484 25452
rect 8536 25440 8542 25492
rect 8846 25440 8852 25492
rect 8904 25480 8910 25492
rect 9033 25483 9091 25489
rect 9033 25480 9045 25483
rect 8904 25452 9045 25480
rect 8904 25440 8910 25452
rect 9033 25449 9045 25452
rect 9079 25449 9091 25483
rect 9033 25443 9091 25449
rect 2685 25415 2743 25421
rect 2685 25381 2697 25415
rect 2731 25412 2743 25415
rect 2774 25412 2780 25424
rect 2731 25384 2780 25412
rect 2731 25381 2743 25384
rect 2685 25375 2743 25381
rect 2774 25372 2780 25384
rect 2832 25412 2838 25424
rect 7561 25415 7619 25421
rect 2832 25384 4660 25412
rect 2832 25372 2838 25384
rect 3053 25347 3111 25353
rect 3053 25313 3065 25347
rect 3099 25344 3111 25347
rect 3418 25344 3424 25356
rect 3099 25316 3424 25344
rect 3099 25313 3111 25316
rect 3053 25307 3111 25313
rect 3418 25304 3424 25316
rect 3476 25304 3482 25356
rect 4430 25344 4436 25356
rect 4391 25316 4436 25344
rect 4430 25304 4436 25316
rect 4488 25304 4494 25356
rect 3436 25208 3464 25304
rect 4632 25288 4660 25384
rect 7561 25381 7573 25415
rect 7607 25412 7619 25415
rect 8389 25415 8447 25421
rect 8389 25412 8401 25415
rect 7607 25384 8401 25412
rect 7607 25381 7619 25384
rect 7561 25375 7619 25381
rect 8389 25381 8401 25384
rect 8435 25412 8447 25415
rect 8662 25412 8668 25424
rect 8435 25384 8668 25412
rect 8435 25381 8447 25384
rect 8389 25375 8447 25381
rect 8662 25372 8668 25384
rect 8720 25372 8726 25424
rect 11238 25412 11244 25424
rect 10428 25384 11244 25412
rect 5718 25304 5724 25356
rect 5776 25344 5782 25356
rect 5813 25347 5871 25353
rect 5813 25344 5825 25347
rect 5776 25316 5825 25344
rect 5776 25304 5782 25316
rect 5813 25313 5825 25316
rect 5859 25344 5871 25347
rect 6086 25344 6092 25356
rect 5859 25316 6092 25344
rect 5859 25313 5871 25316
rect 5813 25307 5871 25313
rect 6086 25304 6092 25316
rect 6144 25304 6150 25356
rect 8202 25304 8208 25356
rect 8260 25344 8266 25356
rect 8754 25344 8760 25356
rect 8260 25316 8760 25344
rect 8260 25304 8266 25316
rect 8754 25304 8760 25316
rect 8812 25304 8818 25356
rect 4522 25276 4528 25288
rect 4483 25248 4528 25276
rect 4522 25236 4528 25248
rect 4580 25236 4586 25288
rect 4614 25236 4620 25288
rect 4672 25276 4678 25288
rect 4709 25279 4767 25285
rect 4709 25276 4721 25279
rect 4672 25248 4721 25276
rect 4672 25236 4678 25248
rect 4709 25245 4721 25248
rect 4755 25276 4767 25279
rect 5166 25276 5172 25288
rect 4755 25248 5172 25276
rect 4755 25245 4767 25248
rect 4709 25239 4767 25245
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 7929 25279 7987 25285
rect 7929 25245 7941 25279
rect 7975 25276 7987 25279
rect 8662 25276 8668 25288
rect 7975 25248 8668 25276
rect 7975 25245 7987 25248
rect 7929 25239 7987 25245
rect 8662 25236 8668 25248
rect 8720 25236 8726 25288
rect 10318 25276 10324 25288
rect 10231 25248 10324 25276
rect 10318 25236 10324 25248
rect 10376 25276 10382 25288
rect 10428 25276 10456 25384
rect 11238 25372 11244 25384
rect 11296 25372 11302 25424
rect 10594 25353 10600 25356
rect 10588 25307 10600 25353
rect 10652 25344 10658 25356
rect 10652 25316 10688 25344
rect 10594 25304 10600 25307
rect 10652 25304 10658 25316
rect 10376 25248 10456 25276
rect 10376 25236 10382 25248
rect 5629 25211 5687 25217
rect 5629 25208 5641 25211
rect 3436 25180 5641 25208
rect 5629 25177 5641 25180
rect 5675 25208 5687 25211
rect 6178 25208 6184 25220
rect 5675 25180 6184 25208
rect 5675 25177 5687 25180
rect 5629 25171 5687 25177
rect 6178 25168 6184 25180
rect 6236 25168 6242 25220
rect 7650 25168 7656 25220
rect 7708 25208 7714 25220
rect 8021 25211 8079 25217
rect 8021 25208 8033 25211
rect 7708 25180 8033 25208
rect 7708 25168 7714 25180
rect 8021 25177 8033 25180
rect 8067 25177 8079 25211
rect 8021 25171 8079 25177
rect 7193 25143 7251 25149
rect 7193 25109 7205 25143
rect 7239 25140 7251 25143
rect 7282 25140 7288 25152
rect 7239 25112 7288 25140
rect 7239 25109 7251 25112
rect 7193 25103 7251 25109
rect 7282 25100 7288 25112
rect 7340 25100 7346 25152
rect 9674 25100 9680 25152
rect 9732 25140 9738 25152
rect 9858 25140 9864 25152
rect 9732 25112 9864 25140
rect 9732 25100 9738 25112
rect 9858 25100 9864 25112
rect 9916 25100 9922 25152
rect 10042 25140 10048 25152
rect 10003 25112 10048 25140
rect 10042 25100 10048 25112
rect 10100 25140 10106 25152
rect 11701 25143 11759 25149
rect 11701 25140 11713 25143
rect 10100 25112 11713 25140
rect 10100 25100 10106 25112
rect 11701 25109 11713 25112
rect 11747 25109 11759 25143
rect 11701 25103 11759 25109
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 4430 24896 4436 24948
rect 4488 24936 4494 24948
rect 4709 24939 4767 24945
rect 4709 24936 4721 24939
rect 4488 24908 4721 24936
rect 4488 24896 4494 24908
rect 4709 24905 4721 24908
rect 4755 24905 4767 24939
rect 6086 24936 6092 24948
rect 6047 24908 6092 24936
rect 4709 24899 4767 24905
rect 6086 24896 6092 24908
rect 6144 24896 6150 24948
rect 8478 24896 8484 24948
rect 8536 24936 8542 24948
rect 8757 24939 8815 24945
rect 8757 24936 8769 24939
rect 8536 24908 8769 24936
rect 8536 24896 8542 24908
rect 8757 24905 8769 24908
rect 8803 24905 8815 24939
rect 8757 24899 8815 24905
rect 3881 24871 3939 24877
rect 3881 24837 3893 24871
rect 3927 24868 3939 24871
rect 4614 24868 4620 24880
rect 3927 24840 4620 24868
rect 3927 24837 3939 24840
rect 3881 24831 3939 24837
rect 4614 24828 4620 24840
rect 4672 24828 4678 24880
rect 9416 24840 10916 24868
rect 9416 24812 9444 24840
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 4249 24803 4307 24809
rect 4249 24769 4261 24803
rect 4295 24800 4307 24803
rect 5258 24800 5264 24812
rect 4295 24772 5264 24800
rect 4295 24769 4307 24772
rect 4249 24763 4307 24769
rect 5258 24760 5264 24772
rect 5316 24760 5322 24812
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24800 6699 24803
rect 7650 24800 7656 24812
rect 6687 24772 7656 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 7650 24760 7656 24772
rect 7708 24760 7714 24812
rect 7745 24803 7803 24809
rect 7745 24769 7757 24803
rect 7791 24769 7803 24803
rect 7745 24763 7803 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 3513 24735 3571 24741
rect 1443 24704 2268 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 2240 24605 2268 24704
rect 3513 24701 3525 24735
rect 3559 24732 3571 24735
rect 4522 24732 4528 24744
rect 3559 24704 4528 24732
rect 3559 24701 3571 24704
rect 3513 24695 3571 24701
rect 4522 24692 4528 24704
rect 4580 24692 4586 24744
rect 7760 24732 7788 24763
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 8573 24803 8631 24809
rect 8573 24800 8585 24803
rect 8444 24772 8585 24800
rect 8444 24760 8450 24772
rect 8573 24769 8585 24772
rect 8619 24800 8631 24803
rect 9217 24803 9275 24809
rect 9217 24800 9229 24803
rect 8619 24772 9229 24800
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 9217 24769 9229 24772
rect 9263 24769 9275 24803
rect 9398 24800 9404 24812
rect 9359 24772 9404 24800
rect 9217 24763 9275 24769
rect 9398 24760 9404 24772
rect 9456 24760 9462 24812
rect 9858 24760 9864 24812
rect 9916 24800 9922 24812
rect 10888 24809 10916 24840
rect 10137 24803 10195 24809
rect 10137 24800 10149 24803
rect 9916 24772 10149 24800
rect 9916 24760 9922 24772
rect 10137 24769 10149 24772
rect 10183 24800 10195 24803
rect 10781 24803 10839 24809
rect 10781 24800 10793 24803
rect 10183 24772 10793 24800
rect 10183 24769 10195 24772
rect 10137 24763 10195 24769
rect 10781 24769 10793 24772
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10873 24803 10931 24809
rect 10873 24769 10885 24803
rect 10919 24800 10931 24803
rect 11333 24803 11391 24809
rect 11333 24800 11345 24803
rect 10919 24772 11345 24800
rect 10919 24769 10931 24772
rect 10873 24763 10931 24769
rect 11333 24769 11345 24772
rect 11379 24800 11391 24803
rect 11422 24800 11428 24812
rect 11379 24772 11428 24800
rect 11379 24769 11391 24772
rect 11333 24763 11391 24769
rect 11422 24760 11428 24772
rect 11480 24760 11486 24812
rect 7024 24704 7788 24732
rect 4246 24624 4252 24676
rect 4304 24664 4310 24676
rect 4617 24667 4675 24673
rect 4617 24664 4629 24667
rect 4304 24636 4629 24664
rect 4304 24624 4310 24636
rect 4617 24633 4629 24636
rect 4663 24664 4675 24667
rect 5077 24667 5135 24673
rect 5077 24664 5089 24667
rect 4663 24636 5089 24664
rect 4663 24633 4675 24636
rect 4617 24627 4675 24633
rect 5077 24633 5089 24636
rect 5123 24664 5135 24667
rect 5442 24664 5448 24676
rect 5123 24636 5448 24664
rect 5123 24633 5135 24636
rect 5077 24627 5135 24633
rect 5442 24624 5448 24636
rect 5500 24624 5506 24676
rect 2225 24599 2283 24605
rect 2225 24565 2237 24599
rect 2271 24596 2283 24599
rect 2406 24596 2412 24608
rect 2271 24568 2412 24596
rect 2271 24565 2283 24568
rect 2225 24559 2283 24565
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5224 24568 5733 24596
rect 5224 24556 5230 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 5721 24559 5779 24565
rect 6914 24556 6920 24608
rect 6972 24596 6978 24608
rect 7024 24605 7052 24704
rect 9861 24667 9919 24673
rect 9861 24633 9873 24667
rect 9907 24664 9919 24667
rect 10410 24664 10416 24676
rect 9907 24636 10416 24664
rect 9907 24633 9919 24636
rect 9861 24627 9919 24633
rect 10410 24624 10416 24636
rect 10468 24664 10474 24676
rect 10689 24667 10747 24673
rect 10689 24664 10701 24667
rect 10468 24636 10701 24664
rect 10468 24624 10474 24636
rect 10689 24633 10701 24636
rect 10735 24664 10747 24667
rect 11330 24664 11336 24676
rect 10735 24636 11336 24664
rect 10735 24633 10747 24636
rect 10689 24627 10747 24633
rect 11330 24624 11336 24636
rect 11388 24624 11394 24676
rect 7009 24599 7067 24605
rect 7009 24596 7021 24599
rect 6972 24568 7021 24596
rect 6972 24556 6978 24568
rect 7009 24565 7021 24568
rect 7055 24565 7067 24599
rect 7190 24596 7196 24608
rect 7151 24568 7196 24596
rect 7009 24559 7067 24565
rect 7190 24556 7196 24568
rect 7248 24556 7254 24608
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 7561 24599 7619 24605
rect 7561 24596 7573 24599
rect 7340 24568 7573 24596
rect 7340 24556 7346 24568
rect 7561 24565 7573 24568
rect 7607 24596 7619 24599
rect 7650 24596 7656 24608
rect 7607 24568 7656 24596
rect 7607 24565 7619 24568
rect 7561 24559 7619 24565
rect 7650 24556 7656 24568
rect 7708 24556 7714 24608
rect 8297 24599 8355 24605
rect 8297 24565 8309 24599
rect 8343 24596 8355 24599
rect 8570 24596 8576 24608
rect 8343 24568 8576 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 8570 24556 8576 24568
rect 8628 24596 8634 24608
rect 9125 24599 9183 24605
rect 9125 24596 9137 24599
rect 8628 24568 9137 24596
rect 8628 24556 8634 24568
rect 9125 24565 9137 24568
rect 9171 24596 9183 24599
rect 9490 24596 9496 24608
rect 9171 24568 9496 24596
rect 9171 24565 9183 24568
rect 9125 24559 9183 24565
rect 9490 24556 9496 24568
rect 9548 24556 9554 24608
rect 10318 24596 10324 24608
rect 10279 24568 10324 24596
rect 10318 24556 10324 24568
rect 10376 24556 10382 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 4341 24395 4399 24401
rect 4341 24361 4353 24395
rect 4387 24392 4399 24395
rect 4430 24392 4436 24404
rect 4387 24364 4436 24392
rect 4387 24361 4399 24364
rect 4341 24355 4399 24361
rect 4430 24352 4436 24364
rect 4488 24352 4494 24404
rect 4522 24352 4528 24404
rect 4580 24392 4586 24404
rect 4709 24395 4767 24401
rect 4709 24392 4721 24395
rect 4580 24364 4721 24392
rect 4580 24352 4586 24364
rect 4709 24361 4721 24364
rect 4755 24361 4767 24395
rect 4709 24355 4767 24361
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 9398 24392 9404 24404
rect 9171 24364 9404 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9398 24352 9404 24364
rect 9456 24352 9462 24404
rect 9674 24392 9680 24404
rect 9635 24364 9680 24392
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 10594 24352 10600 24404
rect 10652 24392 10658 24404
rect 10689 24395 10747 24401
rect 10689 24392 10701 24395
rect 10652 24364 10701 24392
rect 10652 24352 10658 24364
rect 10689 24361 10701 24364
rect 10735 24361 10747 24395
rect 10689 24355 10747 24361
rect 3970 24216 3976 24268
rect 4028 24256 4034 24268
rect 5077 24259 5135 24265
rect 5077 24256 5089 24259
rect 4028 24228 5089 24256
rect 4028 24216 4034 24228
rect 5077 24225 5089 24228
rect 5123 24256 5135 24259
rect 5534 24256 5540 24268
rect 5123 24228 5540 24256
rect 5123 24225 5135 24228
rect 5077 24219 5135 24225
rect 5534 24216 5540 24228
rect 5592 24216 5598 24268
rect 6822 24216 6828 24268
rect 6880 24256 6886 24268
rect 7368 24259 7426 24265
rect 7368 24256 7380 24259
rect 6880 24228 7380 24256
rect 6880 24216 6886 24228
rect 7368 24225 7380 24228
rect 7414 24256 7426 24259
rect 8662 24256 8668 24268
rect 7414 24228 8668 24256
rect 7414 24225 7426 24228
rect 7368 24219 7426 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 9674 24216 9680 24268
rect 9732 24256 9738 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9732 24228 10057 24256
rect 9732 24216 9738 24228
rect 10045 24225 10057 24228
rect 10091 24225 10103 24259
rect 10045 24219 10103 24225
rect 10137 24259 10195 24265
rect 10137 24225 10149 24259
rect 10183 24256 10195 24259
rect 10318 24256 10324 24268
rect 10183 24228 10324 24256
rect 10183 24225 10195 24228
rect 10137 24219 10195 24225
rect 4246 24148 4252 24200
rect 4304 24188 4310 24200
rect 5169 24191 5227 24197
rect 5169 24188 5181 24191
rect 4304 24160 5181 24188
rect 4304 24148 4310 24160
rect 5092 24132 5120 24160
rect 5169 24157 5181 24160
rect 5215 24157 5227 24191
rect 5169 24151 5227 24157
rect 5258 24148 5264 24200
rect 5316 24188 5322 24200
rect 5316 24160 5361 24188
rect 5316 24148 5322 24160
rect 6178 24148 6184 24200
rect 6236 24188 6242 24200
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 6236 24160 7113 24188
rect 6236 24148 6242 24160
rect 7101 24157 7113 24160
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 5074 24080 5080 24132
rect 5132 24080 5138 24132
rect 10060 24120 10088 24219
rect 10318 24216 10324 24228
rect 10376 24256 10382 24268
rect 10870 24256 10876 24268
rect 10376 24228 10876 24256
rect 10376 24216 10382 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10778 24188 10784 24200
rect 10275 24160 10784 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 10318 24120 10324 24132
rect 10060 24092 10324 24120
rect 10318 24080 10324 24092
rect 10376 24080 10382 24132
rect 6914 24052 6920 24064
rect 6875 24024 6920 24052
rect 6914 24012 6920 24024
rect 6972 24052 6978 24064
rect 8481 24055 8539 24061
rect 8481 24052 8493 24055
rect 6972 24024 8493 24052
rect 6972 24012 6978 24024
rect 8481 24021 8493 24024
rect 8527 24021 8539 24055
rect 8481 24015 8539 24021
rect 11149 24055 11207 24061
rect 11149 24021 11161 24055
rect 11195 24052 11207 24055
rect 11238 24052 11244 24064
rect 11195 24024 11244 24052
rect 11195 24021 11207 24024
rect 11149 24015 11207 24021
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 3881 23851 3939 23857
rect 3881 23817 3893 23851
rect 3927 23848 3939 23851
rect 3970 23848 3976 23860
rect 3927 23820 3976 23848
rect 3927 23817 3939 23820
rect 3881 23811 3939 23817
rect 3970 23808 3976 23820
rect 4028 23808 4034 23860
rect 4246 23848 4252 23860
rect 4207 23820 4252 23848
rect 4246 23808 4252 23820
rect 4304 23808 4310 23860
rect 4798 23808 4804 23860
rect 4856 23848 4862 23860
rect 4893 23851 4951 23857
rect 4893 23848 4905 23851
rect 4856 23820 4905 23848
rect 4856 23808 4862 23820
rect 4893 23817 4905 23820
rect 4939 23817 4951 23851
rect 4893 23811 4951 23817
rect 5077 23851 5135 23857
rect 5077 23817 5089 23851
rect 5123 23848 5135 23851
rect 5166 23848 5172 23860
rect 5123 23820 5172 23848
rect 5123 23817 5135 23820
rect 5077 23811 5135 23817
rect 5166 23808 5172 23820
rect 5224 23808 5230 23860
rect 6178 23848 6184 23860
rect 6139 23820 6184 23848
rect 6178 23808 6184 23820
rect 6236 23848 6242 23860
rect 6641 23851 6699 23857
rect 6236 23820 6592 23848
rect 6236 23808 6242 23820
rect 4617 23783 4675 23789
rect 4617 23749 4629 23783
rect 4663 23780 4675 23783
rect 5350 23780 5356 23792
rect 4663 23752 5356 23780
rect 4663 23749 4675 23752
rect 4617 23743 4675 23749
rect 5350 23740 5356 23752
rect 5408 23780 5414 23792
rect 5408 23752 5672 23780
rect 5408 23740 5414 23752
rect 4798 23672 4804 23724
rect 4856 23712 4862 23724
rect 5644 23721 5672 23752
rect 5537 23715 5595 23721
rect 5537 23712 5549 23715
rect 4856 23684 5549 23712
rect 4856 23672 4862 23684
rect 5537 23681 5549 23684
rect 5583 23681 5595 23715
rect 5537 23675 5595 23681
rect 5629 23715 5687 23721
rect 5629 23681 5641 23715
rect 5675 23681 5687 23715
rect 6564 23712 6592 23820
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 6822 23848 6828 23860
rect 6687 23820 6828 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 6822 23808 6828 23820
rect 6880 23808 6886 23860
rect 9858 23808 9864 23860
rect 9916 23848 9922 23860
rect 10137 23851 10195 23857
rect 10137 23848 10149 23851
rect 9916 23820 10149 23848
rect 9916 23808 9922 23820
rect 10137 23817 10149 23820
rect 10183 23817 10195 23851
rect 10137 23811 10195 23817
rect 10781 23851 10839 23857
rect 10781 23817 10793 23851
rect 10827 23848 10839 23851
rect 10870 23848 10876 23860
rect 10827 23820 10876 23848
rect 10827 23817 10839 23820
rect 10781 23811 10839 23817
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 9309 23783 9367 23789
rect 9309 23780 9321 23783
rect 8076 23752 9321 23780
rect 8076 23740 8082 23752
rect 9309 23749 9321 23752
rect 9355 23749 9367 23783
rect 9309 23743 9367 23749
rect 6825 23715 6883 23721
rect 6825 23712 6837 23715
rect 6564 23684 6837 23712
rect 5629 23675 5687 23681
rect 6825 23681 6837 23684
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 5552 23644 5580 23675
rect 8386 23672 8392 23724
rect 8444 23712 8450 23724
rect 8662 23712 8668 23724
rect 8444 23684 8668 23712
rect 8444 23672 8450 23684
rect 8662 23672 8668 23684
rect 8720 23712 8726 23724
rect 8849 23715 8907 23721
rect 8849 23712 8861 23715
rect 8720 23684 8861 23712
rect 8720 23672 8726 23684
rect 8849 23681 8861 23684
rect 8895 23712 8907 23715
rect 9858 23712 9864 23724
rect 8895 23684 9864 23712
rect 8895 23681 8907 23684
rect 8849 23675 8907 23681
rect 9858 23672 9864 23684
rect 9916 23712 9922 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9916 23684 9965 23712
rect 9916 23672 9922 23684
rect 9953 23681 9965 23684
rect 9999 23712 10011 23715
rect 10778 23712 10784 23724
rect 9999 23684 10784 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 5994 23644 6000 23656
rect 5552 23616 6000 23644
rect 5994 23604 6000 23616
rect 6052 23604 6058 23656
rect 9217 23647 9275 23653
rect 9217 23613 9229 23647
rect 9263 23644 9275 23647
rect 9674 23644 9680 23656
rect 9263 23616 9680 23644
rect 9263 23613 9275 23616
rect 9217 23607 9275 23613
rect 9674 23604 9680 23616
rect 9732 23644 9738 23656
rect 10226 23644 10232 23656
rect 9732 23616 10232 23644
rect 9732 23604 9738 23616
rect 10226 23604 10232 23616
rect 10284 23604 10290 23656
rect 6914 23536 6920 23588
rect 6972 23576 6978 23588
rect 7092 23579 7150 23585
rect 7092 23576 7104 23579
rect 6972 23548 7104 23576
rect 6972 23536 6978 23548
rect 7092 23545 7104 23548
rect 7138 23576 7150 23579
rect 7650 23576 7656 23588
rect 7138 23548 7656 23576
rect 7138 23545 7150 23548
rect 7092 23539 7150 23545
rect 7650 23536 7656 23548
rect 7708 23536 7714 23588
rect 9582 23576 9588 23588
rect 7760 23548 9588 23576
rect 5166 23468 5172 23520
rect 5224 23508 5230 23520
rect 5445 23511 5503 23517
rect 5445 23508 5457 23511
rect 5224 23480 5457 23508
rect 5224 23468 5230 23480
rect 5445 23477 5457 23480
rect 5491 23508 5503 23511
rect 7466 23508 7472 23520
rect 5491 23480 7472 23508
rect 5491 23477 5503 23480
rect 5445 23471 5503 23477
rect 7466 23468 7472 23480
rect 7524 23508 7530 23520
rect 7760 23508 7788 23548
rect 9582 23536 9588 23548
rect 9640 23536 9646 23588
rect 10778 23536 10784 23588
rect 10836 23576 10842 23588
rect 11054 23576 11060 23588
rect 10836 23548 11060 23576
rect 10836 23536 10842 23548
rect 11054 23536 11060 23548
rect 11112 23536 11118 23588
rect 7524 23480 7788 23508
rect 7524 23468 7530 23480
rect 8110 23468 8116 23520
rect 8168 23508 8174 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 8168 23480 8217 23508
rect 8168 23468 8174 23480
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 8205 23471 8263 23477
rect 9306 23468 9312 23520
rect 9364 23508 9370 23520
rect 9769 23511 9827 23517
rect 9769 23508 9781 23511
rect 9364 23480 9781 23508
rect 9364 23468 9370 23480
rect 9769 23477 9781 23480
rect 9815 23508 9827 23511
rect 10137 23511 10195 23517
rect 10137 23508 10149 23511
rect 9815 23480 10149 23508
rect 9815 23477 9827 23480
rect 9769 23471 9827 23477
rect 10137 23477 10149 23480
rect 10183 23477 10195 23511
rect 10318 23508 10324 23520
rect 10279 23480 10324 23508
rect 10137 23471 10195 23477
rect 10318 23468 10324 23480
rect 10376 23468 10382 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 4801 23307 4859 23313
rect 4801 23273 4813 23307
rect 4847 23304 4859 23307
rect 5258 23304 5264 23316
rect 4847 23276 5264 23304
rect 4847 23273 4859 23276
rect 4801 23267 4859 23273
rect 5258 23264 5264 23276
rect 5316 23304 5322 23316
rect 6733 23307 6791 23313
rect 6733 23304 6745 23307
rect 5316 23276 6745 23304
rect 5316 23264 5322 23276
rect 6733 23273 6745 23276
rect 6779 23273 6791 23307
rect 6733 23267 6791 23273
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 8294 23304 8300 23316
rect 7248 23276 8300 23304
rect 7248 23264 7254 23276
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 5166 23236 5172 23248
rect 5127 23208 5172 23236
rect 5166 23196 5172 23208
rect 5224 23196 5230 23248
rect 5350 23196 5356 23248
rect 5408 23236 5414 23248
rect 5598 23239 5656 23245
rect 5598 23236 5610 23239
rect 5408 23208 5610 23236
rect 5408 23196 5414 23208
rect 5598 23205 5610 23208
rect 5644 23205 5656 23239
rect 5598 23199 5656 23205
rect 11330 23196 11336 23248
rect 11388 23245 11394 23248
rect 11388 23239 11452 23245
rect 11388 23205 11406 23239
rect 11440 23205 11452 23239
rect 11388 23199 11452 23205
rect 11388 23196 11394 23199
rect 6178 23168 6184 23180
rect 5368 23140 6184 23168
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 5368 23109 5396 23140
rect 6178 23128 6184 23140
rect 6236 23168 6242 23180
rect 7285 23171 7343 23177
rect 7285 23168 7297 23171
rect 6236 23140 7297 23168
rect 6236 23128 6242 23140
rect 7285 23137 7297 23140
rect 7331 23137 7343 23171
rect 8202 23168 8208 23180
rect 8163 23140 8208 23168
rect 7285 23131 7343 23137
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 11149 23171 11207 23177
rect 11149 23137 11161 23171
rect 11195 23168 11207 23171
rect 11238 23168 11244 23180
rect 11195 23140 11244 23168
rect 11195 23137 11207 23140
rect 11149 23131 11207 23137
rect 11238 23128 11244 23140
rect 11296 23128 11302 23180
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 4212 23072 5365 23100
rect 4212 23060 4218 23072
rect 5353 23069 5365 23072
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 8110 23060 8116 23112
rect 8168 23100 8174 23112
rect 8389 23103 8447 23109
rect 8389 23100 8401 23103
rect 8168 23072 8401 23100
rect 8168 23060 8174 23072
rect 8389 23069 8401 23072
rect 8435 23069 8447 23103
rect 8389 23063 8447 23069
rect 7834 22964 7840 22976
rect 7795 22936 7840 22964
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 8846 22924 8852 22976
rect 8904 22964 8910 22976
rect 9306 22964 9312 22976
rect 8904 22936 9312 22964
rect 8904 22924 8910 22936
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 10226 22964 10232 22976
rect 10187 22936 10232 22964
rect 10226 22924 10232 22936
rect 10284 22924 10290 22976
rect 10594 22924 10600 22976
rect 10652 22964 10658 22976
rect 12529 22967 12587 22973
rect 12529 22964 12541 22967
rect 10652 22936 12541 22964
rect 10652 22924 10658 22936
rect 12529 22933 12541 22936
rect 12575 22933 12587 22967
rect 12529 22927 12587 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 4985 22763 5043 22769
rect 4985 22729 4997 22763
rect 5031 22760 5043 22763
rect 5350 22760 5356 22772
rect 5031 22732 5356 22760
rect 5031 22729 5043 22732
rect 4985 22723 5043 22729
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 5592 22732 6837 22760
rect 5592 22720 5598 22732
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 6825 22723 6883 22729
rect 7190 22720 7196 22772
rect 7248 22760 7254 22772
rect 7466 22760 7472 22772
rect 7248 22732 7472 22760
rect 7248 22720 7254 22732
rect 7466 22720 7472 22732
rect 7524 22720 7530 22772
rect 8294 22760 8300 22772
rect 8255 22732 8300 22760
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 5368 22692 5396 22720
rect 5629 22695 5687 22701
rect 5629 22692 5641 22695
rect 5368 22664 5641 22692
rect 5629 22661 5641 22664
rect 5675 22692 5687 22695
rect 5718 22692 5724 22704
rect 5675 22664 5724 22692
rect 5675 22661 5687 22664
rect 5629 22655 5687 22661
rect 5718 22652 5724 22664
rect 5776 22692 5782 22704
rect 6181 22695 6239 22701
rect 6181 22692 6193 22695
rect 5776 22664 6193 22692
rect 5776 22652 5782 22664
rect 6181 22661 6193 22664
rect 6227 22692 6239 22695
rect 6227 22664 7420 22692
rect 6227 22661 6239 22664
rect 6181 22655 6239 22661
rect 2222 22624 2228 22636
rect 1412 22596 2228 22624
rect 1412 22565 1440 22596
rect 2222 22584 2228 22596
rect 2280 22584 2286 22636
rect 7392 22633 7420 22664
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22593 7435 22627
rect 7377 22587 7435 22593
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 10042 22624 10048 22636
rect 9815 22596 10048 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 10042 22584 10048 22596
rect 10100 22624 10106 22636
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 10100 22596 10425 22624
rect 10100 22584 10106 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 10413 22587 10471 22593
rect 11808 22596 13093 22624
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22525 1455 22559
rect 1397 22519 1455 22525
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22556 3663 22559
rect 3694 22556 3700 22568
rect 3651 22528 3700 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 3694 22516 3700 22528
rect 3752 22556 3758 22568
rect 4154 22556 4160 22568
rect 3752 22528 4160 22556
rect 3752 22516 3758 22528
rect 4154 22516 4160 22528
rect 4212 22516 4218 22568
rect 7193 22559 7251 22565
rect 7193 22525 7205 22559
rect 7239 22556 7251 22559
rect 7282 22556 7288 22568
rect 7239 22528 7288 22556
rect 7239 22525 7251 22528
rect 7193 22519 7251 22525
rect 7282 22516 7288 22528
rect 7340 22516 7346 22568
rect 10226 22556 10232 22568
rect 10187 22528 10232 22556
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 1670 22488 1676 22500
rect 1631 22460 1676 22488
rect 1670 22448 1676 22460
rect 1728 22448 1734 22500
rect 3850 22491 3908 22497
rect 3850 22488 3862 22491
rect 3436 22460 3862 22488
rect 3436 22432 3464 22460
rect 3850 22457 3862 22460
rect 3896 22457 3908 22491
rect 10321 22491 10379 22497
rect 10321 22488 10333 22491
rect 3850 22451 3908 22457
rect 9416 22460 10333 22488
rect 9416 22432 9444 22460
rect 10321 22457 10333 22460
rect 10367 22457 10379 22491
rect 10321 22451 10379 22457
rect 3418 22420 3424 22432
rect 3379 22392 3424 22420
rect 3418 22380 3424 22392
rect 3476 22380 3482 22432
rect 6641 22423 6699 22429
rect 6641 22389 6653 22423
rect 6687 22420 6699 22423
rect 7006 22420 7012 22432
rect 6687 22392 7012 22420
rect 6687 22389 6699 22392
rect 6641 22383 6699 22389
rect 7006 22380 7012 22392
rect 7064 22420 7070 22432
rect 7285 22423 7343 22429
rect 7285 22420 7297 22423
rect 7064 22392 7297 22420
rect 7064 22380 7070 22392
rect 7285 22389 7297 22392
rect 7331 22389 7343 22423
rect 7834 22420 7840 22432
rect 7795 22392 7840 22420
rect 7285 22383 7343 22389
rect 7834 22380 7840 22392
rect 7892 22420 7898 22432
rect 8110 22420 8116 22432
rect 7892 22392 8116 22420
rect 7892 22380 7898 22392
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 8662 22420 8668 22432
rect 8623 22392 8668 22420
rect 8662 22380 8668 22392
rect 8720 22380 8726 22432
rect 9398 22420 9404 22432
rect 9359 22392 9404 22420
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 9858 22420 9864 22432
rect 9819 22392 9864 22420
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 11241 22423 11299 22429
rect 11241 22389 11253 22423
rect 11287 22420 11299 22423
rect 11330 22420 11336 22432
rect 11287 22392 11336 22420
rect 11287 22389 11299 22392
rect 11241 22383 11299 22389
rect 11330 22380 11336 22392
rect 11388 22420 11394 22432
rect 11808 22429 11836 22596
rect 13081 22593 13093 22596
rect 13127 22624 13139 22627
rect 13354 22624 13360 22636
rect 13127 22596 13360 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 12158 22448 12164 22500
rect 12216 22488 12222 22500
rect 12253 22491 12311 22497
rect 12253 22488 12265 22491
rect 12216 22460 12265 22488
rect 12216 22448 12222 22460
rect 12253 22457 12265 22460
rect 12299 22488 12311 22491
rect 12897 22491 12955 22497
rect 12897 22488 12909 22491
rect 12299 22460 12909 22488
rect 12299 22457 12311 22460
rect 12253 22451 12311 22457
rect 12897 22457 12909 22460
rect 12943 22488 12955 22491
rect 13078 22488 13084 22500
rect 12943 22460 13084 22488
rect 12943 22457 12955 22460
rect 12897 22451 12955 22457
rect 13078 22448 13084 22460
rect 13136 22448 13142 22500
rect 11793 22423 11851 22429
rect 11793 22420 11805 22423
rect 11388 22392 11805 22420
rect 11388 22380 11394 22392
rect 11793 22389 11805 22392
rect 11839 22389 11851 22423
rect 11793 22383 11851 22389
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12437 22423 12495 22429
rect 12437 22420 12449 22423
rect 12032 22392 12449 22420
rect 12032 22380 12038 22392
rect 12437 22389 12449 22392
rect 12483 22389 12495 22423
rect 12802 22420 12808 22432
rect 12763 22392 12808 22420
rect 12437 22383 12495 22389
rect 12802 22380 12808 22392
rect 12860 22380 12866 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2406 22216 2412 22228
rect 2367 22188 2412 22216
rect 2406 22176 2412 22188
rect 2464 22176 2470 22228
rect 5074 22216 5080 22228
rect 5035 22188 5080 22216
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 6917 22219 6975 22225
rect 6917 22185 6929 22219
rect 6963 22216 6975 22219
rect 7282 22216 7288 22228
rect 6963 22188 7288 22216
rect 6963 22185 6975 22188
rect 6917 22179 6975 22185
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 8018 22216 8024 22228
rect 7979 22188 8024 22216
rect 8018 22176 8024 22188
rect 8076 22176 8082 22228
rect 9398 22176 9404 22228
rect 9456 22216 9462 22228
rect 9677 22219 9735 22225
rect 9677 22216 9689 22219
rect 9456 22188 9689 22216
rect 9456 22176 9462 22188
rect 9677 22185 9689 22188
rect 9723 22185 9735 22219
rect 9677 22179 9735 22185
rect 10226 22176 10232 22228
rect 10284 22216 10290 22228
rect 11241 22219 11299 22225
rect 11241 22216 11253 22219
rect 10284 22188 11253 22216
rect 10284 22176 10290 22188
rect 11241 22185 11253 22188
rect 11287 22185 11299 22219
rect 11241 22179 11299 22185
rect 11609 22219 11667 22225
rect 11609 22185 11621 22219
rect 11655 22216 11667 22219
rect 11974 22216 11980 22228
rect 11655 22188 11980 22216
rect 11655 22185 11667 22188
rect 11609 22179 11667 22185
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12986 22176 12992 22228
rect 13044 22216 13050 22228
rect 13173 22219 13231 22225
rect 13173 22216 13185 22219
rect 13044 22188 13185 22216
rect 13044 22176 13050 22188
rect 13173 22185 13185 22188
rect 13219 22185 13231 22219
rect 13173 22179 13231 22185
rect 3694 22148 3700 22160
rect 2608 22120 3700 22148
rect 2317 22083 2375 22089
rect 2317 22049 2329 22083
rect 2363 22080 2375 22083
rect 2498 22080 2504 22092
rect 2363 22052 2504 22080
rect 2363 22049 2375 22052
rect 2317 22043 2375 22049
rect 2498 22040 2504 22052
rect 2556 22080 2562 22092
rect 2608 22080 2636 22120
rect 3694 22108 3700 22120
rect 3752 22108 3758 22160
rect 5445 22151 5503 22157
rect 5445 22117 5457 22151
rect 5491 22148 5503 22151
rect 5534 22148 5540 22160
rect 5491 22120 5540 22148
rect 5491 22117 5503 22120
rect 5445 22111 5503 22117
rect 5534 22108 5540 22120
rect 5592 22108 5598 22160
rect 7006 22108 7012 22160
rect 7064 22148 7070 22160
rect 7558 22148 7564 22160
rect 7064 22120 7564 22148
rect 7064 22108 7070 22120
rect 7558 22108 7564 22120
rect 7616 22108 7622 22160
rect 10134 22108 10140 22160
rect 10192 22148 10198 22160
rect 11701 22151 11759 22157
rect 10192 22120 10272 22148
rect 10192 22108 10198 22120
rect 2556 22052 2636 22080
rect 2556 22040 2562 22052
rect 2682 22040 2688 22092
rect 2740 22080 2746 22092
rect 2777 22083 2835 22089
rect 2777 22080 2789 22083
rect 2740 22052 2789 22080
rect 2740 22040 2746 22052
rect 2777 22049 2789 22052
rect 2823 22049 2835 22083
rect 2777 22043 2835 22049
rect 3418 22040 3424 22092
rect 3476 22040 3482 22092
rect 6178 22080 6184 22092
rect 6139 22052 6184 22080
rect 6178 22040 6184 22052
rect 6236 22040 6242 22092
rect 7469 22083 7527 22089
rect 7469 22049 7481 22083
rect 7515 22080 7527 22083
rect 7929 22083 7987 22089
rect 7929 22080 7941 22083
rect 7515 22052 7941 22080
rect 7515 22049 7527 22052
rect 7469 22043 7527 22049
rect 7929 22049 7941 22052
rect 7975 22080 7987 22083
rect 8478 22080 8484 22092
rect 7975 22052 8484 22080
rect 7975 22049 7987 22052
rect 7929 22043 7987 22049
rect 8478 22040 8484 22052
rect 8536 22040 8542 22092
rect 9493 22083 9551 22089
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 10042 22080 10048 22092
rect 9539 22052 10048 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 2866 22012 2872 22024
rect 2827 21984 2872 22012
rect 2866 21972 2872 21984
rect 2924 21972 2930 22024
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 22012 3111 22015
rect 3234 22012 3240 22024
rect 3099 21984 3240 22012
rect 3099 21981 3111 21984
rect 3053 21975 3111 21981
rect 2406 21904 2412 21956
rect 2464 21944 2470 21956
rect 3068 21944 3096 21975
rect 3234 21972 3240 21984
rect 3292 22012 3298 22024
rect 3436 22012 3464 22040
rect 10244 22024 10272 22120
rect 11701 22117 11713 22151
rect 11747 22148 11759 22151
rect 11882 22148 11888 22160
rect 11747 22120 11888 22148
rect 11747 22117 11759 22120
rect 11701 22111 11759 22117
rect 11882 22108 11888 22120
rect 11940 22108 11946 22160
rect 12437 22151 12495 22157
rect 12437 22117 12449 22151
rect 12483 22148 12495 22151
rect 12802 22148 12808 22160
rect 12483 22120 12808 22148
rect 12483 22117 12495 22120
rect 12437 22111 12495 22117
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 10612 22052 11836 22080
rect 10612 22024 10640 22052
rect 3292 21984 3464 22012
rect 3292 21972 3298 21984
rect 5166 21972 5172 22024
rect 5224 22012 5230 22024
rect 5537 22015 5595 22021
rect 5537 22012 5549 22015
rect 5224 21984 5549 22012
rect 5224 21972 5230 21984
rect 5537 21981 5549 21984
rect 5583 21981 5595 22015
rect 5718 22012 5724 22024
rect 5679 21984 5724 22012
rect 5537 21975 5595 21981
rect 5718 21972 5724 21984
rect 5776 21972 5782 22024
rect 8110 22012 8116 22024
rect 8071 21984 8116 22012
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 10134 22012 10140 22024
rect 10095 21984 10140 22012
rect 10134 21972 10140 21984
rect 10192 21972 10198 22024
rect 10226 21972 10232 22024
rect 10284 21972 10290 22024
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10594 22012 10600 22024
rect 10367 21984 10600 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 10686 21972 10692 22024
rect 10744 22012 10750 22024
rect 10870 22012 10876 22024
rect 10744 21984 10876 22012
rect 10744 21972 10750 21984
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 11808 22021 11836 22052
rect 12618 22040 12624 22092
rect 12676 22080 12682 22092
rect 12894 22080 12900 22092
rect 12676 22052 12900 22080
rect 12676 22040 12682 22052
rect 12894 22040 12900 22052
rect 12952 22040 12958 22092
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 12250 21972 12256 22024
rect 12308 22012 12314 22024
rect 12434 22012 12440 22024
rect 12308 21984 12440 22012
rect 12308 21972 12314 21984
rect 12434 21972 12440 21984
rect 12492 22012 12498 22024
rect 13170 22012 13176 22024
rect 12492 21984 13176 22012
rect 12492 21972 12498 21984
rect 13170 21972 13176 21984
rect 13228 22012 13234 22024
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 13228 21984 13277 22012
rect 13228 21972 13234 21984
rect 13265 21981 13277 21984
rect 13311 21981 13323 22015
rect 13265 21975 13323 21981
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 13412 21984 13461 22012
rect 13412 21972 13418 21984
rect 13449 21981 13461 21984
rect 13495 22012 13507 22015
rect 13630 22012 13636 22024
rect 13495 21984 13636 22012
rect 13495 21981 13507 21984
rect 13449 21975 13507 21981
rect 13630 21972 13636 21984
rect 13688 21972 13694 22024
rect 2464 21916 3096 21944
rect 7561 21947 7619 21953
rect 2464 21904 2470 21916
rect 7561 21913 7573 21947
rect 7607 21944 7619 21947
rect 8202 21944 8208 21956
rect 7607 21916 8208 21944
rect 7607 21913 7619 21916
rect 7561 21907 7619 21913
rect 8202 21904 8208 21916
rect 8260 21944 8266 21956
rect 8573 21947 8631 21953
rect 8573 21944 8585 21947
rect 8260 21916 8585 21944
rect 8260 21904 8266 21916
rect 8573 21913 8585 21916
rect 8619 21913 8631 21947
rect 8573 21907 8631 21913
rect 11882 21904 11888 21956
rect 11940 21944 11946 21956
rect 12805 21947 12863 21953
rect 12805 21944 12817 21947
rect 11940 21916 12817 21944
rect 11940 21904 11946 21916
rect 12805 21913 12817 21916
rect 12851 21913 12863 21947
rect 12805 21907 12863 21913
rect 13078 21904 13084 21956
rect 13136 21944 13142 21956
rect 13136 21916 13400 21944
rect 13136 21904 13142 21916
rect 13372 21888 13400 21916
rect 1394 21836 1400 21888
rect 1452 21876 1458 21888
rect 9858 21876 9864 21888
rect 1452 21848 9864 21876
rect 1452 21836 1458 21848
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 10686 21876 10692 21888
rect 10647 21848 10692 21876
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 11149 21879 11207 21885
rect 11149 21845 11161 21879
rect 11195 21876 11207 21879
rect 11238 21876 11244 21888
rect 11195 21848 11244 21876
rect 11195 21845 11207 21848
rect 11149 21839 11207 21845
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 13354 21836 13360 21888
rect 13412 21836 13418 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 2406 21672 2412 21684
rect 2367 21644 2412 21672
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 3234 21632 3240 21684
rect 3292 21672 3298 21684
rect 3881 21675 3939 21681
rect 3881 21672 3893 21675
rect 3292 21644 3893 21672
rect 3292 21632 3298 21644
rect 3881 21641 3893 21644
rect 3927 21641 3939 21675
rect 3881 21635 3939 21641
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 5813 21675 5871 21681
rect 5813 21672 5825 21675
rect 5776 21644 5825 21672
rect 5776 21632 5782 21644
rect 5813 21641 5825 21644
rect 5859 21641 5871 21675
rect 7650 21672 7656 21684
rect 7563 21644 7656 21672
rect 5813 21635 5871 21641
rect 7650 21632 7656 21644
rect 7708 21672 7714 21684
rect 8110 21672 8116 21684
rect 7708 21644 8116 21672
rect 7708 21632 7714 21644
rect 8110 21632 8116 21644
rect 8168 21632 8174 21684
rect 8478 21672 8484 21684
rect 8439 21644 8484 21672
rect 8478 21632 8484 21644
rect 8536 21632 8542 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 10100 21644 10241 21672
rect 10100 21632 10106 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 11241 21675 11299 21681
rect 11241 21672 11253 21675
rect 10652 21644 11253 21672
rect 10652 21632 10658 21644
rect 11241 21641 11253 21644
rect 11287 21641 11299 21675
rect 11974 21672 11980 21684
rect 11935 21644 11980 21672
rect 11241 21635 11299 21641
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12342 21672 12348 21684
rect 12124 21644 12348 21672
rect 12124 21632 12130 21644
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 12986 21672 12992 21684
rect 12947 21644 12992 21672
rect 12986 21632 12992 21644
rect 13044 21632 13050 21684
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 13265 21675 13323 21681
rect 13265 21672 13277 21675
rect 13228 21644 13277 21672
rect 13228 21632 13234 21644
rect 13265 21641 13277 21644
rect 13311 21641 13323 21675
rect 13630 21672 13636 21684
rect 13591 21644 13636 21672
rect 13265 21635 13323 21641
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 7285 21607 7343 21613
rect 7285 21573 7297 21607
rect 7331 21604 7343 21607
rect 8018 21604 8024 21616
rect 7331 21576 8024 21604
rect 7331 21573 7343 21576
rect 7285 21567 7343 21573
rect 8018 21564 8024 21576
rect 8076 21564 8082 21616
rect 9950 21564 9956 21616
rect 10008 21604 10014 21616
rect 10612 21604 10640 21632
rect 10008 21576 10640 21604
rect 11701 21607 11759 21613
rect 10008 21564 10014 21576
rect 11701 21573 11713 21607
rect 11747 21604 11759 21607
rect 11882 21604 11888 21616
rect 11747 21576 11888 21604
rect 11747 21573 11759 21576
rect 11701 21567 11759 21573
rect 11882 21564 11888 21576
rect 11940 21564 11946 21616
rect 2498 21536 2504 21548
rect 2459 21508 2504 21536
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 7929 21539 7987 21545
rect 7929 21505 7941 21539
rect 7975 21536 7987 21539
rect 8386 21536 8392 21548
rect 7975 21508 8392 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 8386 21496 8392 21508
rect 8444 21536 8450 21548
rect 9033 21539 9091 21545
rect 9033 21536 9045 21539
rect 8444 21508 9045 21536
rect 8444 21496 8450 21508
rect 9033 21505 9045 21508
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 9769 21539 9827 21545
rect 9769 21505 9781 21539
rect 9815 21536 9827 21539
rect 10870 21536 10876 21548
rect 9815 21508 10876 21536
rect 9815 21505 9827 21508
rect 9769 21499 9827 21505
rect 10870 21496 10876 21508
rect 10928 21536 10934 21548
rect 11330 21536 11336 21548
rect 10928 21508 11336 21536
rect 10928 21496 10934 21508
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 12437 21539 12495 21545
rect 12437 21505 12449 21539
rect 12483 21536 12495 21539
rect 12802 21536 12808 21548
rect 12483 21508 12808 21536
rect 12483 21505 12495 21508
rect 12437 21499 12495 21505
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 8662 21428 8668 21480
rect 8720 21468 8726 21480
rect 8849 21471 8907 21477
rect 8849 21468 8861 21471
rect 8720 21440 8861 21468
rect 8720 21428 8726 21440
rect 8849 21437 8861 21440
rect 8895 21437 8907 21471
rect 8849 21431 8907 21437
rect 2041 21403 2099 21409
rect 2041 21369 2053 21403
rect 2087 21400 2099 21403
rect 2222 21400 2228 21412
rect 2087 21372 2228 21400
rect 2087 21369 2099 21372
rect 2041 21363 2099 21369
rect 2222 21360 2228 21372
rect 2280 21400 2286 21412
rect 2768 21403 2826 21409
rect 2768 21400 2780 21403
rect 2280 21372 2780 21400
rect 2280 21360 2286 21372
rect 2768 21369 2780 21372
rect 2814 21400 2826 21403
rect 3142 21400 3148 21412
rect 2814 21372 3148 21400
rect 2814 21369 2826 21372
rect 2768 21363 2826 21369
rect 3142 21360 3148 21372
rect 3200 21360 3206 21412
rect 10042 21360 10048 21412
rect 10100 21400 10106 21412
rect 10137 21403 10195 21409
rect 10137 21400 10149 21403
rect 10100 21372 10149 21400
rect 10100 21360 10106 21372
rect 10137 21369 10149 21372
rect 10183 21400 10195 21403
rect 10594 21400 10600 21412
rect 10183 21372 10600 21400
rect 10183 21369 10195 21372
rect 10137 21363 10195 21369
rect 10594 21360 10600 21372
rect 10652 21360 10658 21412
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 5166 21332 5172 21344
rect 5127 21304 5172 21332
rect 5166 21292 5172 21304
rect 5224 21292 5230 21344
rect 5534 21332 5540 21344
rect 5447 21304 5540 21332
rect 5534 21292 5540 21304
rect 5592 21332 5598 21344
rect 6086 21332 6092 21344
rect 5592 21304 6092 21332
rect 5592 21292 5598 21304
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 8389 21335 8447 21341
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8941 21335 8999 21341
rect 8941 21332 8953 21335
rect 8435 21304 8953 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8941 21301 8953 21304
rect 8987 21332 8999 21335
rect 9306 21332 9312 21344
rect 8987 21304 9312 21332
rect 8987 21301 8999 21304
rect 8941 21295 8999 21301
rect 9306 21292 9312 21304
rect 9364 21332 9370 21344
rect 9858 21332 9864 21344
rect 9364 21304 9864 21332
rect 9364 21292 9370 21304
rect 9858 21292 9864 21304
rect 9916 21292 9922 21344
rect 10686 21332 10692 21344
rect 10647 21304 10692 21332
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 1670 21088 1676 21140
rect 1728 21128 1734 21140
rect 2409 21131 2467 21137
rect 2409 21128 2421 21131
rect 1728 21100 2421 21128
rect 1728 21088 1734 21100
rect 2409 21097 2421 21100
rect 2455 21128 2467 21131
rect 2866 21128 2872 21140
rect 2455 21100 2872 21128
rect 2455 21097 2467 21100
rect 2409 21091 2467 21097
rect 2866 21088 2872 21100
rect 2924 21088 2930 21140
rect 8573 21131 8631 21137
rect 8573 21097 8585 21131
rect 8619 21128 8631 21131
rect 8662 21128 8668 21140
rect 8619 21100 8668 21128
rect 8619 21097 8631 21100
rect 8573 21091 8631 21097
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 10134 21128 10140 21140
rect 9539 21100 10140 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 10134 21088 10140 21100
rect 10192 21128 10198 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 10192 21100 10333 21128
rect 10192 21088 10198 21100
rect 10321 21097 10333 21100
rect 10367 21097 10379 21131
rect 10321 21091 10379 21097
rect 10686 21088 10692 21140
rect 10744 21128 10750 21140
rect 11885 21131 11943 21137
rect 11885 21128 11897 21131
rect 10744 21100 11897 21128
rect 10744 21088 10750 21100
rect 11885 21097 11897 21100
rect 11931 21097 11943 21131
rect 12342 21128 12348 21140
rect 12303 21100 12348 21128
rect 11885 21091 11943 21097
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 2777 21063 2835 21069
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 2958 21060 2964 21072
rect 2823 21032 2964 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 2958 21020 2964 21032
rect 3016 21020 3022 21072
rect 4433 21063 4491 21069
rect 4433 21029 4445 21063
rect 4479 21060 4491 21063
rect 4706 21060 4712 21072
rect 4479 21032 4712 21060
rect 4479 21029 4491 21032
rect 4433 21023 4491 21029
rect 4706 21020 4712 21032
rect 4764 21060 4770 21072
rect 5442 21060 5448 21072
rect 4764 21032 5448 21060
rect 4764 21020 4770 21032
rect 5442 21020 5448 21032
rect 5500 21020 5506 21072
rect 9950 21060 9956 21072
rect 9911 21032 9956 21060
rect 9950 21020 9956 21032
rect 10008 21020 10014 21072
rect 2869 20995 2927 21001
rect 2869 20961 2881 20995
rect 2915 20992 2927 20995
rect 3050 20992 3056 21004
rect 2915 20964 3056 20992
rect 2915 20961 2927 20964
rect 2869 20955 2927 20961
rect 3050 20952 3056 20964
rect 3108 20952 3114 21004
rect 4522 20992 4528 21004
rect 4483 20964 4528 20992
rect 4522 20952 4528 20964
rect 4580 20952 4586 21004
rect 6178 20952 6184 21004
rect 6236 20992 6242 21004
rect 6457 20995 6515 21001
rect 6457 20992 6469 20995
rect 6236 20964 6469 20992
rect 6236 20952 6242 20964
rect 6457 20961 6469 20964
rect 6503 20961 6515 20995
rect 6457 20955 6515 20961
rect 6546 20952 6552 21004
rect 6604 20992 6610 21004
rect 6713 20995 6771 21001
rect 6713 20992 6725 20995
rect 6604 20964 6725 20992
rect 6604 20952 6610 20964
rect 6713 20961 6725 20964
rect 6759 20992 6771 20995
rect 7834 20992 7840 21004
rect 6759 20964 7840 20992
rect 6759 20961 6771 20964
rect 6713 20955 6771 20961
rect 7834 20952 7840 20964
rect 7892 20952 7898 21004
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 10410 20992 10416 21004
rect 9824 20964 10416 20992
rect 9824 20952 9830 20964
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 10502 20952 10508 21004
rect 10560 20992 10566 21004
rect 10689 20995 10747 21001
rect 10689 20992 10701 20995
rect 10560 20964 10701 20992
rect 10560 20952 10566 20964
rect 10689 20961 10701 20964
rect 10735 20961 10747 20995
rect 10689 20955 10747 20961
rect 12066 20952 12072 21004
rect 12124 20992 12130 21004
rect 12253 20995 12311 21001
rect 12253 20992 12265 20995
rect 12124 20964 12265 20992
rect 12124 20952 12130 20964
rect 12253 20961 12265 20964
rect 12299 20961 12311 20995
rect 12253 20955 12311 20961
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20893 3019 20927
rect 4614 20924 4620 20936
rect 4575 20896 4620 20924
rect 2961 20887 3019 20893
rect 2976 20856 3004 20887
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 10778 20924 10784 20936
rect 10739 20896 10784 20924
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 10870 20884 10876 20936
rect 10928 20924 10934 20936
rect 12437 20927 12495 20933
rect 10928 20896 10973 20924
rect 10928 20884 10934 20896
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 3142 20856 3148 20868
rect 2976 20828 3148 20856
rect 3142 20816 3148 20828
rect 3200 20856 3206 20868
rect 4632 20856 4660 20884
rect 3200 20828 4660 20856
rect 3200 20816 3206 20828
rect 11606 20816 11612 20868
rect 11664 20856 11670 20868
rect 12452 20856 12480 20887
rect 11664 20828 12480 20856
rect 11664 20816 11670 20828
rect 2317 20791 2375 20797
rect 2317 20757 2329 20791
rect 2363 20788 2375 20791
rect 2682 20788 2688 20800
rect 2363 20760 2688 20788
rect 2363 20757 2375 20760
rect 2317 20751 2375 20757
rect 2682 20748 2688 20760
rect 2740 20788 2746 20800
rect 4065 20791 4123 20797
rect 4065 20788 4077 20791
rect 2740 20760 4077 20788
rect 2740 20748 2746 20760
rect 4065 20757 4077 20760
rect 4111 20757 4123 20791
rect 7834 20788 7840 20800
rect 7795 20760 7840 20788
rect 4065 20751 4123 20757
rect 7834 20748 7840 20760
rect 7892 20748 7898 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 1857 20587 1915 20593
rect 1857 20553 1869 20587
rect 1903 20584 1915 20587
rect 2958 20584 2964 20596
rect 1903 20556 2964 20584
rect 1903 20553 1915 20556
rect 1857 20547 1915 20553
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 4522 20544 4528 20596
rect 4580 20584 4586 20596
rect 4985 20587 5043 20593
rect 4985 20584 4997 20587
rect 4580 20556 4997 20584
rect 4580 20544 4586 20556
rect 4985 20553 4997 20556
rect 5031 20553 5043 20587
rect 4985 20547 5043 20553
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 5629 20587 5687 20593
rect 5629 20584 5641 20587
rect 5592 20556 5641 20584
rect 5592 20544 5598 20556
rect 5629 20553 5641 20556
rect 5675 20553 5687 20587
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 5629 20547 5687 20553
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 11606 20584 11612 20596
rect 11567 20556 11612 20584
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 12342 20584 12348 20596
rect 12023 20556 12348 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 2222 20516 2228 20528
rect 2183 20488 2228 20516
rect 2222 20476 2228 20488
rect 2280 20476 2286 20528
rect 4065 20519 4123 20525
rect 4065 20485 4077 20519
rect 4111 20516 4123 20519
rect 4614 20516 4620 20528
rect 4111 20488 4620 20516
rect 4111 20485 4123 20488
rect 4065 20479 4123 20485
rect 4614 20476 4620 20488
rect 4672 20476 4678 20528
rect 6178 20476 6184 20528
rect 6236 20516 6242 20528
rect 7009 20519 7067 20525
rect 7009 20516 7021 20519
rect 6236 20488 7021 20516
rect 6236 20476 6242 20488
rect 7009 20485 7021 20488
rect 7055 20485 7067 20519
rect 7009 20479 7067 20485
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2556 20420 2697 20448
rect 2556 20408 2562 20420
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 10091 20420 11161 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 11149 20417 11161 20420
rect 11195 20448 11207 20451
rect 11422 20448 11428 20460
rect 11195 20420 11428 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 11422 20408 11428 20420
rect 11480 20448 11486 20460
rect 11624 20448 11652 20544
rect 12066 20476 12072 20528
rect 12124 20516 12130 20528
rect 12621 20519 12679 20525
rect 12621 20516 12633 20519
rect 12124 20488 12633 20516
rect 12124 20476 12130 20488
rect 12621 20485 12633 20488
rect 12667 20485 12679 20519
rect 12621 20479 12679 20485
rect 11480 20420 11652 20448
rect 11480 20408 11486 20420
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8110 20380 8116 20392
rect 8067 20352 8116 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10060 20352 10885 20380
rect 10060 20324 10088 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 2593 20315 2651 20321
rect 2593 20281 2605 20315
rect 2639 20312 2651 20315
rect 2866 20312 2872 20324
rect 2639 20284 2872 20312
rect 2639 20281 2651 20284
rect 2593 20275 2651 20281
rect 2866 20272 2872 20284
rect 2924 20321 2930 20324
rect 2924 20315 2988 20321
rect 2924 20281 2942 20315
rect 2976 20281 2988 20315
rect 2924 20275 2988 20281
rect 7929 20315 7987 20321
rect 7929 20281 7941 20315
rect 7975 20312 7987 20315
rect 8266 20315 8324 20321
rect 8266 20312 8278 20315
rect 7975 20284 8278 20312
rect 7975 20281 7987 20284
rect 7929 20275 7987 20281
rect 8266 20281 8278 20284
rect 8312 20312 8324 20315
rect 8478 20312 8484 20324
rect 8312 20284 8484 20312
rect 8312 20281 8324 20284
rect 8266 20275 8324 20281
rect 2924 20272 2930 20275
rect 8478 20272 8484 20284
rect 8536 20272 8542 20324
rect 10042 20272 10048 20324
rect 10100 20272 10106 20324
rect 10965 20315 11023 20321
rect 10965 20312 10977 20315
rect 10336 20284 10977 20312
rect 4982 20204 4988 20256
rect 5040 20244 5046 20256
rect 5169 20247 5227 20253
rect 5169 20244 5181 20247
rect 5040 20216 5181 20244
rect 5040 20204 5046 20216
rect 5169 20213 5181 20216
rect 5215 20213 5227 20247
rect 9398 20244 9404 20256
rect 9359 20216 9404 20244
rect 5169 20207 5227 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 10134 20204 10140 20256
rect 10192 20244 10198 20256
rect 10336 20253 10364 20284
rect 10965 20281 10977 20284
rect 11011 20281 11023 20315
rect 10965 20275 11023 20281
rect 10321 20247 10379 20253
rect 10321 20244 10333 20247
rect 10192 20216 10333 20244
rect 10192 20204 10198 20216
rect 10321 20213 10333 20216
rect 10367 20213 10379 20247
rect 10502 20244 10508 20256
rect 10463 20216 10508 20244
rect 10321 20207 10379 20213
rect 10502 20204 10508 20216
rect 10560 20204 10566 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 2498 20000 2504 20052
rect 2556 20040 2562 20052
rect 3329 20043 3387 20049
rect 3329 20040 3341 20043
rect 2556 20012 3341 20040
rect 2556 20000 2562 20012
rect 3329 20009 3341 20012
rect 3375 20009 3387 20043
rect 4522 20040 4528 20052
rect 4483 20012 4528 20040
rect 3329 20003 3387 20009
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 4890 20040 4896 20052
rect 4851 20012 4896 20040
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 6236 20012 6377 20040
rect 6236 20000 6242 20012
rect 6365 20009 6377 20012
rect 6411 20009 6423 20043
rect 6365 20003 6423 20009
rect 7653 20043 7711 20049
rect 7653 20009 7665 20043
rect 7699 20040 7711 20043
rect 7834 20040 7840 20052
rect 7699 20012 7840 20040
rect 7699 20009 7711 20012
rect 7653 20003 7711 20009
rect 2866 19932 2872 19984
rect 2924 19972 2930 19984
rect 2961 19975 3019 19981
rect 2961 19972 2973 19975
rect 2924 19944 2973 19972
rect 2924 19932 2930 19944
rect 2961 19941 2973 19944
rect 3007 19972 3019 19975
rect 3510 19972 3516 19984
rect 3007 19944 3516 19972
rect 3007 19941 3019 19944
rect 2961 19935 3019 19941
rect 3510 19932 3516 19944
rect 3568 19972 3574 19984
rect 4341 19975 4399 19981
rect 4341 19972 4353 19975
rect 3568 19944 4353 19972
rect 3568 19932 3574 19944
rect 4341 19941 4353 19944
rect 4387 19941 4399 19975
rect 4341 19935 4399 19941
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 4356 19904 4384 19935
rect 6914 19904 6920 19916
rect 4356 19876 5120 19904
rect 6875 19876 6920 19904
rect 5092 19848 5120 19876
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 7009 19907 7067 19913
rect 7009 19873 7021 19907
rect 7055 19904 7067 19907
rect 7282 19904 7288 19916
rect 7055 19876 7288 19904
rect 7055 19873 7067 19876
rect 7009 19867 7067 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 4246 19796 4252 19848
rect 4304 19836 4310 19848
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 4304 19808 4997 19836
rect 4304 19796 4310 19808
rect 4985 19805 4997 19808
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 5074 19796 5080 19848
rect 5132 19836 5138 19848
rect 5132 19808 5225 19836
rect 5132 19796 5138 19808
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 7156 19808 7205 19836
rect 7156 19796 7162 19808
rect 7193 19805 7205 19808
rect 7239 19836 7251 19839
rect 7668 19836 7696 20003
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 10229 20043 10287 20049
rect 10229 20009 10241 20043
rect 10275 20040 10287 20043
rect 10410 20040 10416 20052
rect 10275 20012 10416 20040
rect 10275 20009 10287 20012
rect 10229 20003 10287 20009
rect 10410 20000 10416 20012
rect 10468 20040 10474 20052
rect 10778 20040 10784 20052
rect 10468 20012 10784 20040
rect 10468 20000 10474 20012
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 10965 20043 11023 20049
rect 10965 20040 10977 20043
rect 10928 20012 10977 20040
rect 10928 20000 10934 20012
rect 10965 20009 10977 20012
rect 11011 20040 11023 20043
rect 12529 20043 12587 20049
rect 12529 20040 12541 20043
rect 11011 20012 12541 20040
rect 11011 20009 11023 20012
rect 10965 20003 11023 20009
rect 12529 20009 12541 20012
rect 12575 20009 12587 20043
rect 12529 20003 12587 20009
rect 9493 19975 9551 19981
rect 9493 19941 9505 19975
rect 9539 19972 9551 19975
rect 10502 19972 10508 19984
rect 9539 19944 10508 19972
rect 9539 19941 9551 19944
rect 9493 19935 9551 19941
rect 10502 19932 10508 19944
rect 10560 19932 10566 19984
rect 11422 19981 11428 19984
rect 11416 19972 11428 19981
rect 11383 19944 11428 19972
rect 11416 19935 11428 19944
rect 11422 19932 11428 19935
rect 11480 19932 11486 19984
rect 11238 19864 11244 19916
rect 11296 19864 11302 19916
rect 7239 19808 7696 19836
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 10192 19808 10517 19836
rect 10192 19796 10198 19808
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 10870 19796 10876 19848
rect 10928 19836 10934 19848
rect 11149 19839 11207 19845
rect 11149 19836 11161 19839
rect 10928 19808 11161 19836
rect 10928 19796 10934 19808
rect 11149 19805 11161 19808
rect 11195 19836 11207 19839
rect 11256 19836 11284 19864
rect 11195 19808 11284 19836
rect 11195 19805 11207 19808
rect 11149 19799 11207 19805
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 6549 19771 6607 19777
rect 6549 19768 6561 19771
rect 5776 19740 6561 19768
rect 5776 19728 5782 19740
rect 6549 19737 6561 19740
rect 6595 19737 6607 19771
rect 6549 19731 6607 19737
rect 2501 19703 2559 19709
rect 2501 19669 2513 19703
rect 2547 19700 2559 19703
rect 2682 19700 2688 19712
rect 2547 19672 2688 19700
rect 2547 19669 2559 19672
rect 2501 19663 2559 19669
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 8110 19700 8116 19712
rect 8071 19672 8116 19700
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 1581 19499 1639 19505
rect 1581 19496 1593 19499
rect 1452 19468 1593 19496
rect 1452 19456 1458 19468
rect 1581 19465 1593 19468
rect 1627 19465 1639 19499
rect 2958 19496 2964 19508
rect 2919 19468 2964 19496
rect 1581 19459 1639 19465
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 10689 19499 10747 19505
rect 10689 19465 10701 19499
rect 10735 19496 10747 19499
rect 11054 19496 11060 19508
rect 10735 19468 11060 19496
rect 10735 19465 10747 19468
rect 10689 19459 10747 19465
rect 11054 19456 11060 19468
rect 11112 19496 11118 19508
rect 11333 19499 11391 19505
rect 11333 19496 11345 19499
rect 11112 19468 11345 19496
rect 11112 19456 11118 19468
rect 11333 19465 11345 19468
rect 11379 19496 11391 19499
rect 11422 19496 11428 19508
rect 11379 19468 11428 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 11422 19456 11428 19468
rect 11480 19456 11486 19508
rect 5442 19388 5448 19440
rect 5500 19388 5506 19440
rect 10870 19388 10876 19440
rect 10928 19428 10934 19440
rect 11609 19431 11667 19437
rect 11609 19428 11621 19431
rect 10928 19400 11621 19428
rect 10928 19388 10934 19400
rect 11609 19397 11621 19400
rect 11655 19397 11667 19431
rect 11609 19391 11667 19397
rect 3510 19360 3516 19372
rect 3471 19332 3516 19360
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 5074 19320 5080 19372
rect 5132 19360 5138 19372
rect 5169 19363 5227 19369
rect 5169 19360 5181 19363
rect 5132 19332 5181 19360
rect 5132 19320 5138 19332
rect 5169 19329 5181 19332
rect 5215 19360 5227 19363
rect 5460 19360 5488 19388
rect 5215 19332 5488 19360
rect 5215 19329 5227 19332
rect 5169 19323 5227 19329
rect 6178 19320 6184 19372
rect 6236 19360 6242 19372
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6236 19332 6837 19360
rect 6236 19320 6242 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 3050 19292 3056 19304
rect 2915 19264 3056 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 3050 19252 3056 19264
rect 3108 19292 3114 19304
rect 3326 19292 3332 19304
rect 3108 19264 3332 19292
rect 3108 19252 3114 19264
rect 3326 19252 3332 19264
rect 3384 19252 3390 19304
rect 4982 19292 4988 19304
rect 4943 19264 4988 19292
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 6546 19292 6552 19304
rect 6507 19264 6552 19292
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 7098 19301 7104 19304
rect 7092 19292 7104 19301
rect 7059 19264 7104 19292
rect 7092 19255 7104 19264
rect 7098 19252 7104 19255
rect 7156 19252 7162 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9272 19264 9321 19292
rect 9272 19252 9278 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 4525 19227 4583 19233
rect 4525 19193 4537 19227
rect 4571 19224 4583 19227
rect 4890 19224 4896 19236
rect 4571 19196 4896 19224
rect 4571 19193 4583 19196
rect 4525 19187 4583 19193
rect 4890 19184 4896 19196
rect 4948 19184 4954 19236
rect 6086 19184 6092 19236
rect 6144 19224 6150 19236
rect 6273 19227 6331 19233
rect 6273 19224 6285 19227
rect 6144 19196 6285 19224
rect 6144 19184 6150 19196
rect 6273 19193 6285 19196
rect 6319 19224 6331 19227
rect 6822 19224 6828 19236
rect 6319 19196 6828 19224
rect 6319 19193 6331 19196
rect 6273 19187 6331 19193
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 9398 19224 9404 19236
rect 9140 19196 9404 19224
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3384 19128 3433 19156
rect 3384 19116 3390 19128
rect 3421 19125 3433 19128
rect 3467 19125 3479 19159
rect 3421 19119 3479 19125
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4246 19156 4252 19168
rect 4203 19128 4252 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 4617 19159 4675 19165
rect 4617 19125 4629 19159
rect 4663 19156 4675 19159
rect 4706 19156 4712 19168
rect 4663 19128 4712 19156
rect 4663 19125 4675 19128
rect 4617 19119 4675 19125
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5074 19156 5080 19168
rect 5035 19128 5080 19156
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 5629 19159 5687 19165
rect 5629 19156 5641 19159
rect 5592 19128 5641 19156
rect 5592 19116 5598 19128
rect 5629 19125 5641 19128
rect 5675 19125 5687 19159
rect 8202 19156 8208 19168
rect 8163 19128 8208 19156
rect 5629 19119 5687 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 9140 19165 9168 19196
rect 9398 19184 9404 19196
rect 9456 19224 9462 19236
rect 9554 19227 9612 19233
rect 9554 19224 9566 19227
rect 9456 19196 9566 19224
rect 9456 19184 9462 19196
rect 9554 19193 9566 19196
rect 9600 19193 9612 19227
rect 9554 19187 9612 19193
rect 9125 19159 9183 19165
rect 9125 19156 9137 19159
rect 8444 19128 9137 19156
rect 8444 19116 8450 19128
rect 9125 19125 9137 19128
rect 9171 19125 9183 19159
rect 9125 19119 9183 19125
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 4982 18952 4988 18964
rect 4943 18924 4988 18952
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 5718 18952 5724 18964
rect 5679 18924 5724 18952
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 6641 18955 6699 18961
rect 6641 18921 6653 18955
rect 6687 18952 6699 18955
rect 7098 18952 7104 18964
rect 6687 18924 7104 18952
rect 6687 18921 6699 18924
rect 6641 18915 6699 18921
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 9214 18912 9220 18964
rect 9272 18952 9278 18964
rect 9309 18955 9367 18961
rect 9309 18952 9321 18955
rect 9272 18924 9321 18952
rect 9272 18912 9278 18924
rect 9309 18921 9321 18924
rect 9355 18921 9367 18955
rect 10410 18952 10416 18964
rect 10371 18924 10416 18952
rect 9309 18915 9367 18921
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 10873 18955 10931 18961
rect 10873 18952 10885 18955
rect 10744 18924 10885 18952
rect 10744 18912 10750 18924
rect 10873 18921 10885 18924
rect 10919 18921 10931 18955
rect 10873 18915 10931 18921
rect 4709 18887 4767 18893
rect 4709 18853 4721 18887
rect 4755 18884 4767 18887
rect 5074 18884 5080 18896
rect 4755 18856 5080 18884
rect 4755 18853 4767 18856
rect 4709 18847 4767 18853
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 5534 18776 5540 18828
rect 5592 18816 5598 18828
rect 5629 18819 5687 18825
rect 5629 18816 5641 18819
rect 5592 18788 5641 18816
rect 5592 18776 5598 18788
rect 5629 18785 5641 18788
rect 5675 18785 5687 18819
rect 5629 18779 5687 18785
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6144 18788 6837 18816
rect 6144 18776 6150 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 10870 18816 10876 18828
rect 10827 18788 10876 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 4706 18708 4712 18760
rect 4764 18748 4770 18760
rect 5905 18751 5963 18757
rect 5905 18748 5917 18751
rect 4764 18720 5917 18748
rect 4764 18708 4770 18720
rect 5905 18717 5917 18720
rect 5951 18748 5963 18751
rect 7282 18748 7288 18760
rect 5951 18720 7288 18748
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 11054 18748 11060 18760
rect 11015 18720 11060 18748
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 3053 18615 3111 18621
rect 3053 18581 3065 18615
rect 3099 18612 3111 18615
rect 3326 18612 3332 18624
rect 3099 18584 3332 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 5258 18612 5264 18624
rect 5219 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 7834 18572 7840 18624
rect 7892 18612 7898 18624
rect 8113 18615 8171 18621
rect 8113 18612 8125 18615
rect 7892 18584 8125 18612
rect 7892 18572 7898 18584
rect 8113 18581 8125 18584
rect 8159 18581 8171 18615
rect 8113 18575 8171 18581
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3053 18411 3111 18417
rect 3053 18408 3065 18411
rect 2832 18380 3065 18408
rect 2832 18368 2838 18380
rect 3053 18377 3065 18380
rect 3099 18377 3111 18411
rect 4706 18408 4712 18420
rect 4667 18380 4712 18408
rect 3053 18371 3111 18377
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 4982 18368 4988 18420
rect 5040 18408 5046 18420
rect 5994 18408 6000 18420
rect 5040 18380 6000 18408
rect 5040 18368 5046 18380
rect 5994 18368 6000 18380
rect 6052 18408 6058 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6052 18380 6561 18408
rect 6052 18368 6058 18380
rect 6549 18377 6561 18380
rect 6595 18408 6607 18411
rect 10505 18411 10563 18417
rect 6595 18380 7236 18408
rect 6595 18377 6607 18380
rect 6549 18371 6607 18377
rect 5077 18343 5135 18349
rect 5077 18309 5089 18343
rect 5123 18340 5135 18343
rect 5534 18340 5540 18352
rect 5123 18312 5540 18340
rect 5123 18309 5135 18312
rect 5077 18303 5135 18309
rect 5534 18300 5540 18312
rect 5592 18340 5598 18352
rect 6822 18340 6828 18352
rect 5592 18312 6828 18340
rect 5592 18300 5598 18312
rect 6822 18300 6828 18312
rect 6880 18300 6886 18352
rect 3142 18232 3148 18284
rect 3200 18272 3206 18284
rect 3510 18272 3516 18284
rect 3200 18244 3516 18272
rect 3200 18232 3206 18244
rect 3510 18232 3516 18244
rect 3568 18272 3574 18284
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 3568 18244 3617 18272
rect 3568 18232 3574 18244
rect 3605 18241 3617 18244
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5316 18244 5641 18272
rect 5316 18232 5322 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3007 18176 3433 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 3421 18173 3433 18176
rect 3467 18204 3479 18207
rect 3694 18204 3700 18216
rect 3467 18176 3700 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 3694 18164 3700 18176
rect 3752 18164 3758 18216
rect 5736 18204 5764 18235
rect 7208 18213 7236 18380
rect 10505 18377 10517 18411
rect 10551 18408 10563 18411
rect 10686 18408 10692 18420
rect 10551 18380 10692 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 11149 18411 11207 18417
rect 11149 18408 11161 18411
rect 11112 18380 11161 18408
rect 11112 18368 11118 18380
rect 11149 18377 11161 18380
rect 11195 18377 11207 18411
rect 11149 18371 11207 18377
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 7340 18244 7481 18272
rect 7340 18232 7346 18244
rect 7469 18241 7481 18244
rect 7515 18272 7527 18275
rect 8202 18272 8208 18284
rect 7515 18244 8208 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 4540 18176 5764 18204
rect 7193 18207 7251 18213
rect 2593 18139 2651 18145
rect 2593 18105 2605 18139
rect 2639 18136 2651 18139
rect 2639 18108 3556 18136
rect 2639 18105 2651 18108
rect 2593 18099 2651 18105
rect 3528 18080 3556 18108
rect 4540 18080 4568 18176
rect 7193 18173 7205 18207
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 5537 18139 5595 18145
rect 5537 18105 5549 18139
rect 5583 18136 5595 18139
rect 5626 18136 5632 18148
rect 5583 18108 5632 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 5626 18096 5632 18108
rect 5684 18136 5690 18148
rect 5684 18108 6868 18136
rect 5684 18096 5690 18108
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 4341 18071 4399 18077
rect 4341 18037 4353 18071
rect 4387 18068 4399 18071
rect 4522 18068 4528 18080
rect 4387 18040 4528 18068
rect 4387 18037 4399 18040
rect 4341 18031 4399 18037
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 6086 18028 6092 18080
rect 6144 18068 6150 18080
rect 6840 18077 6868 18108
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 6144 18040 6193 18068
rect 6144 18028 6150 18040
rect 6181 18037 6193 18040
rect 6227 18037 6239 18071
rect 6181 18031 6239 18037
rect 6825 18071 6883 18077
rect 6825 18037 6837 18071
rect 6871 18037 6883 18071
rect 6825 18031 6883 18037
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 7156 18040 7297 18068
rect 7156 18028 7162 18040
rect 7285 18037 7297 18040
rect 7331 18068 7343 18071
rect 8018 18068 8024 18080
rect 7331 18040 8024 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 8113 18071 8171 18077
rect 8113 18037 8125 18071
rect 8159 18068 8171 18071
rect 8294 18068 8300 18080
rect 8159 18040 8300 18068
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9306 18068 9312 18080
rect 9171 18040 9312 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 10870 18068 10876 18080
rect 10831 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 3142 17864 3148 17876
rect 3103 17836 3148 17864
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 5442 17864 5448 17876
rect 5403 17836 5448 17864
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 5718 17824 5724 17876
rect 5776 17864 5782 17876
rect 5997 17867 6055 17873
rect 5997 17864 6009 17867
rect 5776 17836 6009 17864
rect 5776 17824 5782 17836
rect 5997 17833 6009 17836
rect 6043 17833 6055 17867
rect 7282 17864 7288 17876
rect 7243 17836 7288 17864
rect 5997 17827 6055 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 7975 17836 8493 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 8481 17833 8493 17836
rect 8527 17864 8539 17867
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 8527 17836 9689 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 9677 17827 9735 17833
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 8389 17799 8447 17805
rect 8389 17796 8401 17799
rect 8352 17768 8401 17796
rect 8352 17756 8358 17768
rect 8389 17765 8401 17768
rect 8435 17765 8447 17799
rect 8389 17759 8447 17765
rect 10226 17756 10232 17808
rect 10284 17756 10290 17808
rect 4338 17737 4344 17740
rect 3789 17731 3847 17737
rect 3789 17697 3801 17731
rect 3835 17728 3847 17731
rect 4332 17728 4344 17737
rect 3835 17700 4344 17728
rect 3835 17697 3847 17700
rect 3789 17691 3847 17697
rect 4332 17691 4344 17700
rect 4338 17688 4344 17691
rect 4396 17688 4402 17740
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9732 17700 10057 17728
rect 9732 17688 9738 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10244 17728 10272 17756
rect 10410 17728 10416 17740
rect 10183 17700 10416 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 3234 17620 3240 17672
rect 3292 17660 3298 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3292 17632 4077 17660
rect 3292 17620 3298 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 8536 17632 8585 17660
rect 8536 17620 8542 17632
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 10008 17632 10241 17660
rect 10008 17620 10014 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 6917 17527 6975 17533
rect 6917 17493 6929 17527
rect 6963 17524 6975 17527
rect 7098 17524 7104 17536
rect 6963 17496 7104 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7800 17496 8033 17524
rect 7800 17484 7806 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 3568 17292 3709 17320
rect 3568 17280 3574 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 5258 17320 5264 17332
rect 5219 17292 5264 17320
rect 3697 17283 3755 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5626 17320 5632 17332
rect 5587 17292 5632 17320
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 8941 17323 8999 17329
rect 8941 17320 8953 17323
rect 8352 17292 8953 17320
rect 8352 17280 8358 17292
rect 8941 17289 8953 17292
rect 8987 17289 8999 17323
rect 8941 17283 8999 17289
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 9732 17292 9965 17320
rect 9732 17280 9738 17292
rect 9953 17289 9965 17292
rect 9999 17320 10011 17323
rect 10502 17320 10508 17332
rect 9999 17292 10508 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 11974 17252 11980 17264
rect 11204 17224 11980 17252
rect 11204 17212 11210 17224
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 3970 17184 3976 17196
rect 3651 17156 3976 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 3970 17144 3976 17156
rect 4028 17184 4034 17196
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 4028 17156 4169 17184
rect 4028 17144 4034 17156
rect 4157 17153 4169 17156
rect 4203 17153 4215 17187
rect 4338 17184 4344 17196
rect 4251 17156 4344 17184
rect 4157 17147 4215 17153
rect 4338 17144 4344 17156
rect 4396 17184 4402 17196
rect 7285 17187 7343 17193
rect 4396 17156 4844 17184
rect 4396 17144 4402 17156
rect 3970 17008 3976 17060
rect 4028 17048 4034 17060
rect 4065 17051 4123 17057
rect 4065 17048 4077 17051
rect 4028 17020 4077 17048
rect 4028 17008 4034 17020
rect 4065 17017 4077 17020
rect 4111 17017 4123 17051
rect 4065 17011 4123 17017
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 4816 16989 4844 17156
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7331 17156 7941 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7929 17153 7941 17156
rect 7975 17184 7987 17187
rect 8386 17184 8392 17196
rect 7975 17156 8392 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8527 17156 9597 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 9585 17153 9597 17156
rect 9631 17184 9643 17187
rect 9950 17184 9956 17196
rect 9631 17156 9956 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 8496 17116 8524 17147
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 9306 17116 9312 17128
rect 8352 17088 8524 17116
rect 9267 17088 9312 17116
rect 8352 17076 8358 17088
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 7558 17048 7564 17060
rect 6687 17020 7564 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7558 17008 7564 17020
rect 7616 17048 7622 17060
rect 7837 17051 7895 17057
rect 7837 17048 7849 17051
rect 7616 17020 7849 17048
rect 7616 17008 7622 17020
rect 7837 17017 7849 17020
rect 7883 17017 7895 17051
rect 7837 17011 7895 17017
rect 4801 16983 4859 16989
rect 4801 16949 4813 16983
rect 4847 16980 4859 16983
rect 5442 16980 5448 16992
rect 4847 16952 5448 16980
rect 4847 16949 4859 16952
rect 4801 16943 4859 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 8849 16983 8907 16989
rect 8849 16949 8861 16983
rect 8895 16980 8907 16983
rect 9398 16980 9404 16992
rect 8895 16952 9404 16980
rect 8895 16949 8907 16952
rect 8849 16943 8907 16949
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10410 16980 10416 16992
rect 10371 16952 10416 16980
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 3789 16779 3847 16785
rect 3789 16745 3801 16779
rect 3835 16776 3847 16779
rect 3970 16776 3976 16788
rect 3835 16748 3976 16776
rect 3835 16745 3847 16748
rect 3789 16739 3847 16745
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 5166 16776 5172 16788
rect 5127 16748 5172 16776
rect 5166 16736 5172 16748
rect 5224 16776 5230 16788
rect 5534 16776 5540 16788
rect 5224 16748 5540 16776
rect 5224 16736 5230 16748
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 7558 16776 7564 16788
rect 7519 16748 7564 16776
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8573 16779 8631 16785
rect 8573 16776 8585 16779
rect 8536 16748 8585 16776
rect 8536 16736 8542 16748
rect 8573 16745 8585 16748
rect 8619 16745 8631 16779
rect 8573 16739 8631 16745
rect 9033 16779 9091 16785
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9306 16776 9312 16788
rect 9079 16748 9312 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 1670 16708 1676 16720
rect 1631 16680 1676 16708
rect 1670 16668 1676 16680
rect 1728 16668 1734 16720
rect 2866 16668 2872 16720
rect 2924 16708 2930 16720
rect 2961 16711 3019 16717
rect 2961 16708 2973 16711
rect 2924 16680 2973 16708
rect 2924 16668 2930 16680
rect 2961 16677 2973 16680
rect 3007 16677 3019 16711
rect 2961 16671 3019 16677
rect 7101 16711 7159 16717
rect 7101 16677 7113 16711
rect 7147 16708 7159 16711
rect 7742 16708 7748 16720
rect 7147 16680 7748 16708
rect 7147 16677 7159 16680
rect 7101 16671 7159 16677
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 2674 16643 2732 16649
rect 2674 16640 2686 16643
rect 2608 16612 2686 16640
rect 2608 16504 2636 16612
rect 2674 16609 2686 16612
rect 2720 16609 2732 16643
rect 5074 16640 5080 16652
rect 5035 16612 5080 16640
rect 2674 16603 2732 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16640 6791 16643
rect 6822 16640 6828 16652
rect 6779 16612 6828 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7469 16643 7527 16649
rect 7469 16609 7481 16643
rect 7515 16640 7527 16643
rect 7926 16640 7932 16652
rect 7515 16612 7788 16640
rect 7887 16612 7932 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 5258 16572 5264 16584
rect 5219 16544 5264 16572
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 7760 16572 7788 16612
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8018 16600 8024 16652
rect 8076 16640 8082 16652
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 8076 16612 8121 16640
rect 9600 16612 10241 16640
rect 8076 16600 8082 16612
rect 8036 16572 8064 16600
rect 9600 16584 9628 16612
rect 10229 16609 10241 16612
rect 10275 16640 10287 16643
rect 11054 16640 11060 16652
rect 10275 16612 11060 16640
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11324 16643 11382 16649
rect 11324 16609 11336 16643
rect 11370 16640 11382 16643
rect 11606 16640 11612 16652
rect 11370 16612 11612 16640
rect 11370 16609 11382 16612
rect 11324 16603 11382 16609
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 7760 16544 8064 16572
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16572 8263 16575
rect 8478 16572 8484 16584
rect 8251 16544 8484 16572
rect 8251 16541 8263 16544
rect 8205 16535 8263 16541
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 9582 16532 9588 16584
rect 9640 16532 9646 16584
rect 2774 16504 2780 16516
rect 2608 16476 2780 16504
rect 2774 16464 2780 16476
rect 2832 16504 2838 16516
rect 4709 16507 4767 16513
rect 4709 16504 4721 16507
rect 2832 16476 4721 16504
rect 2832 16464 2838 16476
rect 4709 16473 4721 16476
rect 4755 16473 4767 16507
rect 9950 16504 9956 16516
rect 9863 16476 9956 16504
rect 4709 16467 4767 16473
rect 9950 16464 9956 16476
rect 10008 16504 10014 16516
rect 10318 16504 10324 16516
rect 10008 16476 10324 16504
rect 10008 16464 10014 16476
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 4341 16439 4399 16445
rect 4341 16405 4353 16439
rect 4387 16436 4399 16439
rect 4522 16436 4528 16448
rect 4387 16408 4528 16436
rect 4387 16405 4399 16408
rect 4341 16399 4399 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 12492 16408 12537 16436
rect 12492 16396 12498 16408
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 1394 16192 1400 16244
rect 1452 16232 1458 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1452 16204 1593 16232
rect 1452 16192 1458 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 2774 16232 2780 16244
rect 2735 16204 2780 16232
rect 1581 16195 1639 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5592 16204 6193 16232
rect 5592 16192 5598 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 8478 16232 8484 16244
rect 8439 16204 8484 16232
rect 6181 16195 6239 16201
rect 8478 16192 8484 16204
rect 8536 16232 8542 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8536 16204 9045 16232
rect 8536 16192 8542 16204
rect 9033 16201 9045 16204
rect 9079 16201 9091 16235
rect 9033 16195 9091 16201
rect 9306 16192 9312 16244
rect 9364 16232 9370 16244
rect 9490 16232 9496 16244
rect 9364 16204 9496 16232
rect 9364 16192 9370 16204
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 11146 16232 11152 16244
rect 10744 16204 11152 16232
rect 10744 16192 10750 16204
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16096 9551 16099
rect 9539 16068 9720 16096
rect 9539 16065 9551 16068
rect 9493 16059 9551 16065
rect 3234 15988 3240 16040
rect 3292 16028 3298 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3292 16000 3433 16028
rect 3292 15988 3298 16000
rect 3421 15997 3433 16000
rect 3467 16028 3479 16031
rect 3970 16028 3976 16040
rect 3467 16000 3976 16028
rect 3467 15997 3479 16000
rect 3421 15991 3479 15997
rect 3970 15988 3976 16000
rect 4028 16028 4034 16040
rect 4249 16031 4307 16037
rect 4249 16028 4261 16031
rect 4028 16000 4261 16028
rect 4028 15988 4034 16000
rect 4249 15997 4261 16000
rect 4295 15997 4307 16031
rect 4249 15991 4307 15997
rect 6822 15988 6828 16040
rect 6880 16028 6886 16040
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 6880 16000 7113 16028
rect 6880 15988 6886 16000
rect 7101 15997 7113 16000
rect 7147 16028 7159 16031
rect 8754 16028 8760 16040
rect 7147 16000 8760 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 8754 15988 8760 16000
rect 8812 16028 8818 16040
rect 9582 16028 9588 16040
rect 8812 16000 9588 16028
rect 8812 15988 8818 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9692 16028 9720 16068
rect 9858 16037 9864 16040
rect 9852 16028 9864 16037
rect 9692 16000 9864 16028
rect 9852 15991 9864 16000
rect 9858 15988 9864 15991
rect 9916 15988 9922 16040
rect 4522 15969 4528 15972
rect 4516 15960 4528 15969
rect 4483 15932 4528 15960
rect 4516 15923 4528 15932
rect 4522 15920 4528 15923
rect 4580 15920 4586 15972
rect 7374 15969 7380 15972
rect 7368 15960 7380 15969
rect 7335 15932 7380 15960
rect 7368 15923 7380 15932
rect 7374 15920 7380 15923
rect 7432 15920 7438 15972
rect 11606 15960 11612 15972
rect 11519 15932 11612 15960
rect 11606 15920 11612 15932
rect 11664 15960 11670 15972
rect 12250 15960 12256 15972
rect 11664 15932 12256 15960
rect 11664 15920 11670 15932
rect 12250 15920 12256 15932
rect 12308 15920 12314 15972
rect 3786 15892 3792 15904
rect 3747 15864 3792 15892
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 4154 15892 4160 15904
rect 4115 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15892 4218 15904
rect 5258 15892 5264 15904
rect 4212 15864 5264 15892
rect 4212 15852 4218 15864
rect 5258 15852 5264 15864
rect 5316 15892 5322 15904
rect 5629 15895 5687 15901
rect 5629 15892 5641 15895
rect 5316 15864 5641 15892
rect 5316 15852 5322 15864
rect 5629 15861 5641 15864
rect 5675 15861 5687 15895
rect 5629 15855 5687 15861
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7926 15892 7932 15904
rect 6687 15864 7932 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 9548 15864 10977 15892
rect 9548 15852 9554 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11112 15864 11897 15892
rect 11112 15852 11118 15864
rect 11885 15861 11897 15864
rect 11931 15861 11943 15895
rect 11885 15855 11943 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7340 15660 7573 15688
rect 7340 15648 7346 15660
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 7561 15651 7619 15657
rect 7653 15691 7711 15697
rect 7653 15657 7665 15691
rect 7699 15688 7711 15691
rect 7926 15688 7932 15700
rect 7699 15660 7932 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8294 15688 8300 15700
rect 8159 15660 8300 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8294 15648 8300 15660
rect 8352 15688 8358 15700
rect 8662 15688 8668 15700
rect 8352 15660 8668 15688
rect 8352 15648 8358 15660
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10042 15648 10048 15700
rect 10100 15648 10106 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11425 15691 11483 15697
rect 11425 15688 11437 15691
rect 11112 15660 11437 15688
rect 11112 15648 11118 15660
rect 11425 15657 11437 15660
rect 11471 15657 11483 15691
rect 11425 15651 11483 15657
rect 7466 15580 7472 15632
rect 7524 15620 7530 15632
rect 8021 15623 8079 15629
rect 8021 15620 8033 15623
rect 7524 15592 8033 15620
rect 7524 15580 7530 15592
rect 8021 15589 8033 15592
rect 8067 15589 8079 15623
rect 8021 15583 8079 15589
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 4321 15555 4379 15561
rect 4321 15552 4333 15555
rect 4212 15524 4333 15552
rect 4212 15512 4218 15524
rect 4321 15521 4333 15524
rect 4367 15521 4379 15555
rect 4321 15515 4379 15521
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15552 7251 15555
rect 7374 15552 7380 15564
rect 7239 15524 7380 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7374 15512 7380 15524
rect 7432 15552 7438 15564
rect 7432 15524 8248 15552
rect 7432 15512 7438 15524
rect 8220 15496 8248 15524
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10060 15561 10088 15648
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9732 15524 10057 15552
rect 9732 15512 9738 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 4028 15456 4077 15484
rect 4028 15444 4034 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 6546 15484 6552 15496
rect 6507 15456 6552 15484
rect 4065 15447 4123 15453
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8260 15456 8305 15484
rect 8260 15444 8266 15456
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9640 15456 10149 15484
rect 9640 15444 9646 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10137 15447 10195 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 11440 15484 11468 15651
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11865 15555 11923 15561
rect 11865 15552 11877 15555
rect 11572 15524 11877 15552
rect 11572 15512 11578 15524
rect 11865 15521 11877 15524
rect 11911 15521 11923 15555
rect 11865 15515 11923 15521
rect 11609 15487 11667 15493
rect 11609 15484 11621 15487
rect 11440 15456 11621 15484
rect 11609 15453 11621 15456
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 8754 15308 8760 15360
rect 8812 15348 8818 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8812 15320 9137 15348
rect 8812 15308 8818 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9125 15311 9183 15317
rect 12250 15308 12256 15360
rect 12308 15348 12314 15360
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12308 15320 13001 15348
rect 12308 15308 12314 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 4154 15144 4160 15156
rect 4115 15116 4160 15144
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 5074 15104 5080 15156
rect 5132 15144 5138 15156
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 5132 15116 5181 15144
rect 5132 15104 5138 15116
rect 5169 15113 5181 15116
rect 5215 15113 5227 15147
rect 5169 15107 5227 15113
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 7650 15144 7656 15156
rect 7524 15116 7656 15144
rect 7524 15104 7530 15116
rect 7650 15104 7656 15116
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 7837 15107 7895 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 10376 15116 10517 15144
rect 10376 15104 10382 15116
rect 10505 15113 10517 15116
rect 10551 15144 10563 15147
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 10551 15116 11069 15144
rect 10551 15113 10563 15116
rect 10505 15107 10563 15113
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11514 15144 11520 15156
rect 11475 15116 11520 15144
rect 11057 15107 11115 15113
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 12158 15144 12164 15156
rect 12119 15116 12164 15144
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 5920 15048 6837 15076
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4580 14980 5089 15008
rect 4580 14968 4586 14980
rect 5077 14977 5089 14980
rect 5123 15008 5135 15011
rect 5810 15008 5816 15020
rect 5123 14980 5816 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14940 4767 14943
rect 5537 14943 5595 14949
rect 5537 14940 5549 14943
rect 4755 14912 5549 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 5537 14909 5549 14912
rect 5583 14940 5595 14943
rect 5920 14940 5948 15048
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 6825 15039 6883 15045
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 13078 15076 13084 15088
rect 12952 15048 13084 15076
rect 12952 15036 12958 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7340 14980 7389 15008
rect 7340 14968 7346 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12768 14980 13001 15008
rect 12768 14968 12774 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 5583 14912 5948 14940
rect 6273 14943 6331 14949
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 6273 14909 6285 14943
rect 6319 14940 6331 14943
rect 6546 14940 6552 14952
rect 6319 14912 6552 14940
rect 6319 14909 6331 14912
rect 6273 14903 6331 14909
rect 6546 14900 6552 14912
rect 6604 14940 6610 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6604 14912 7205 14940
rect 6604 14900 6610 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 8754 14940 8760 14952
rect 8352 14912 8760 14940
rect 8352 14900 8358 14912
rect 8754 14900 8760 14912
rect 8812 14940 8818 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8812 14912 9137 14940
rect 8812 14900 8818 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 12158 14900 12164 14952
rect 12216 14940 12222 14952
rect 12216 14912 12940 14940
rect 12216 14900 12222 14912
rect 9030 14872 9036 14884
rect 8943 14844 9036 14872
rect 9030 14832 9036 14844
rect 9088 14872 9094 14884
rect 9392 14875 9450 14881
rect 9392 14872 9404 14875
rect 9088 14844 9404 14872
rect 9088 14832 9094 14844
rect 9392 14841 9404 14844
rect 9438 14872 9450 14875
rect 9490 14872 9496 14884
rect 9438 14844 9496 14872
rect 9438 14841 9450 14844
rect 9392 14835 9450 14841
rect 9490 14832 9496 14844
rect 9548 14832 9554 14884
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14872 11943 14875
rect 12802 14872 12808 14884
rect 11931 14844 12808 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 12912 14816 12940 14912
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5316 14776 5641 14804
rect 5316 14764 5322 14776
rect 5629 14773 5641 14776
rect 5675 14773 5687 14807
rect 5629 14767 5687 14773
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 5776 14776 6561 14804
rect 5776 14764 5782 14776
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 6595 14776 7297 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7285 14773 7297 14776
rect 7331 14804 7343 14807
rect 9214 14804 9220 14816
rect 7331 14776 9220 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12216 14776 12449 14804
rect 12216 14764 12222 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12894 14804 12900 14816
rect 12855 14776 12900 14804
rect 12437 14767 12495 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 5868 14572 7297 14600
rect 5868 14560 5874 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 7285 14563 7343 14569
rect 7929 14603 7987 14609
rect 7929 14569 7941 14603
rect 7975 14600 7987 14603
rect 8202 14600 8208 14612
rect 7975 14572 8208 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 8849 14603 8907 14609
rect 8849 14569 8861 14603
rect 8895 14600 8907 14603
rect 9030 14600 9036 14612
rect 8895 14572 9036 14600
rect 8895 14569 8907 14572
rect 8849 14563 8907 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9582 14600 9588 14612
rect 9539 14572 9588 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 11609 14603 11667 14609
rect 11609 14569 11621 14603
rect 11655 14600 11667 14603
rect 12069 14603 12127 14609
rect 12069 14600 12081 14603
rect 11655 14572 12081 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 12069 14569 12081 14572
rect 12115 14600 12127 14603
rect 12158 14600 12164 14612
rect 12115 14572 12164 14600
rect 12115 14569 12127 14572
rect 12069 14563 12127 14569
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12710 14600 12716 14612
rect 12671 14572 12716 14600
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12860 14572 13277 14600
rect 12860 14560 12866 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 1670 14532 1676 14544
rect 1631 14504 1676 14532
rect 1670 14492 1676 14504
rect 1728 14492 1734 14544
rect 6178 14473 6184 14476
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 6172 14464 6184 14473
rect 1443 14436 1716 14464
rect 6091 14436 6184 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1688 14408 1716 14436
rect 6172 14427 6184 14436
rect 6236 14464 6242 14476
rect 7282 14464 7288 14476
rect 6236 14436 7288 14464
rect 6178 14424 6184 14427
rect 6236 14424 6242 14436
rect 7282 14424 7288 14436
rect 7340 14424 7346 14476
rect 10502 14464 10508 14476
rect 10463 14436 10508 14464
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 10652 14436 10697 14464
rect 10652 14424 10658 14436
rect 1670 14356 1676 14408
rect 1728 14356 1734 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 5592 14368 5917 14396
rect 5592 14356 5598 14368
rect 5905 14365 5917 14368
rect 5951 14365 5963 14399
rect 10686 14396 10692 14408
rect 10647 14368 10692 14396
rect 5905 14359 5963 14365
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12308 14368 12353 14396
rect 12308 14356 12314 14368
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 9953 14331 10011 14337
rect 9953 14328 9965 14331
rect 9732 14300 9965 14328
rect 9732 14288 9738 14300
rect 9953 14297 9965 14300
rect 9999 14328 10011 14331
rect 10318 14328 10324 14340
rect 9999 14300 10324 14328
rect 9999 14297 10011 14300
rect 9953 14291 10011 14297
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 10502 14288 10508 14340
rect 10560 14328 10566 14340
rect 11701 14331 11759 14337
rect 11701 14328 11713 14331
rect 10560 14300 11713 14328
rect 10560 14288 10566 14300
rect 11701 14297 11713 14300
rect 11747 14297 11759 14331
rect 11701 14291 11759 14297
rect 5258 14260 5264 14272
rect 5219 14232 5264 14260
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 10134 14260 10140 14272
rect 10095 14232 10140 14260
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 11112 14232 11161 14260
rect 11112 14220 11118 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 5316 14028 6837 14056
rect 5316 14016 5322 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 8110 14056 8116 14068
rect 7524 14028 8116 14056
rect 7524 14016 7530 14028
rect 8110 14016 8116 14028
rect 8168 14056 8174 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8168 14028 8585 14056
rect 8168 14016 8174 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 8573 14019 8631 14025
rect 8757 14059 8815 14065
rect 8757 14025 8769 14059
rect 8803 14056 8815 14059
rect 9582 14056 9588 14068
rect 8803 14028 9588 14056
rect 8803 14025 8815 14028
rect 8757 14019 8815 14025
rect 1670 13988 1676 14000
rect 1631 13960 1676 13988
rect 1670 13948 1676 13960
rect 1728 13948 1734 14000
rect 5626 13948 5632 14000
rect 5684 13988 5690 14000
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 5684 13960 6561 13988
rect 5684 13948 5690 13960
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 5905 13923 5963 13929
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 6178 13920 6184 13932
rect 5951 13892 6184 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 5534 13852 5540 13864
rect 5495 13824 5540 13852
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 6564 13852 6592 13951
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7248 13892 7297 13920
rect 7248 13880 7254 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7374 13880 7380 13932
rect 7432 13920 7438 13932
rect 8588 13920 8616 14019
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10594 14056 10600 14068
rect 10555 14028 10600 14056
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11572 14028 11805 14056
rect 11572 14016 11578 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 11793 14019 11851 14025
rect 8662 13948 8668 14000
rect 8720 13988 8726 14000
rect 9122 13988 9128 14000
rect 8720 13960 9128 13988
rect 8720 13948 8726 13960
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 10229 13991 10287 13997
rect 10229 13957 10241 13991
rect 10275 13988 10287 13991
rect 10704 13988 10732 14016
rect 10275 13960 10732 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 7432 13892 7477 13920
rect 8588 13892 9229 13920
rect 7432 13880 7438 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9490 13920 9496 13932
rect 9447 13892 9496 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 10744 13892 11161 13920
rect 10744 13880 10750 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11808 13920 11836 14019
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 12216 14028 12449 14056
rect 12216 14016 12222 14028
rect 12437 14025 12449 14028
rect 12483 14056 12495 14059
rect 13449 14059 13507 14065
rect 13449 14056 13461 14059
rect 12483 14028 13461 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 13449 14025 13461 14028
rect 13495 14025 13507 14059
rect 13449 14019 13507 14025
rect 12710 13920 12716 13932
rect 11808 13892 12716 13920
rect 11149 13883 11207 13889
rect 12710 13880 12716 13892
rect 12768 13920 12774 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12768 13892 13001 13920
rect 12768 13880 12774 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 9861 13855 9919 13861
rect 6564 13824 6868 13852
rect 6840 13784 6868 13824
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 11054 13852 11060 13864
rect 9907 13824 10916 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 6840 13756 7205 13784
rect 7193 13753 7205 13756
rect 7239 13753 7251 13787
rect 7193 13747 7251 13753
rect 9125 13787 9183 13793
rect 9125 13753 9137 13787
rect 9171 13784 9183 13787
rect 9306 13784 9312 13796
rect 9171 13756 9312 13784
rect 9171 13753 9183 13756
rect 9125 13747 9183 13753
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 10888 13728 10916 13824
rect 10980 13824 11060 13852
rect 10980 13793 11008 13824
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13078 13852 13084 13864
rect 12943 13824 13084 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 10965 13787 11023 13793
rect 10965 13753 10977 13787
rect 11011 13753 11023 13787
rect 10965 13747 11023 13753
rect 12805 13787 12863 13793
rect 12805 13753 12817 13787
rect 12851 13784 12863 13787
rect 12986 13784 12992 13796
rect 12851 13756 12992 13784
rect 12851 13753 12863 13756
rect 12805 13747 12863 13753
rect 10870 13716 10876 13728
rect 10783 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13716 10934 13728
rect 11057 13719 11115 13725
rect 11057 13716 11069 13719
rect 10928 13688 11069 13716
rect 10928 13676 10934 13688
rect 11057 13685 11069 13688
rect 11103 13685 11115 13719
rect 11057 13679 11115 13685
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 12820 13716 12848 13747
rect 12986 13744 12992 13756
rect 13044 13784 13050 13796
rect 13814 13784 13820 13796
rect 13044 13756 13820 13784
rect 13044 13744 13050 13756
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 12299 13688 12848 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 6914 13512 6920 13524
rect 6827 13484 6920 13512
rect 6914 13472 6920 13484
rect 6972 13512 6978 13524
rect 7190 13512 7196 13524
rect 6972 13484 7196 13512
rect 6972 13472 6978 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 8849 13515 8907 13521
rect 8849 13512 8861 13515
rect 8720 13484 8861 13512
rect 8720 13472 8726 13484
rect 8849 13481 8861 13484
rect 8895 13512 8907 13515
rect 9306 13512 9312 13524
rect 8895 13484 9312 13512
rect 8895 13481 8907 13484
rect 8849 13475 8907 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 11054 13512 11060 13524
rect 10919 13484 11060 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11422 13512 11428 13524
rect 11287 13484 11428 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13354 13512 13360 13524
rect 13044 13484 13360 13512
rect 13044 13472 13050 13484
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 10229 13447 10287 13453
rect 10229 13413 10241 13447
rect 10275 13444 10287 13447
rect 10594 13444 10600 13456
rect 10275 13416 10600 13444
rect 10275 13413 10287 13416
rect 10229 13407 10287 13413
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 10704 13444 10732 13472
rect 11885 13447 11943 13453
rect 11885 13444 11897 13447
rect 10704 13416 11897 13444
rect 11885 13413 11897 13416
rect 11931 13444 11943 13447
rect 12250 13444 12256 13456
rect 11931 13416 12256 13444
rect 11931 13413 11943 13416
rect 11885 13407 11943 13413
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 12802 13444 12808 13456
rect 12575 13416 12808 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 12802 13404 12808 13416
rect 12860 13444 12866 13456
rect 13078 13444 13084 13456
rect 12860 13416 13084 13444
rect 12860 13404 12866 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11296 13280 11345 13308
rect 11296 13268 11302 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11514 13308 11520 13320
rect 11475 13280 11520 13308
rect 11333 13271 11391 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4062 13172 4068 13184
rect 3476 13144 4068 13172
rect 3476 13132 3482 13144
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 7926 13172 7932 13184
rect 7887 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13172 7990 13184
rect 8294 13172 8300 13184
rect 7984 13144 8300 13172
rect 7984 13132 7990 13144
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 10229 12971 10287 12977
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 10502 12968 10508 12980
rect 10275 12940 10508 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 11422 12968 11428 12980
rect 11011 12940 11428 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11572 12940 11621 12968
rect 11572 12928 11578 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 11609 12931 11667 12937
rect 11440 12900 11468 12928
rect 12250 12900 12256 12912
rect 11440 12872 12256 12900
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 10318 12792 10324 12844
rect 10376 12832 10382 12844
rect 10502 12832 10508 12844
rect 10376 12804 10508 12832
rect 10376 12792 10382 12804
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 7926 12764 7932 12776
rect 7887 12736 7932 12764
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8202 12705 8208 12708
rect 7837 12699 7895 12705
rect 7837 12665 7849 12699
rect 7883 12696 7895 12699
rect 8174 12699 8208 12705
rect 8174 12696 8186 12699
rect 7883 12668 8186 12696
rect 7883 12665 7895 12668
rect 7837 12659 7895 12665
rect 8174 12665 8186 12668
rect 8260 12696 8266 12708
rect 8260 12668 8322 12696
rect 8174 12659 8208 12665
rect 8202 12656 8208 12659
rect 8260 12656 8266 12668
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11333 12699 11391 12705
rect 11333 12696 11345 12699
rect 11296 12668 11345 12696
rect 11296 12656 11302 12668
rect 11333 12665 11345 12668
rect 11379 12696 11391 12699
rect 11422 12696 11428 12708
rect 11379 12668 11428 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9490 12628 9496 12640
rect 9355 12600 9496 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 11514 12588 11520 12640
rect 11572 12628 11578 12640
rect 12618 12628 12624 12640
rect 11572 12600 12624 12628
rect 11572 12588 11578 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 5810 12424 5816 12436
rect 5684 12396 5816 12424
rect 5684 12384 5690 12396
rect 5810 12384 5816 12396
rect 5868 12384 5874 12436
rect 9766 12384 9772 12436
rect 9824 12384 9830 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 9916 12396 10272 12424
rect 9916 12384 9922 12396
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8662 12356 8668 12368
rect 8352 12328 8668 12356
rect 8352 12316 8358 12328
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 9784 12356 9812 12384
rect 10244 12368 10272 12396
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 9784 12328 10057 12356
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 10226 12316 10232 12368
rect 10284 12316 10290 12368
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 11146 12356 11152 12368
rect 10744 12328 11152 12356
rect 10744 12316 10750 12328
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 4614 12288 4620 12300
rect 4575 12260 4620 12288
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7975 12260 8401 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8389 12257 8401 12260
rect 8435 12288 8447 12291
rect 9582 12288 9588 12300
rect 8435 12260 9588 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10597 12291 10655 12297
rect 10597 12288 10609 12291
rect 9916 12260 10609 12288
rect 9916 12248 9922 12260
rect 10597 12257 10609 12260
rect 10643 12288 10655 12291
rect 10873 12291 10931 12297
rect 10873 12288 10885 12291
rect 10643 12260 10885 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 10873 12257 10885 12260
rect 10919 12257 10931 12291
rect 10873 12251 10931 12257
rect 11238 12248 11244 12300
rect 11296 12288 11302 12300
rect 11405 12291 11463 12297
rect 11405 12288 11417 12291
rect 11296 12260 11417 12288
rect 11296 12248 11302 12260
rect 11405 12257 11417 12260
rect 11451 12257 11463 12291
rect 11405 12251 11463 12257
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 4246 12220 4252 12232
rect 3927 12192 4252 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4396 12192 4721 12220
rect 4396 12180 4402 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4890 12220 4896 12232
rect 4803 12192 4896 12220
rect 4709 12183 4767 12189
rect 4890 12180 4896 12192
rect 4948 12220 4954 12232
rect 5718 12220 5724 12232
rect 4948 12192 5724 12220
rect 4948 12180 4954 12192
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 8754 12220 8760 12232
rect 8711 12192 8760 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 8680 12152 8708 12183
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 11146 12220 11152 12232
rect 10704 12192 11152 12220
rect 10042 12152 10048 12164
rect 8260 12124 8708 12152
rect 10003 12124 10048 12152
rect 8260 12112 8266 12124
rect 10042 12112 10048 12124
rect 10100 12152 10106 12164
rect 10704 12161 10732 12192
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 10100 12124 10149 12152
rect 10100 12112 10106 12124
rect 10137 12121 10149 12124
rect 10183 12121 10195 12155
rect 10137 12115 10195 12121
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12121 10747 12155
rect 10689 12115 10747 12121
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 4120 12056 4261 12084
rect 4120 12044 4126 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 4249 12047 4307 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12618 12084 12624 12096
rect 12575 12056 12624 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 3789 11883 3847 11889
rect 3789 11849 3801 11883
rect 3835 11880 3847 11883
rect 4890 11880 4896 11892
rect 3835 11852 4896 11880
rect 3835 11849 3847 11852
rect 3789 11843 3847 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 7926 11880 7932 11892
rect 7668 11852 7932 11880
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 7668 11753 7696 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 8628 11852 10149 11880
rect 8628 11840 8634 11852
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 11238 11880 11244 11892
rect 11199 11852 11244 11880
rect 10137 11843 10195 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 12434 11880 12440 11892
rect 12395 11852 12440 11880
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 9950 11812 9956 11824
rect 9911 11784 9956 11812
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 7653 11747 7711 11753
rect 4203 11716 4384 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 4246 11676 4252 11688
rect 4207 11648 4252 11676
rect 1397 11639 1455 11645
rect 1412 11608 1440 11639
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 4356 11676 4384 11716
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 12158 11744 12164 11756
rect 12119 11716 12164 11744
rect 10689 11707 10747 11713
rect 4522 11685 4528 11688
rect 4505 11679 4528 11685
rect 4505 11676 4517 11679
rect 4356 11648 4517 11676
rect 4505 11645 4517 11648
rect 4580 11676 4586 11688
rect 7561 11679 7619 11685
rect 4580 11648 4653 11676
rect 4505 11639 4528 11645
rect 4522 11636 4528 11639
rect 4580 11636 4586 11648
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 7920 11679 7978 11685
rect 7920 11676 7932 11679
rect 7607 11648 7932 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 7920 11645 7932 11648
rect 7966 11676 7978 11679
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 7966 11648 9689 11676
rect 7966 11645 7978 11648
rect 7920 11639 7978 11645
rect 9677 11645 9689 11648
rect 9723 11676 9735 11679
rect 10502 11676 10508 11688
rect 9723 11648 10508 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 10704 11676 10732 11707
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12676 11716 13001 11744
rect 12676 11704 12682 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 10560 11648 10732 11676
rect 10560 11636 10566 11648
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 13078 11676 13084 11688
rect 12584 11648 13084 11676
rect 12584 11636 12590 11648
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 2222 11608 2228 11620
rect 1412 11580 2228 11608
rect 2222 11568 2228 11580
rect 2280 11568 2286 11620
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11608 3479 11611
rect 4338 11608 4344 11620
rect 3467 11580 4344 11608
rect 3467 11577 3479 11580
rect 3421 11571 3479 11577
rect 4338 11568 4344 11580
rect 4396 11568 4402 11620
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11608 7251 11611
rect 7239 11580 7880 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 5718 11540 5724 11552
rect 5675 11512 5724 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 7852 11540 7880 11580
rect 10042 11568 10048 11620
rect 10100 11608 10106 11620
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 10100 11580 10609 11608
rect 10100 11568 10106 11580
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 10597 11571 10655 11577
rect 11808 11580 12909 11608
rect 8754 11540 8760 11552
rect 7852 11512 8760 11540
rect 8754 11500 8760 11512
rect 8812 11540 8818 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8812 11512 9045 11540
rect 8812 11500 8818 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 9033 11503 9091 11509
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10008 11512 10517 11540
rect 10008 11500 10014 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11808 11549 11836 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11112 11512 11805 11540
rect 11112 11500 11118 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12216 11512 12817 11540
rect 12216 11500 12222 11512
rect 12805 11509 12817 11512
rect 12851 11540 12863 11543
rect 13722 11540 13728 11552
rect 12851 11512 13728 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 4801 11339 4859 11345
rect 4801 11336 4813 11339
rect 4304 11308 4813 11336
rect 4304 11296 4310 11308
rect 4801 11305 4813 11308
rect 4847 11305 4859 11339
rect 7742 11336 7748 11348
rect 7703 11308 7748 11336
rect 4801 11299 4859 11305
rect 3881 11271 3939 11277
rect 3881 11237 3893 11271
rect 3927 11268 3939 11271
rect 4614 11268 4620 11280
rect 3927 11240 4620 11268
rect 3927 11237 3939 11240
rect 3881 11231 3939 11237
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 4816 11268 4844 11299
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8018 11296 8024 11348
rect 8076 11336 8082 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 8076 11308 8125 11336
rect 8076 11296 8082 11308
rect 8113 11305 8125 11308
rect 8159 11336 8171 11339
rect 8159 11308 8248 11336
rect 8159 11305 8171 11308
rect 8113 11299 8171 11305
rect 5442 11268 5448 11280
rect 4816 11240 5448 11268
rect 4522 11200 4528 11212
rect 4483 11172 4528 11200
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 5092 11209 5120 11240
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 6822 11228 6828 11280
rect 6880 11268 6886 11280
rect 7101 11271 7159 11277
rect 7101 11268 7113 11271
rect 6880 11240 7113 11268
rect 6880 11228 6886 11240
rect 7101 11237 7113 11240
rect 7147 11268 7159 11271
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 7147 11240 7665 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 7653 11237 7665 11240
rect 7699 11268 7711 11271
rect 7926 11268 7932 11280
rect 7699 11240 7932 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 8220 11268 8248 11308
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8536 11308 8769 11336
rect 8536 11296 8542 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9950 11336 9956 11348
rect 9548 11308 9956 11336
rect 9548 11296 9554 11308
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 11238 11336 11244 11348
rect 11103 11308 11244 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12618 11336 12624 11348
rect 12575 11308 12624 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 8570 11268 8576 11280
rect 8220 11240 8576 11268
rect 8570 11228 8576 11240
rect 8628 11228 8634 11280
rect 11146 11268 11152 11280
rect 9692 11240 11152 11268
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5344 11203 5402 11209
rect 5344 11169 5356 11203
rect 5390 11200 5402 11203
rect 5718 11200 5724 11212
rect 5390 11172 5724 11200
rect 5390 11169 5402 11172
rect 5344 11163 5402 11169
rect 5000 11132 5028 11163
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 8202 11132 8208 11144
rect 4172 11104 5028 11132
rect 8163 11104 8208 11132
rect 3053 10999 3111 11005
rect 3053 10965 3065 10999
rect 3099 10996 3111 10999
rect 3326 10996 3332 11008
rect 3099 10968 3332 10996
rect 3099 10965 3111 10968
rect 3053 10959 3111 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4172 10996 4200 11104
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 8312 11064 8340 11095
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9692 11141 9720 11240
rect 11146 11228 11152 11240
rect 11204 11268 11210 11280
rect 11609 11271 11667 11277
rect 11609 11268 11621 11271
rect 11204 11240 11621 11268
rect 11204 11228 11210 11240
rect 11609 11237 11621 11240
rect 11655 11237 11667 11271
rect 11609 11231 11667 11237
rect 9950 11209 9956 11212
rect 9944 11200 9956 11209
rect 9911 11172 9956 11200
rect 9944 11163 9956 11172
rect 9950 11160 9956 11163
rect 10008 11160 10014 11212
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9640 11104 9689 11132
rect 9640 11092 9646 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 7984 11036 8340 11064
rect 7984 11024 7990 11036
rect 6454 10996 6460 11008
rect 4028 10968 4200 10996
rect 6415 10968 6460 10996
rect 4028 10956 4034 10968
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 4614 10792 4620 10804
rect 4571 10764 4620 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5905 10795 5963 10801
rect 5905 10792 5917 10795
rect 5592 10764 5917 10792
rect 5592 10752 5598 10764
rect 5905 10761 5917 10764
rect 5951 10761 5963 10795
rect 5905 10755 5963 10761
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 8628 10764 8769 10792
rect 8628 10752 8634 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 9582 10792 9588 10804
rect 9447 10764 9588 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 10962 10792 10968 10804
rect 10643 10764 10968 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 6454 10724 6460 10736
rect 3528 10696 6460 10724
rect 3528 10665 3556 10696
rect 6454 10684 6460 10696
rect 6512 10724 6518 10736
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 6512 10696 6561 10724
rect 6512 10684 6518 10696
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 2915 10628 3525 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4580 10628 5089 10656
rect 4580 10616 4586 10628
rect 5077 10625 5089 10628
rect 5123 10625 5135 10659
rect 6564 10656 6592 10687
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 9677 10727 9735 10733
rect 9677 10724 9689 10727
rect 7984 10696 9689 10724
rect 7984 10684 7990 10696
rect 9677 10693 9689 10696
rect 9723 10724 9735 10727
rect 9950 10724 9956 10736
rect 9723 10696 9956 10724
rect 9723 10693 9735 10696
rect 9677 10687 9735 10693
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 10505 10727 10563 10733
rect 10505 10693 10517 10727
rect 10551 10724 10563 10727
rect 10686 10724 10692 10736
rect 10551 10696 10692 10724
rect 10551 10693 10563 10696
rect 10505 10687 10563 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 6564 10628 6960 10656
rect 5077 10619 5135 10625
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3108 10560 3433 10588
rect 3108 10548 3114 10560
rect 3421 10557 3433 10560
rect 3467 10588 3479 10591
rect 4062 10588 4068 10600
rect 3467 10560 4068 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6932 10588 6960 10628
rect 7081 10591 7139 10597
rect 7081 10588 7093 10591
rect 6932 10560 7093 10588
rect 7081 10557 7093 10560
rect 7127 10557 7139 10591
rect 10704 10588 10732 10684
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 11238 10656 11244 10668
rect 10836 10628 11244 10656
rect 10836 10616 10842 10628
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 10704 10560 11069 10588
rect 7081 10551 7139 10557
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 4985 10523 5043 10529
rect 4985 10489 4997 10523
rect 5031 10520 5043 10523
rect 5074 10520 5080 10532
rect 5031 10492 5080 10520
rect 5031 10489 5043 10492
rect 4985 10483 5043 10489
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 2958 10452 2964 10464
rect 2919 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3970 10452 3976 10464
rect 3931 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4890 10452 4896 10464
rect 4479 10424 4896 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 5718 10452 5724 10464
rect 5675 10424 5724 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 7616 10424 8217 10452
rect 7616 10412 7622 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 9640 10424 10149 10452
rect 9640 10412 9646 10424
rect 10137 10421 10149 10424
rect 10183 10452 10195 10455
rect 10594 10452 10600 10464
rect 10183 10424 10600 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 10594 10412 10600 10424
rect 10652 10452 10658 10464
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 10652 10424 10977 10452
rect 10652 10412 10658 10424
rect 10965 10421 10977 10424
rect 11011 10421 11023 10455
rect 10965 10415 11023 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 3384 10220 5089 10248
rect 3384 10208 3390 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5077 10211 5135 10217
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6638 10248 6644 10260
rect 6052 10220 6644 10248
rect 6052 10208 6058 10220
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7558 10248 7564 10260
rect 7519 10220 7564 10248
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 7193 10183 7251 10189
rect 7193 10149 7205 10183
rect 7239 10180 7251 10183
rect 7374 10180 7380 10192
rect 7239 10152 7380 10180
rect 7239 10149 7251 10152
rect 7193 10143 7251 10149
rect 7374 10140 7380 10152
rect 7432 10180 7438 10192
rect 8110 10180 8116 10192
rect 7432 10152 8116 10180
rect 7432 10140 7438 10152
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8588 10180 8616 10211
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10042 10248 10048 10260
rect 9732 10220 10048 10248
rect 9732 10208 9738 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10226 10248 10232 10260
rect 10183 10220 10232 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10778 10248 10784 10260
rect 10739 10220 10784 10248
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 9858 10180 9864 10192
rect 8588 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3326 10112 3332 10124
rect 3200 10084 3332 10112
rect 3200 10072 3206 10084
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 4982 10072 4988 10124
rect 5040 10112 5046 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5040 10084 5457 10112
rect 5040 10072 5046 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 8570 10072 8576 10124
rect 8628 10112 8634 10124
rect 8757 10115 8815 10121
rect 8757 10112 8769 10115
rect 8628 10084 8769 10112
rect 8628 10072 8634 10084
rect 8757 10081 8769 10084
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4212 10016 4629 10044
rect 4212 10004 4218 10016
rect 4617 10013 4629 10016
rect 4663 10044 4675 10047
rect 5074 10044 5080 10056
rect 4663 10016 5080 10044
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5224 10016 5549 10044
rect 5224 10004 5230 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5537 10007 5595 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 6638 10044 6644 10056
rect 6599 10016 6644 10044
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 10502 10044 10508 10056
rect 10367 10016 10508 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 9677 9979 9735 9985
rect 9677 9945 9689 9979
rect 9723 9976 9735 9979
rect 9766 9976 9772 9988
rect 9723 9948 9772 9976
rect 9723 9945 9735 9948
rect 9677 9939 9735 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 4982 9908 4988 9920
rect 4943 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 4522 9704 4528 9716
rect 4387 9676 4528 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 5776 9676 6193 9704
rect 5776 9664 5782 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 6181 9667 6239 9673
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 8573 9707 8631 9713
rect 8573 9704 8585 9707
rect 8352 9676 8585 9704
rect 8352 9664 8358 9676
rect 8573 9673 8585 9676
rect 8619 9673 8631 9707
rect 10042 9704 10048 9716
rect 10003 9676 10048 9704
rect 8573 9667 8631 9673
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 5442 9636 5448 9648
rect 3384 9608 5448 9636
rect 3384 9596 3390 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 9766 9636 9772 9648
rect 9679 9608 9772 9636
rect 9766 9596 9772 9608
rect 9824 9636 9830 9648
rect 10226 9636 10232 9648
rect 9824 9608 10232 9636
rect 9824 9596 9830 9608
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 5718 9568 5724 9580
rect 4580 9540 5724 9568
rect 4580 9528 4586 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7098 9568 7104 9580
rect 6687 9540 7104 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 8754 9568 8760 9580
rect 8527 9540 8760 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 8754 9528 8760 9540
rect 8812 9568 8818 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8812 9540 9137 9568
rect 8812 9528 8818 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 4706 9500 4712 9512
rect 4619 9472 4712 9500
rect 4706 9460 4712 9472
rect 4764 9500 4770 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 4764 9472 5641 9500
rect 4764 9460 4770 9472
rect 5629 9469 5641 9472
rect 5675 9500 5687 9503
rect 6822 9500 6828 9512
rect 5675 9472 6828 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7374 9500 7380 9512
rect 7335 9472 7380 9500
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 8662 9500 8668 9512
rect 8444 9472 8668 9500
rect 8444 9460 8450 9472
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5123 9404 5580 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 5166 9364 5172 9376
rect 5127 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5552 9373 5580 9404
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 8021 9435 8079 9441
rect 8021 9432 8033 9435
rect 6972 9404 8033 9432
rect 6972 9392 6978 9404
rect 8021 9401 8033 9404
rect 8067 9432 8079 9435
rect 9033 9435 9091 9441
rect 9033 9432 9045 9435
rect 8067 9404 9045 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 9033 9401 9045 9404
rect 9079 9401 9091 9435
rect 9033 9395 9091 9401
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7466 9364 7472 9376
rect 7156 9336 7472 9364
rect 7156 9324 7162 9336
rect 7466 9324 7472 9336
rect 7524 9364 7530 9376
rect 7926 9364 7932 9376
rect 7524 9336 7932 9364
rect 7524 9324 7530 9336
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 8720 9336 8953 9364
rect 8720 9324 8726 9336
rect 8941 9333 8953 9336
rect 8987 9333 8999 9367
rect 10502 9364 10508 9376
rect 10463 9336 10508 9364
rect 8941 9327 8999 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 4338 9160 4344 9172
rect 4299 9132 4344 9160
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 5721 9163 5779 9169
rect 5721 9160 5733 9163
rect 5224 9132 5733 9160
rect 5224 9120 5230 9132
rect 5721 9129 5733 9132
rect 5767 9129 5779 9163
rect 5721 9123 5779 9129
rect 6181 9163 6239 9169
rect 6181 9129 6193 9163
rect 6227 9160 6239 9163
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 6227 9132 6469 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 6457 9129 6469 9132
rect 6503 9160 6515 9163
rect 7466 9160 7472 9172
rect 6503 9132 7472 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 7466 9120 7472 9132
rect 7524 9160 7530 9172
rect 8570 9160 8576 9172
rect 7524 9132 8576 9160
rect 7524 9120 7530 9132
rect 8570 9120 8576 9132
rect 8628 9160 8634 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8628 9132 9045 9160
rect 8628 9120 8634 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 5445 9095 5503 9101
rect 5445 9061 5457 9095
rect 5491 9092 5503 9095
rect 5534 9092 5540 9104
rect 5491 9064 5540 9092
rect 5491 9061 5503 9064
rect 5445 9055 5503 9061
rect 5534 9052 5540 9064
rect 5592 9092 5598 9104
rect 6638 9092 6644 9104
rect 5592 9064 6644 9092
rect 5592 9052 5598 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 7000 9095 7058 9101
rect 7000 9061 7012 9095
rect 7046 9092 7058 9095
rect 7098 9092 7104 9104
rect 7046 9064 7104 9092
rect 7046 9061 7058 9064
rect 7000 9055 7058 9061
rect 7098 9052 7104 9064
rect 7156 9092 7162 9104
rect 7558 9092 7564 9104
rect 7156 9064 7564 9092
rect 7156 9052 7162 9064
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 4488 8996 4721 9024
rect 4488 8984 4494 8996
rect 4709 8993 4721 8996
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 6181 9027 6239 9033
rect 6181 9024 6193 9027
rect 6135 8996 6193 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 6181 8993 6193 8996
rect 6227 8993 6239 9027
rect 6181 8987 6239 8993
rect 4798 8956 4804 8968
rect 4759 8928 4804 8956
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 6730 8956 6736 8968
rect 6691 8928 6736 8956
rect 4893 8919 4951 8925
rect 4522 8848 4528 8900
rect 4580 8888 4586 8900
rect 4908 8888 4936 8919
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 4580 8860 4936 8888
rect 4580 8848 4586 8860
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 4028 8792 5917 8820
rect 4028 8780 4034 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 8110 8820 8116 8832
rect 8071 8792 8116 8820
rect 5905 8783 5963 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8662 8820 8668 8832
rect 8352 8792 8668 8820
rect 8352 8780 8358 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10410 8820 10416 8832
rect 10091 8792 10416 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4430 8616 4436 8628
rect 4391 8588 4436 8616
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 5040 8588 5181 8616
rect 5040 8576 5046 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 9125 8619 9183 8625
rect 9125 8585 9137 8619
rect 9171 8616 9183 8619
rect 9398 8616 9404 8628
rect 9171 8588 9404 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 7392 8520 7941 8548
rect 5718 8480 5724 8492
rect 5679 8452 5724 8480
rect 5718 8440 5724 8452
rect 5776 8480 5782 8492
rect 6178 8480 6184 8492
rect 5776 8452 6184 8480
rect 5776 8440 5782 8452
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7392 8489 7420 8520
rect 7929 8517 7941 8520
rect 7975 8517 7987 8551
rect 7929 8511 7987 8517
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7064 8452 7389 8480
rect 7064 8440 7070 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7558 8480 7564 8492
rect 7471 8452 7564 8480
rect 7377 8443 7435 8449
rect 7558 8440 7564 8452
rect 7616 8480 7622 8492
rect 8110 8480 8116 8492
rect 7616 8452 8116 8480
rect 7616 8440 7622 8452
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 2409 8415 2467 8421
rect 2409 8381 2421 8415
rect 2455 8412 2467 8415
rect 2498 8412 2504 8424
rect 2455 8384 2504 8412
rect 2455 8381 2467 8384
rect 2409 8375 2467 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 5534 8412 5540 8424
rect 5495 8384 5540 8412
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 6638 8412 6644 8424
rect 5684 8384 5729 8412
rect 6551 8384 6644 8412
rect 5684 8372 5690 8384
rect 6638 8372 6644 8384
rect 6696 8412 6702 8424
rect 7282 8412 7288 8424
rect 6696 8384 7288 8412
rect 6696 8372 6702 8384
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 9140 8412 9168 8579
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 10594 8480 10600 8492
rect 9539 8452 10364 8480
rect 10555 8452 10600 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 8527 8384 9168 8412
rect 9769 8415 9827 8421
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 9858 8412 9864 8424
rect 9815 8384 9864 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10336 8421 10364 8452
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10962 8412 10968 8424
rect 10367 8384 10968 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 2317 8347 2375 8353
rect 2317 8313 2329 8347
rect 2363 8344 2375 8347
rect 2590 8344 2596 8356
rect 2363 8316 2596 8344
rect 2363 8313 2375 8316
rect 2317 8307 2375 8313
rect 2590 8304 2596 8316
rect 2648 8353 2654 8356
rect 2648 8347 2712 8353
rect 2648 8313 2666 8347
rect 2700 8313 2712 8347
rect 2648 8307 2712 8313
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5644 8344 5672 8372
rect 10410 8344 10416 8356
rect 5123 8316 5672 8344
rect 10371 8316 10416 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 2648 8304 2654 8307
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 3789 8279 3847 8285
rect 3789 8276 3801 8279
rect 3568 8248 3801 8276
rect 3568 8236 3574 8248
rect 3789 8245 3801 8248
rect 3835 8245 3847 8279
rect 6914 8276 6920 8288
rect 6875 8248 6920 8276
rect 3789 8239 3847 8245
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 8389 8279 8447 8285
rect 8389 8245 8401 8279
rect 8435 8276 8447 8279
rect 8478 8276 8484 8288
rect 8435 8248 8484 8276
rect 8435 8245 8447 8248
rect 8389 8239 8447 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8662 8276 8668 8288
rect 8623 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9582 8276 9588 8288
rect 9088 8248 9588 8276
rect 9088 8236 9094 8248
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 9950 8276 9956 8288
rect 9911 8248 9956 8276
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4522 8072 4528 8084
rect 4479 8044 4528 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 4798 8072 4804 8084
rect 4759 8044 4804 8072
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 6236 8044 6377 8072
rect 6236 8032 6242 8044
rect 6365 8041 6377 8044
rect 6411 8041 6423 8075
rect 6365 8035 6423 8041
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7098 8072 7104 8084
rect 7055 8044 7104 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 8021 8075 8079 8081
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 8294 8072 8300 8084
rect 8067 8044 8300 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 9030 8072 9036 8084
rect 8991 8044 9036 8072
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10134 8072 10140 8084
rect 10091 8044 10140 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10134 8032 10140 8044
rect 10192 8072 10198 8084
rect 10594 8072 10600 8084
rect 10192 8044 10600 8072
rect 10192 8032 10198 8044
rect 10594 8032 10600 8044
rect 10652 8072 10658 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 10652 8044 11989 8072
rect 10652 8032 10658 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 1670 8004 1676 8016
rect 1631 7976 1676 8004
rect 1670 7964 1676 7976
rect 1728 7964 1734 8016
rect 7377 8007 7435 8013
rect 7377 7973 7389 8007
rect 7423 8004 7435 8007
rect 7558 8004 7564 8016
rect 7423 7976 7564 8004
rect 7423 7973 7435 7976
rect 7377 7967 7435 7973
rect 7558 7964 7564 7976
rect 7616 7964 7622 8016
rect 9858 7964 9864 8016
rect 9916 8004 9922 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9916 7976 10333 8004
rect 9916 7964 9922 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2406 7936 2412 7948
rect 1443 7908 2412 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 5258 7945 5264 7948
rect 5252 7936 5264 7945
rect 5219 7908 5264 7936
rect 5252 7899 5264 7908
rect 5258 7896 5264 7899
rect 5316 7896 5322 7948
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 7834 7936 7840 7948
rect 7699 7908 7840 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 10864 7939 10922 7945
rect 10864 7905 10876 7939
rect 10910 7936 10922 7939
rect 11790 7936 11796 7948
rect 10910 7908 11796 7936
rect 10910 7905 10922 7908
rect 10864 7899 10922 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 4982 7868 4988 7880
rect 4943 7840 4988 7868
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 8478 7868 8484 7880
rect 8439 7840 8484 7868
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 8588 7800 8616 7831
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 10597 7871 10655 7877
rect 10597 7868 10609 7871
rect 9640 7840 10609 7868
rect 9640 7828 9646 7840
rect 10597 7837 10609 7840
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 8352 7772 8616 7800
rect 8352 7760 8358 7772
rect 2498 7732 2504 7744
rect 2411 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7732 2562 7744
rect 3329 7735 3387 7741
rect 3329 7732 3341 7735
rect 2556 7704 3341 7732
rect 2556 7692 2562 7704
rect 3329 7701 3341 7704
rect 3375 7732 3387 7735
rect 3418 7732 3424 7744
rect 3375 7704 3424 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 2406 7528 2412 7540
rect 2367 7500 2412 7528
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 3108 7500 3157 7528
rect 3108 7488 3114 7500
rect 3145 7497 3157 7500
rect 3191 7528 3203 7531
rect 3510 7528 3516 7540
rect 3191 7500 3516 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 7834 7528 7840 7540
rect 6319 7500 7840 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7528 11854 7540
rect 12434 7528 12440 7540
rect 11848 7500 12440 7528
rect 11848 7488 11854 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 5684 7432 6561 7460
rect 5684 7420 5690 7432
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 7374 7460 7380 7472
rect 7335 7432 7380 7460
rect 6549 7423 6607 7429
rect 3510 7333 3516 7336
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 3237 7327 3295 7333
rect 1443 7296 2084 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2056 7200 2084 7296
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 3504 7324 3516 7333
rect 3471 7296 3516 7324
rect 3237 7287 3295 7293
rect 3504 7287 3516 7296
rect 3252 7256 3280 7287
rect 3510 7284 3516 7287
rect 3568 7284 3574 7336
rect 6564 7324 6592 7423
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 6730 7324 6736 7336
rect 6564 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7392 7324 7420 7420
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9398 7392 9404 7404
rect 8987 7364 9404 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9815 7364 9996 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 7392 7296 8677 7324
rect 3418 7256 3424 7268
rect 3252 7228 3424 7256
rect 3418 7216 3424 7228
rect 3476 7256 3482 7268
rect 4982 7256 4988 7268
rect 3476 7228 4988 7256
rect 3476 7216 3482 7228
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5040 7228 5549 7256
rect 5040 7216 5046 7228
rect 5537 7225 5549 7228
rect 5583 7225 5595 7259
rect 5537 7219 5595 7225
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 7392 7256 7420 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9640 7296 9873 7324
rect 9640 7284 9646 7296
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9968 7324 9996 7364
rect 10134 7333 10140 7336
rect 10128 7324 10140 7333
rect 9968 7296 10140 7324
rect 9861 7287 9919 7293
rect 10128 7287 10140 7296
rect 8757 7259 8815 7265
rect 8757 7256 8769 7259
rect 5960 7228 7420 7256
rect 8128 7228 8769 7256
rect 5960 7216 5966 7228
rect 1394 7148 1400 7200
rect 1452 7188 1458 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 1452 7160 1593 7188
rect 1452 7148 1458 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 1581 7151 1639 7157
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7188 4678 7200
rect 5169 7191 5227 7197
rect 5169 7188 5181 7191
rect 4672 7160 5181 7188
rect 4672 7148 4678 7160
rect 5169 7157 5181 7160
rect 5215 7188 5227 7191
rect 5258 7188 5264 7200
rect 5215 7160 5264 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 7006 7188 7012 7200
rect 6967 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7834 7188 7840 7200
rect 7795 7160 7840 7188
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 8128 7197 8156 7228
rect 8757 7225 8769 7228
rect 8803 7225 8815 7259
rect 9876 7256 9904 7287
rect 10134 7284 10140 7287
rect 10192 7284 10198 7336
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 9876 7228 12173 7256
rect 8757 7219 8815 7225
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 8076 7160 8125 7188
rect 8076 7148 8082 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8113 7151 8171 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 11020 7160 11253 7188
rect 11020 7148 11026 7160
rect 11241 7157 11253 7160
rect 11287 7157 11299 7191
rect 11241 7151 11299 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 4617 6987 4675 6993
rect 4617 6953 4629 6987
rect 4663 6984 4675 6987
rect 4798 6984 4804 6996
rect 4663 6956 4804 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 4985 6987 5043 6993
rect 4985 6953 4997 6987
rect 5031 6984 5043 6987
rect 5074 6984 5080 6996
rect 5031 6956 5080 6984
rect 5031 6953 5043 6956
rect 4985 6947 5043 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6457 6987 6515 6993
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 6822 6984 6828 6996
rect 6503 6956 6828 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8021 6987 8079 6993
rect 8021 6953 8033 6987
rect 8067 6984 8079 6987
rect 8478 6984 8484 6996
rect 8067 6956 8484 6984
rect 8067 6953 8079 6956
rect 8021 6947 8079 6953
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 9582 6984 9588 6996
rect 9539 6956 9588 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 12529 6987 12587 6993
rect 12529 6984 12541 6987
rect 12032 6956 12541 6984
rect 12032 6944 12038 6956
rect 12529 6953 12541 6956
rect 12575 6953 12587 6987
rect 12529 6947 12587 6953
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 6917 6919 6975 6925
rect 6917 6916 6929 6919
rect 6788 6888 6929 6916
rect 6788 6876 6794 6888
rect 6917 6885 6929 6888
rect 6963 6916 6975 6919
rect 8294 6916 8300 6928
rect 6963 6888 8300 6916
rect 6963 6885 6975 6888
rect 6917 6879 6975 6885
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 8938 6916 8944 6928
rect 8444 6888 8944 6916
rect 8444 6876 8450 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 12676 6888 12721 6916
rect 12676 6876 12682 6888
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1578 6848 1584 6860
rect 1443 6820 1584 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3605 6851 3663 6857
rect 3605 6817 3617 6851
rect 3651 6848 3663 6851
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 3651 6820 3893 6848
rect 3651 6817 3663 6820
rect 3605 6811 3663 6817
rect 3881 6817 3893 6820
rect 3927 6848 3939 6851
rect 3970 6848 3976 6860
rect 3927 6820 3976 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 5442 6848 5448 6860
rect 5123 6820 5448 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6848 6423 6851
rect 6822 6848 6828 6860
rect 6411 6820 6828 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6848 9183 6851
rect 9398 6848 9404 6860
rect 9171 6820 9404 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 2648 6752 4353 6780
rect 2648 6740 2654 6752
rect 4341 6749 4353 6752
rect 4387 6780 4399 6783
rect 4890 6780 4896 6792
rect 4387 6752 4896 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 5184 6712 5212 6743
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6696 6752 7021 6780
rect 6696 6740 6702 6752
rect 7009 6749 7021 6752
rect 7055 6780 7067 6783
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7055 6752 7849 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7837 6749 7849 6752
rect 7883 6780 7895 6783
rect 8202 6780 8208 6792
rect 7883 6752 8208 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8478 6780 8484 6792
rect 8439 6752 8484 6780
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 9140 6780 9168 6811
rect 9398 6808 9404 6820
rect 9456 6848 9462 6860
rect 9950 6857 9956 6860
rect 9944 6848 9956 6857
rect 9456 6820 9956 6848
rect 9456 6808 9462 6820
rect 9944 6811 9956 6820
rect 10008 6848 10014 6860
rect 10962 6848 10968 6860
rect 10008 6820 10968 6848
rect 9950 6808 9956 6811
rect 10008 6808 10014 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 8711 6752 9168 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9640 6752 9689 6780
rect 9640 6740 9646 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 12710 6780 12716 6792
rect 11112 6752 12204 6780
rect 11112 6740 11118 6752
rect 4672 6684 5212 6712
rect 4672 6672 4678 6684
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 8938 6712 8944 6724
rect 5500 6684 8944 6712
rect 5500 6672 5506 6684
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 12176 6721 12204 6752
rect 12452 6752 12716 6780
rect 12452 6724 12480 6752
rect 12710 6740 12716 6752
rect 12768 6780 12774 6792
rect 13354 6780 13360 6792
rect 12768 6752 13360 6780
rect 12768 6740 12774 6752
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 12161 6715 12219 6721
rect 12161 6681 12173 6715
rect 12207 6681 12219 6715
rect 12161 6675 12219 6681
rect 12434 6672 12440 6724
rect 12492 6672 12498 6724
rect 934 6604 940 6656
rect 992 6644 998 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 992 6616 1593 6644
rect 992 6604 998 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1946 6644 1952 6656
rect 1907 6616 1952 6644
rect 1581 6607 1639 6613
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3418 6644 3424 6656
rect 3283 6616 3424 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3418 6604 3424 6616
rect 3476 6644 3482 6656
rect 3697 6647 3755 6653
rect 3697 6644 3709 6647
rect 3476 6616 3709 6644
rect 3476 6604 3482 6616
rect 3697 6613 3709 6616
rect 3743 6613 3755 6647
rect 3697 6607 3755 6613
rect 7561 6647 7619 6653
rect 7561 6613 7573 6647
rect 7607 6644 7619 6647
rect 7742 6644 7748 6656
rect 7607 6616 7748 6644
rect 7607 6613 7619 6616
rect 7561 6607 7619 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 11054 6644 11060 6656
rect 11015 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11974 6644 11980 6656
rect 11935 6616 11980 6644
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13630 6644 13636 6656
rect 12860 6616 13636 6644
rect 12860 6604 12866 6616
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 2096 6412 4261 6440
rect 2096 6400 2102 6412
rect 4249 6409 4261 6412
rect 4295 6440 4307 6443
rect 5074 6440 5080 6452
rect 4295 6412 5080 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5442 6440 5448 6452
rect 5403 6412 5448 6440
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 6730 6440 6736 6452
rect 5951 6412 6736 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 8662 6440 8668 6452
rect 8623 6412 8668 6440
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9950 6440 9956 6452
rect 9815 6412 9956 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 3329 6375 3387 6381
rect 3329 6372 3341 6375
rect 2669 6344 3341 6372
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1544 6276 1593 6304
rect 1544 6264 1550 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2406 6236 2412 6248
rect 1443 6208 2412 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2669 6245 2697 6344
rect 3329 6341 3341 6344
rect 3375 6372 3387 6375
rect 5258 6372 5264 6384
rect 3375 6344 5264 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 6457 6375 6515 6381
rect 6457 6372 6469 6375
rect 5592 6344 6469 6372
rect 5592 6332 5598 6344
rect 6457 6341 6469 6344
rect 6503 6372 6515 6375
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 6503 6344 6561 6372
rect 6503 6341 6515 6344
rect 6457 6335 6515 6341
rect 6549 6341 6561 6344
rect 6595 6341 6607 6375
rect 6549 6335 6607 6341
rect 8573 6375 8631 6381
rect 8573 6341 8585 6375
rect 8619 6372 8631 6375
rect 8754 6372 8760 6384
rect 8619 6344 8760 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 8754 6332 8760 6344
rect 8812 6372 8818 6384
rect 8812 6344 9168 6372
rect 8812 6332 8818 6344
rect 4890 6304 4896 6316
rect 4851 6276 4896 6304
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7558 6304 7564 6316
rect 6319 6276 7564 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7558 6264 7564 6276
rect 7616 6304 7622 6316
rect 9140 6313 9168 6344
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7616 6276 7665 6304
rect 7616 6264 7622 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9784 6304 9812 6403
rect 9950 6400 9956 6412
rect 10008 6440 10014 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 10008 6412 10057 6440
rect 10008 6400 10014 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11296 6412 11805 6440
rect 11296 6400 11302 6412
rect 11793 6409 11805 6412
rect 11839 6440 11851 6443
rect 11839 6412 12940 6440
rect 11839 6409 11851 6412
rect 11793 6403 11851 6409
rect 12912 6313 12940 6412
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 13412 6412 13461 6440
rect 13412 6400 13418 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 9355 6276 9812 6304
rect 12897 6307 12955 6313
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 12897 6273 12909 6307
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 2669 6239 2731 6245
rect 2669 6208 2685 6239
rect 2673 6205 2685 6208
rect 2719 6205 2731 6239
rect 2673 6199 2731 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 3927 6208 4813 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4801 6205 4813 6208
rect 4847 6236 4859 6239
rect 5166 6236 5172 6248
rect 4847 6208 5172 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6236 6515 6239
rect 7466 6236 7472 6248
rect 6503 6208 7472 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7892 6208 8125 6236
rect 7892 6196 7898 6208
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8478 6236 8484 6248
rect 8159 6208 8484 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8478 6196 8484 6208
rect 8536 6236 8542 6248
rect 9490 6236 9496 6248
rect 8536 6208 9496 6236
rect 8536 6196 8542 6208
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 10226 6236 10232 6248
rect 10187 6208 10232 6236
rect 10226 6196 10232 6208
rect 10284 6236 10290 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10284 6208 10793 6236
rect 10284 6196 10290 6208
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12526 6236 12532 6248
rect 12299 6208 12532 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13004 6236 13032 6267
rect 12860 6208 13032 6236
rect 12860 6196 12866 6208
rect 1578 6128 1584 6180
rect 1636 6168 1642 6180
rect 2225 6171 2283 6177
rect 2225 6168 2237 6171
rect 1636 6140 2237 6168
rect 1636 6128 1642 6140
rect 2225 6137 2237 6140
rect 2271 6168 2283 6171
rect 2314 6168 2320 6180
rect 2271 6140 2320 6168
rect 2271 6137 2283 6140
rect 2225 6131 2283 6137
rect 2314 6128 2320 6140
rect 2372 6168 2378 6180
rect 4709 6171 4767 6177
rect 2372 6140 4660 6168
rect 2372 6128 2378 6140
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 2464 6072 2513 6100
rect 2464 6060 2470 6072
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 2501 6063 2559 6069
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2648 6072 2881 6100
rect 2648 6060 2654 6072
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 4338 6100 4344 6112
rect 4299 6072 4344 6100
rect 2869 6063 2927 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 4632 6100 4660 6140
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 4982 6168 4988 6180
rect 4755 6140 4988 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 7561 6171 7619 6177
rect 7561 6168 7573 6171
rect 5184 6140 7573 6168
rect 5184 6100 5212 6140
rect 7561 6137 7573 6140
rect 7607 6168 7619 6171
rect 7742 6168 7748 6180
rect 7607 6140 7748 6168
rect 7607 6137 7619 6140
rect 7561 6131 7619 6137
rect 7742 6128 7748 6140
rect 7800 6168 7806 6180
rect 9033 6171 9091 6177
rect 9033 6168 9045 6171
rect 7800 6140 9045 6168
rect 7800 6128 7806 6140
rect 9033 6137 9045 6140
rect 9079 6168 9091 6171
rect 9306 6168 9312 6180
rect 9079 6140 9312 6168
rect 9079 6137 9091 6140
rect 9033 6131 9091 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9582 6128 9588 6180
rect 9640 6168 9646 6180
rect 11054 6168 11060 6180
rect 9640 6140 11060 6168
rect 9640 6128 9646 6140
rect 11054 6128 11060 6140
rect 11112 6168 11118 6180
rect 11149 6171 11207 6177
rect 11149 6168 11161 6171
rect 11112 6140 11161 6168
rect 11112 6128 11118 6140
rect 11149 6137 11161 6140
rect 11195 6137 11207 6171
rect 12618 6168 12624 6180
rect 11149 6131 11207 6137
rect 12452 6140 12624 6168
rect 7098 6100 7104 6112
rect 4632 6072 5212 6100
rect 7059 6072 7104 6100
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 9732 6072 10425 6100
rect 9732 6060 9738 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 11330 6100 11336 6112
rect 11291 6072 11336 6100
rect 10413 6063 10471 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 12452 6109 12480 6140
rect 12618 6128 12624 6140
rect 12676 6168 12682 6180
rect 13817 6171 13875 6177
rect 13817 6168 13829 6171
rect 12676 6140 13829 6168
rect 12676 6128 12682 6140
rect 13817 6137 13829 6140
rect 13863 6137 13875 6171
rect 13817 6131 13875 6137
rect 12437 6103 12495 6109
rect 12437 6069 12449 6103
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12584 6072 12817 6100
rect 12584 6060 12590 6072
rect 12805 6069 12817 6072
rect 12851 6100 12863 6103
rect 13354 6100 13360 6112
rect 12851 6072 13360 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 3329 5899 3387 5905
rect 3329 5896 3341 5899
rect 2832 5868 3341 5896
rect 2832 5856 2838 5868
rect 3329 5865 3341 5868
rect 3375 5896 3387 5899
rect 4338 5896 4344 5908
rect 3375 5868 4344 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 4614 5896 4620 5908
rect 4575 5868 4620 5896
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 6549 5899 6607 5905
rect 5316 5868 6224 5896
rect 5316 5856 5322 5868
rect 2958 5828 2964 5840
rect 1412 5800 2964 5828
rect 1412 5769 1440 5800
rect 2958 5788 2964 5800
rect 3016 5828 3022 5840
rect 3605 5831 3663 5837
rect 3605 5828 3617 5831
rect 3016 5800 3617 5828
rect 3016 5788 3022 5800
rect 3605 5797 3617 5800
rect 3651 5797 3663 5831
rect 6086 5828 6092 5840
rect 3605 5791 3663 5797
rect 5552 5800 6092 5828
rect 5552 5772 5580 5800
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 6196 5828 6224 5868
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 6638 5896 6644 5908
rect 6595 5868 6644 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6972 5868 7205 5896
rect 6972 5856 6978 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 8386 5896 8392 5908
rect 8159 5868 8392 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 8128 5828 8156 5859
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9306 5896 9312 5908
rect 8987 5868 9312 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11388 5868 12081 5896
rect 11388 5856 11394 5868
rect 12069 5865 12081 5868
rect 12115 5896 12127 5899
rect 12158 5896 12164 5908
rect 12115 5868 12164 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 6196 5800 8156 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 2866 5760 2872 5772
rect 2731 5732 2872 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 4062 5760 4068 5772
rect 4023 5732 4068 5760
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 5534 5760 5540 5772
rect 5495 5732 5540 5760
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5902 5760 5908 5772
rect 5675 5732 5908 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 7098 5760 7104 5772
rect 7059 5732 7104 5760
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8386 5760 8392 5772
rect 8343 5732 8392 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8386 5720 8392 5732
rect 8444 5760 8450 5772
rect 8846 5760 8852 5772
rect 8444 5732 8852 5760
rect 8444 5720 8450 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9766 5760 9772 5772
rect 9723 5732 9772 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 13262 5760 13268 5772
rect 12176 5732 13268 5760
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5661 5779 5695
rect 7282 5692 7288 5704
rect 7243 5664 7288 5692
rect 5721 5655 5779 5661
rect 2501 5627 2559 5633
rect 2501 5593 2513 5627
rect 2547 5624 2559 5627
rect 3142 5624 3148 5636
rect 2547 5596 3148 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 5074 5584 5080 5636
rect 5132 5624 5138 5636
rect 5736 5624 5764 5655
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12176 5701 12204 5732
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11848 5664 12173 5692
rect 11848 5652 11854 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12802 5692 12808 5704
rect 12299 5664 12808 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 5132 5596 5764 5624
rect 9861 5627 9919 5633
rect 5132 5584 5138 5596
rect 9861 5593 9873 5627
rect 9907 5624 9919 5627
rect 10042 5624 10048 5636
rect 9907 5596 10048 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 10321 5627 10379 5633
rect 10321 5593 10333 5627
rect 10367 5624 10379 5627
rect 11701 5627 11759 5633
rect 10367 5596 11376 5624
rect 10367 5593 10379 5596
rect 10321 5587 10379 5593
rect 11348 5568 11376 5596
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 11974 5624 11980 5636
rect 11747 5596 11980 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 2130 5516 2136 5568
rect 2188 5556 2194 5568
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2188 5528 2881 5556
rect 2188 5516 2194 5528
rect 2869 5525 2881 5528
rect 2915 5525 2927 5559
rect 4246 5556 4252 5568
rect 4207 5528 4252 5556
rect 2869 5519 2927 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4982 5556 4988 5568
rect 4943 5528 4988 5556
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 6730 5556 6736 5568
rect 6691 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 10594 5556 10600 5568
rect 10555 5528 10600 5556
rect 10594 5516 10600 5528
rect 10652 5516 10658 5568
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 12268 5556 12296 5655
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 11388 5528 12296 5556
rect 11388 5516 11394 5528
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 13449 5559 13507 5565
rect 13449 5556 13461 5559
rect 12860 5528 13461 5556
rect 12860 5516 12866 5528
rect 13449 5525 13461 5528
rect 13495 5525 13507 5559
rect 13449 5519 13507 5525
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 1946 5352 1952 5364
rect 1907 5324 1952 5352
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 2961 5355 3019 5361
rect 2961 5352 2973 5355
rect 2924 5324 2973 5352
rect 2924 5312 2930 5324
rect 2961 5321 2973 5324
rect 3007 5321 3019 5355
rect 4890 5352 4896 5364
rect 4851 5324 4896 5352
rect 2961 5315 3019 5321
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9398 5352 9404 5364
rect 9263 5324 9404 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 1857 5287 1915 5293
rect 1857 5253 1869 5287
rect 1903 5284 1915 5287
rect 5902 5284 5908 5296
rect 1903 5256 2636 5284
rect 5863 5256 5908 5284
rect 1903 5253 1915 5256
rect 1857 5247 1915 5253
rect 2406 5216 2412 5228
rect 2367 5188 2412 5216
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2608 5225 2636 5256
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5216 2651 5219
rect 3050 5216 3056 5228
rect 2639 5188 3056 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3476 5188 3525 5216
rect 3476 5176 3482 5188
rect 3513 5185 3525 5188
rect 3559 5185 3571 5219
rect 7282 5216 7288 5228
rect 3513 5179 3571 5185
rect 6564 5188 7288 5216
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2682 5148 2688 5160
rect 2363 5120 2688 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 5534 5148 5540 5160
rect 5495 5120 5540 5148
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 3421 5083 3479 5089
rect 3421 5049 3433 5083
rect 3467 5080 3479 5083
rect 3758 5083 3816 5089
rect 3758 5080 3770 5083
rect 3467 5052 3770 5080
rect 3467 5049 3479 5052
rect 3421 5043 3479 5049
rect 3758 5049 3770 5052
rect 3804 5080 3816 5083
rect 5074 5080 5080 5092
rect 3804 5052 5080 5080
rect 3804 5049 3816 5052
rect 3758 5043 3816 5049
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 6564 5021 6592 5188
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 7340 5188 7573 5216
rect 7340 5176 7346 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 9232 5148 9260 5315
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9640 5324 9689 5352
rect 9640 5312 9646 5324
rect 9677 5321 9689 5324
rect 9723 5352 9735 5355
rect 9766 5352 9772 5364
rect 9723 5324 9772 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12158 5352 12164 5364
rect 12119 5324 12164 5352
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 12894 5312 12900 5364
rect 12952 5352 12958 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12952 5324 13001 5352
rect 12952 5312 12958 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 13320 5324 13369 5352
rect 13320 5312 13326 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 13357 5315 13415 5321
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11330 5216 11336 5228
rect 10827 5188 11336 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 8619 5120 9260 5148
rect 12437 5151 12495 5157
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12894 5148 12900 5160
rect 12483 5120 12900 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12894 5108 12900 5120
rect 12952 5108 12958 5160
rect 7377 5083 7435 5089
rect 7377 5049 7389 5083
rect 7423 5080 7435 5083
rect 7558 5080 7564 5092
rect 7423 5052 7564 5080
rect 7423 5049 7435 5052
rect 7377 5043 7435 5049
rect 7558 5040 7564 5052
rect 7616 5040 7622 5092
rect 10045 5083 10103 5089
rect 10045 5049 10057 5083
rect 10091 5080 10103 5083
rect 10091 5052 10548 5080
rect 10091 5049 10103 5052
rect 10045 5043 10103 5049
rect 10520 5024 10548 5052
rect 6273 5015 6331 5021
rect 6273 4981 6285 5015
rect 6319 5012 6331 5015
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6319 4984 6561 5012
rect 6319 4981 6331 4984
rect 6273 4975 6331 4981
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 6549 4975 6607 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7466 5012 7472 5024
rect 7427 4984 7472 5012
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 8754 5012 8760 5024
rect 8715 4984 8760 5012
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 10134 5012 10140 5024
rect 10095 4984 10140 5012
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10502 5012 10508 5024
rect 10463 4984 10508 5012
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 11330 5012 11336 5024
rect 10652 4984 10697 5012
rect 11291 4984 11336 5012
rect 10652 4972 10658 4984
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4212 4780 4261 4808
rect 4212 4768 4218 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 4433 4811 4491 4817
rect 4433 4777 4445 4811
rect 4479 4808 4491 4811
rect 4982 4808 4988 4820
rect 4479 4780 4988 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5994 4808 6000 4820
rect 5955 4780 6000 4808
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 6730 4808 6736 4820
rect 6503 4780 6736 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6972 4780 7021 4808
rect 6972 4768 6978 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 7469 4811 7527 4817
rect 7469 4777 7481 4811
rect 7515 4808 7527 4811
rect 7650 4808 7656 4820
rect 7515 4780 7656 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 7650 4768 7656 4780
rect 7708 4808 7714 4820
rect 8110 4808 8116 4820
rect 7708 4780 8116 4808
rect 7708 4768 7714 4780
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10192 4780 10701 4808
rect 10192 4768 10198 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 11054 4808 11060 4820
rect 11015 4780 11060 4808
rect 10689 4771 10747 4777
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 2498 4740 2504 4752
rect 2363 4712 2504 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 2498 4700 2504 4712
rect 2556 4700 2562 4752
rect 4890 4740 4896 4752
rect 4803 4712 4896 4740
rect 4890 4700 4896 4712
rect 4948 4740 4954 4752
rect 5442 4740 5448 4752
rect 4948 4712 5448 4740
rect 4948 4700 4954 4712
rect 5442 4700 5448 4712
rect 5500 4700 5506 4752
rect 5905 4743 5963 4749
rect 5905 4709 5917 4743
rect 5951 4740 5963 4743
rect 7098 4740 7104 4752
rect 5951 4712 7104 4740
rect 5951 4709 5963 4712
rect 5905 4703 5963 4709
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 8021 4743 8079 4749
rect 8021 4709 8033 4743
rect 8067 4740 8079 4743
rect 8386 4740 8392 4752
rect 8067 4712 8392 4740
rect 8067 4709 8079 4712
rect 8021 4703 8079 4709
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 3142 4672 3148 4684
rect 2823 4644 3148 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 4798 4672 4804 4684
rect 4759 4644 4804 4672
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5776 4644 6377 4672
rect 5776 4632 5782 4644
rect 6365 4641 6377 4644
rect 6411 4672 6423 4675
rect 7006 4672 7012 4684
rect 6411 4644 7012 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 8202 4672 8208 4684
rect 7975 4644 8208 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 10042 4672 10048 4684
rect 9539 4644 10048 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 11330 4672 11336 4684
rect 10336 4644 11336 4672
rect 10336 4616 10364 4644
rect 11330 4632 11336 4644
rect 11388 4672 11394 4684
rect 11497 4675 11555 4681
rect 11497 4672 11509 4675
rect 11388 4644 11509 4672
rect 11388 4632 11394 4644
rect 11497 4641 11509 4644
rect 11543 4641 11555 4675
rect 11497 4635 11555 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2866 4604 2872 4616
rect 1995 4576 2872 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 2961 4567 3019 4573
rect 2498 4496 2504 4548
rect 2556 4536 2562 4548
rect 2976 4536 3004 4567
rect 5074 4564 5080 4576
rect 5132 4604 5138 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5132 4576 5457 4604
rect 5132 4564 5138 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 5445 4567 5503 4573
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8168 4576 8213 4604
rect 8168 4564 8174 4576
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9732 4576 10149 4604
rect 9732 4564 9738 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10318 4604 10324 4616
rect 10231 4576 10324 4604
rect 10137 4567 10195 4573
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11112 4576 11253 4604
rect 11112 4564 11118 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 7558 4536 7564 4548
rect 2556 4508 3004 4536
rect 7471 4508 7564 4536
rect 2556 4496 2562 4508
rect 7558 4496 7564 4508
rect 7616 4536 7622 4548
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 7616 4508 8953 4536
rect 7616 4496 7622 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 3510 4468 3516 4480
rect 3471 4440 3516 4468
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4062 4468 4068 4480
rect 3927 4440 4068 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8573 4471 8631 4477
rect 8573 4468 8585 4471
rect 7524 4440 8585 4468
rect 7524 4428 7530 4440
rect 8573 4437 8585 4440
rect 8619 4437 8631 4471
rect 8573 4431 8631 4437
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 10502 4468 10508 4480
rect 9723 4440 10508 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 10502 4428 10508 4440
rect 10560 4428 10566 4480
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 12621 4471 12679 4477
rect 12621 4468 12633 4471
rect 10744 4440 12633 4468
rect 10744 4428 10750 4440
rect 12621 4437 12633 4440
rect 12667 4468 12679 4471
rect 12710 4468 12716 4480
rect 12667 4440 12716 4468
rect 12667 4437 12679 4440
rect 12621 4431 12679 4437
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2314 4264 2320 4276
rect 2275 4236 2320 4264
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 2924 4236 4353 4264
rect 2924 4224 2930 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 5074 4224 5080 4276
rect 5132 4264 5138 4276
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 5132 4236 5365 4264
rect 5132 4224 5138 4236
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 5353 4227 5411 4233
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 6546 4264 6552 4276
rect 6135 4236 6552 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 7466 4264 7472 4276
rect 7427 4236 7472 4264
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 9769 4267 9827 4273
rect 9769 4233 9781 4267
rect 9815 4264 9827 4267
rect 10318 4264 10324 4276
rect 9815 4236 10324 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 11609 4267 11667 4273
rect 11609 4264 11621 4267
rect 11112 4236 11621 4264
rect 11112 4224 11118 4236
rect 11609 4233 11621 4236
rect 11655 4264 11667 4267
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11655 4236 11989 4264
rect 11655 4233 11667 4236
rect 11609 4227 11667 4233
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 11977 4227 12035 4233
rect 2777 4199 2835 4205
rect 2777 4165 2789 4199
rect 2823 4196 2835 4199
rect 3510 4196 3516 4208
rect 2823 4168 3516 4196
rect 2823 4165 2835 4168
rect 2777 4159 2835 4165
rect 3510 4156 3516 4168
rect 3568 4156 3574 4208
rect 3602 4156 3608 4208
rect 3660 4196 3666 4208
rect 4062 4196 4068 4208
rect 3660 4168 4068 4196
rect 3660 4156 3666 4168
rect 4062 4156 4068 4168
rect 4120 4156 4126 4208
rect 4249 4199 4307 4205
rect 4249 4165 4261 4199
rect 4295 4196 4307 4199
rect 4890 4196 4896 4208
rect 4295 4168 4896 4196
rect 4295 4165 4307 4168
rect 4249 4159 4307 4165
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3108 4100 3341 4128
rect 3108 4088 3114 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 4080 4128 4108 4156
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4080 4100 4813 4128
rect 3329 4091 3387 4097
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5092 4128 5120 4224
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 8110 4196 8116 4208
rect 6972 4168 8116 4196
rect 6972 4156 6978 4168
rect 8036 4137 8064 4168
rect 8110 4156 8116 4168
rect 8168 4196 8174 4208
rect 8168 4168 8248 4196
rect 8168 4156 8174 4168
rect 5031 4100 5120 4128
rect 8021 4131 8079 4137
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 8021 4097 8033 4131
rect 8067 4097 8079 4131
rect 8220 4128 8248 4168
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 8220 4100 8861 4128
rect 8021 4091 8079 4097
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 10502 4128 10508 4140
rect 10463 4100 10508 4128
rect 8849 4091 8907 4097
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10686 4128 10692 4140
rect 10647 4100 10692 4128
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 12986 4128 12992 4140
rect 12452 4100 12992 4128
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1946 4060 1952 4072
rect 1443 4032 1952 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 3568 4032 4721 4060
rect 3568 4020 3574 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4060 7435 4063
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7423 4032 7849 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 7837 4029 7849 4032
rect 7883 4060 7895 4063
rect 8478 4060 8484 4072
rect 7883 4032 8484 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 9030 4060 9036 4072
rect 8991 4032 9036 4060
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 12452 4069 12480 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10192 4032 10425 4060
rect 10192 4020 10198 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 1670 3992 1676 4004
rect 1631 3964 1676 3992
rect 1670 3952 1676 3964
rect 1728 3952 1734 4004
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 3145 3995 3203 4001
rect 3145 3992 3157 3995
rect 2372 3964 3157 3992
rect 2372 3952 2378 3964
rect 3145 3961 3157 3964
rect 3191 3961 3203 3995
rect 3878 3992 3884 4004
rect 3839 3964 3884 3992
rect 3145 3955 3203 3961
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 7929 3995 7987 4001
rect 7929 3992 7941 3995
rect 6564 3964 7941 3992
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 3237 3927 3295 3933
rect 3237 3924 3249 3927
rect 2731 3896 3249 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 3237 3893 3249 3896
rect 3283 3924 3295 3927
rect 3326 3924 3332 3936
rect 3283 3896 3332 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6564 3933 6592 3964
rect 7929 3961 7941 3964
rect 7975 3961 7987 3995
rect 7929 3955 7987 3961
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 8573 3995 8631 4001
rect 8573 3992 8585 3995
rect 8444 3964 8585 3992
rect 8444 3952 8450 3964
rect 8573 3961 8585 3964
rect 8619 3992 8631 3995
rect 9582 3992 9588 4004
rect 8619 3964 9588 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 9582 3952 9588 3964
rect 9640 3952 9646 4004
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6144 3896 6561 3924
rect 6144 3884 6150 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10410 3924 10416 3936
rect 10091 3896 10416 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 11330 3924 11336 3936
rect 11291 3896 11336 3924
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 12618 3924 12624 3936
rect 12579 3896 12624 3924
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 3602 3720 3608 3732
rect 2455 3692 3608 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 4120 3692 4537 3720
rect 4120 3680 4126 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 5074 3720 5080 3732
rect 5035 3692 5080 3720
rect 4525 3683 4583 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6089 3723 6147 3729
rect 6089 3689 6101 3723
rect 6135 3720 6147 3723
rect 6730 3720 6736 3732
rect 6135 3692 6736 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7340 3692 7665 3720
rect 7340 3680 7346 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 10560 3692 10609 3720
rect 10560 3680 10566 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 10597 3683 10655 3689
rect 10686 3680 10692 3732
rect 10744 3680 10750 3732
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 11388 3692 12449 3720
rect 11388 3680 11394 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 12437 3683 12495 3689
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 1302 3652 1308 3664
rect 624 3624 1308 3652
rect 624 3612 630 3624
rect 1302 3612 1308 3624
rect 1360 3612 1366 3664
rect 1673 3655 1731 3661
rect 1673 3621 1685 3655
rect 1719 3652 1731 3655
rect 2774 3652 2780 3664
rect 1719 3624 2780 3652
rect 1719 3621 1731 3624
rect 1673 3615 1731 3621
rect 2774 3612 2780 3624
rect 2832 3652 2838 3664
rect 5810 3652 5816 3664
rect 2832 3624 5816 3652
rect 2832 3612 2838 3624
rect 5810 3612 5816 3624
rect 5868 3612 5874 3664
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 6540 3655 6598 3661
rect 6540 3652 6552 3655
rect 6420 3624 6552 3652
rect 6420 3612 6426 3624
rect 6540 3621 6552 3624
rect 6586 3652 6598 3655
rect 6914 3652 6920 3664
rect 6586 3624 6920 3652
rect 6586 3621 6598 3624
rect 6540 3615 6598 3621
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 10321 3655 10379 3661
rect 10321 3621 10333 3655
rect 10367 3652 10379 3655
rect 10704 3652 10732 3680
rect 10367 3624 10732 3652
rect 10367 3621 10379 3624
rect 10321 3615 10379 3621
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 3568 3556 4445 3584
rect 3568 3544 3574 3556
rect 4433 3553 4445 3556
rect 4479 3584 4491 3587
rect 5258 3584 5264 3596
rect 4479 3556 5264 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9640 3556 9689 3584
rect 9640 3544 9646 3556
rect 9677 3553 9689 3556
rect 9723 3584 9735 3587
rect 10226 3584 10232 3596
rect 9723 3556 10232 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 11054 3584 11060 3596
rect 11015 3556 11060 3584
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11313 3587 11371 3593
rect 11313 3584 11325 3587
rect 11204 3556 11325 3584
rect 11204 3544 11210 3556
rect 11313 3553 11325 3556
rect 11359 3553 11371 3587
rect 11313 3547 11371 3553
rect 12526 3544 12532 3596
rect 12584 3584 12590 3596
rect 13170 3584 13176 3596
rect 12584 3556 13176 3584
rect 12584 3544 12590 3556
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3050 3516 3056 3528
rect 2963 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3516 3114 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3108 3488 3433 3516
rect 3108 3476 3114 3488
rect 3421 3485 3433 3488
rect 3467 3516 3479 3519
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3467 3488 3893 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3881 3485 3893 3488
rect 3927 3516 3939 3519
rect 4614 3516 4620 3528
rect 3927 3488 4620 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 6270 3516 6276 3528
rect 6231 3488 6276 3516
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 12768 3488 13553 3516
rect 12768 3476 12774 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 1854 3408 1860 3460
rect 1912 3448 1918 3460
rect 2590 3448 2596 3460
rect 1912 3420 2596 3448
rect 1912 3408 1918 3420
rect 2590 3408 2596 3420
rect 2648 3408 2654 3460
rect 8294 3448 8300 3460
rect 8207 3420 8300 3448
rect 8294 3408 8300 3420
rect 8352 3448 8358 3460
rect 9398 3448 9404 3460
rect 8352 3420 9404 3448
rect 8352 3408 8358 3420
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 10226 3448 10232 3460
rect 9824 3420 10232 3448
rect 9824 3408 9830 3420
rect 10226 3408 10232 3420
rect 10284 3408 10290 3460
rect 2317 3383 2375 3389
rect 2317 3349 2329 3383
rect 2363 3380 2375 3383
rect 3050 3380 3056 3392
rect 2363 3352 3056 3380
rect 2363 3349 2375 3352
rect 2317 3343 2375 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 4065 3383 4123 3389
rect 4065 3349 4077 3383
rect 4111 3380 4123 3383
rect 4246 3380 4252 3392
rect 4111 3352 4252 3380
rect 4111 3349 4123 3352
rect 4065 3343 4123 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 8536 3352 8585 3380
rect 8536 3340 8542 3352
rect 8573 3349 8585 3352
rect 8619 3380 8631 3383
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8619 3352 8953 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 8941 3343 8999 3349
rect 9861 3383 9919 3389
rect 9861 3349 9873 3383
rect 9907 3380 9919 3383
rect 10134 3380 10140 3392
rect 9907 3352 10140 3380
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2866 3176 2872 3188
rect 2547 3148 2872 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 5442 3176 5448 3188
rect 5132 3148 5448 3176
rect 5132 3136 5138 3148
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3176 7159 3179
rect 7190 3176 7196 3188
rect 7147 3148 7196 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8570 3136 8576 3148
rect 8628 3176 8634 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 8628 3148 9137 3176
rect 8628 3136 8634 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9582 3176 9588 3188
rect 9543 3148 9588 3176
rect 9125 3139 9183 3145
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 3145 3111 3203 3117
rect 3145 3108 3157 3111
rect 2648 3080 3157 3108
rect 2648 3068 2654 3080
rect 3145 3077 3157 3080
rect 3191 3077 3203 3111
rect 3145 3071 3203 3077
rect 3234 3068 3240 3120
rect 3292 3108 3298 3120
rect 3881 3111 3939 3117
rect 3881 3108 3893 3111
rect 3292 3080 3893 3108
rect 3292 3068 3298 3080
rect 3881 3077 3893 3080
rect 3927 3108 3939 3111
rect 4062 3108 4068 3120
rect 3927 3080 4068 3108
rect 3927 3077 3939 3080
rect 3881 3071 3939 3077
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 2774 3040 2780 3052
rect 1688 3012 2780 3040
rect 1422 2975 1480 2981
rect 1422 2941 1434 2975
rect 1468 2972 1480 2975
rect 1688 2972 1716 3012
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 9140 3040 9168 3139
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11480 3148 11805 3176
rect 11480 3136 11486 3148
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 12434 3176 12440 3188
rect 12395 3148 12440 3176
rect 11793 3139 11851 3145
rect 11057 3111 11115 3117
rect 11057 3077 11069 3111
rect 11103 3108 11115 3111
rect 11146 3108 11152 3120
rect 11103 3080 11152 3108
rect 11103 3077 11115 3080
rect 11057 3071 11115 3077
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 11808 3108 11836 3139
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 12710 3108 12716 3120
rect 11808 3080 12716 3108
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 13081 3043 13139 3049
rect 3476 3012 4108 3040
rect 9140 3012 9812 3040
rect 3476 3000 3482 3012
rect 1468 2944 1716 2972
rect 2961 2975 3019 2981
rect 1468 2941 1480 2944
rect 1422 2935 1480 2941
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3970 2972 3976 2984
rect 3007 2944 3976 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 4080 2981 4108 3012
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2972 4123 2975
rect 6270 2972 6276 2984
rect 4111 2944 6276 2972
rect 4111 2941 4123 2944
rect 4065 2935 4123 2941
rect 6270 2932 6276 2944
rect 6328 2972 6334 2984
rect 7190 2972 7196 2984
rect 6328 2944 7196 2972
rect 6328 2932 6334 2944
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7282 2932 7288 2984
rect 7340 2972 7346 2984
rect 7449 2975 7507 2981
rect 7449 2972 7461 2975
rect 7340 2944 7461 2972
rect 7340 2932 7346 2944
rect 7449 2941 7461 2944
rect 7495 2941 7507 2975
rect 7449 2935 7507 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2941 9735 2975
rect 9784 2972 9812 3012
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13446 3040 13452 3052
rect 13127 3012 13452 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14918 3040 14924 3052
rect 13872 3012 14924 3040
rect 13872 3000 13878 3012
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 9933 2975 9991 2981
rect 9933 2972 9945 2975
rect 9784 2944 9945 2972
rect 9677 2935 9735 2941
rect 9933 2941 9945 2944
rect 9979 2941 9991 2975
rect 9933 2935 9991 2941
rect 4332 2907 4390 2913
rect 4332 2873 4344 2907
rect 4378 2904 4390 2907
rect 4614 2904 4620 2916
rect 4378 2876 4620 2904
rect 4378 2873 4390 2876
rect 4332 2867 4390 2873
rect 4614 2864 4620 2876
rect 4672 2904 4678 2916
rect 5074 2904 5080 2916
rect 4672 2876 5080 2904
rect 4672 2864 4678 2876
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 9692 2904 9720 2935
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12768 2944 12817 2972
rect 12768 2932 12774 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 13722 2972 13728 2984
rect 12943 2944 13728 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 11054 2904 11060 2916
rect 9692 2876 11060 2904
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 11422 2864 11428 2916
rect 11480 2904 11486 2916
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 11480 2876 12265 2904
rect 11480 2864 11486 2876
rect 12253 2873 12265 2876
rect 12299 2904 12311 2907
rect 12912 2904 12940 2935
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 12299 2876 12940 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 256 2808 1593 2836
rect 256 2796 262 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 1949 2839 2007 2845
rect 1949 2836 1961 2839
rect 1820 2808 1961 2836
rect 1820 2796 1826 2808
rect 1949 2805 1961 2808
rect 1995 2805 2007 2839
rect 13446 2836 13452 2848
rect 13407 2808 13452 2836
rect 1949 2799 2007 2805
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3050 2632 3056 2644
rect 2915 2604 3056 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3970 2632 3976 2644
rect 3559 2604 3976 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4080 2604 4445 2632
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4080 2564 4108 2604
rect 4433 2601 4445 2604
rect 4479 2632 4491 2635
rect 4706 2632 4712 2644
rect 4479 2604 4712 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5074 2632 5080 2644
rect 5035 2604 5080 2632
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5442 2632 5448 2644
rect 5403 2604 5448 2632
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7190 2632 7196 2644
rect 7103 2604 7196 2632
rect 7190 2592 7196 2604
rect 7248 2632 7254 2644
rect 8478 2632 8484 2644
rect 7248 2604 8484 2632
rect 7248 2592 7254 2604
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 8570 2592 8576 2644
rect 8628 2592 8634 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 9732 2604 10241 2632
rect 9732 2592 9738 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 10229 2595 10287 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 3927 2536 4108 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4246 2524 4252 2576
rect 4304 2564 4310 2576
rect 4525 2567 4583 2573
rect 4525 2564 4537 2567
rect 4304 2536 4537 2564
rect 4304 2524 4310 2536
rect 4525 2533 4537 2536
rect 4571 2564 4583 2567
rect 6549 2567 6607 2573
rect 6549 2564 6561 2567
rect 4571 2536 6561 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 6549 2533 6561 2536
rect 6595 2533 6607 2567
rect 8588 2564 8616 2592
rect 9490 2564 9496 2576
rect 8588 2536 9496 2564
rect 6549 2527 6607 2533
rect 9490 2524 9496 2536
rect 9548 2564 9554 2576
rect 10134 2564 10140 2576
rect 9548 2536 10140 2564
rect 9548 2524 9554 2536
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 10778 2524 10784 2576
rect 10836 2564 10842 2576
rect 12158 2564 12164 2576
rect 10836 2536 12164 2564
rect 10836 2524 10842 2536
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 12452 2564 12480 2592
rect 13081 2567 13139 2573
rect 13081 2564 13093 2567
rect 12452 2536 13093 2564
rect 13081 2533 13093 2536
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 1762 2505 1768 2508
rect 1745 2499 1768 2505
rect 1745 2496 1757 2499
rect 1452 2468 1757 2496
rect 1452 2456 1458 2468
rect 1745 2465 1757 2468
rect 1820 2496 1826 2508
rect 5629 2499 5687 2505
rect 1820 2468 1893 2496
rect 1745 2459 1768 2465
rect 1762 2456 1768 2459
rect 1820 2456 1826 2468
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 7469 2499 7527 2505
rect 5675 2468 6316 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2397 1547 2431
rect 1489 2391 1547 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5442 2428 5448 2440
rect 4755 2400 5448 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 1504 2292 1532 2391
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 6288 2372 6316 2468
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 8018 2496 8024 2508
rect 7515 2468 8024 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 9585 2499 9643 2505
rect 8619 2468 9260 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9232 2437 9260 2468
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9766 2496 9772 2508
rect 9631 2468 9772 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 9824 2468 10609 2496
rect 9824 2456 9830 2468
rect 10597 2465 10609 2468
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11940 2468 11989 2496
rect 11940 2456 11946 2468
rect 11977 2465 11989 2468
rect 12023 2496 12035 2499
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12023 2468 13001 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9950 2428 9956 2440
rect 9263 2400 9956 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10134 2428 10140 2440
rect 10047 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2428 10198 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10192 2400 10701 2428
rect 10192 2388 10198 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11146 2428 11152 2440
rect 10919 2400 11152 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 11146 2388 11152 2400
rect 11204 2428 11210 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11204 2400 11345 2428
rect 11204 2388 11210 2400
rect 11333 2397 11345 2400
rect 11379 2428 11391 2431
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11379 2400 11713 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 11701 2397 11713 2400
rect 11747 2428 11759 2431
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 11747 2400 13277 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 13265 2397 13277 2400
rect 13311 2428 13323 2431
rect 13446 2428 13452 2440
rect 13311 2400 13452 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13446 2388 13452 2400
rect 13504 2428 13510 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13504 2400 13645 2428
rect 13504 2388 13510 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 3142 2320 3148 2372
rect 3200 2360 3206 2372
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 3200 2332 4077 2360
rect 3200 2320 3206 2332
rect 4065 2329 4077 2332
rect 4111 2329 4123 2363
rect 6270 2360 6276 2372
rect 6231 2332 6276 2360
rect 4065 2323 4123 2329
rect 6270 2320 6276 2332
rect 6328 2320 6334 2372
rect 9766 2320 9772 2372
rect 9824 2360 9830 2372
rect 10226 2360 10232 2372
rect 9824 2332 10232 2360
rect 9824 2320 9830 2332
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 3418 2292 3424 2304
rect 1504 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 5810 2292 5816 2304
rect 5771 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 7650 2292 7656 2304
rect 7611 2264 7656 2292
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 5718 1232 5724 1284
rect 5776 1272 5782 1284
rect 7834 1272 7840 1284
rect 5776 1244 7840 1272
rect 5776 1232 5782 1244
rect 7834 1232 7840 1244
rect 7892 1232 7898 1284
rect 6914 552 6920 604
rect 6972 592 6978 604
rect 7098 592 7104 604
rect 6972 564 7104 592
rect 6972 552 6978 564
rect 7098 552 7104 564
rect 7156 552 7162 604
rect 9950 552 9956 604
rect 10008 592 10014 604
rect 10134 592 10140 604
rect 10008 564 10140 592
rect 10008 552 10014 564
rect 10134 552 10140 564
rect 10192 552 10198 604
rect 10594 552 10600 604
rect 10652 592 10658 604
rect 10870 592 10876 604
rect 10652 564 10876 592
rect 10652 552 10658 564
rect 10870 552 10876 564
rect 10928 552 10934 604
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 4528 36320 4580 36372
rect 5540 36363 5592 36372
rect 5540 36329 5549 36363
rect 5549 36329 5583 36363
rect 5583 36329 5592 36363
rect 5540 36320 5592 36329
rect 4252 36227 4304 36236
rect 4252 36193 4261 36227
rect 4261 36193 4295 36227
rect 4295 36193 4304 36227
rect 4252 36184 4304 36193
rect 5448 36184 5500 36236
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 572 35776 624 35828
rect 2596 35776 2648 35828
rect 3976 35776 4028 35828
rect 6184 35776 6236 35828
rect 6920 35776 6972 35828
rect 8024 35708 8076 35760
rect 3240 35572 3292 35624
rect 5540 35504 5592 35556
rect 10324 35572 10376 35624
rect 2228 35436 2280 35488
rect 4252 35436 4304 35488
rect 5448 35479 5500 35488
rect 5448 35445 5457 35479
rect 5457 35445 5491 35479
rect 5491 35445 5500 35479
rect 5448 35436 5500 35445
rect 6000 35436 6052 35488
rect 7472 35479 7524 35488
rect 7472 35445 7481 35479
rect 7481 35445 7515 35479
rect 7515 35445 7524 35479
rect 7472 35436 7524 35445
rect 8300 35436 8352 35488
rect 9220 35479 9272 35488
rect 9220 35445 9229 35479
rect 9229 35445 9263 35479
rect 9263 35445 9272 35479
rect 9220 35436 9272 35445
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 204 35232 256 35284
rect 2136 35232 2188 35284
rect 4160 35232 4212 35284
rect 6644 35232 6696 35284
rect 7748 35232 7800 35284
rect 10140 35232 10192 35284
rect 15384 35232 15436 35284
rect 1860 35096 1912 35148
rect 2504 35139 2556 35148
rect 2504 35105 2513 35139
rect 2513 35105 2547 35139
rect 2547 35105 2556 35139
rect 2504 35096 2556 35105
rect 4068 35139 4120 35148
rect 4068 35105 4077 35139
rect 4077 35105 4111 35139
rect 4111 35105 4120 35139
rect 4068 35096 4120 35105
rect 6184 35096 6236 35148
rect 6920 35139 6972 35148
rect 6920 35105 6929 35139
rect 6929 35105 6963 35139
rect 6963 35105 6972 35139
rect 6920 35096 6972 35105
rect 8392 35139 8444 35148
rect 8392 35105 8401 35139
rect 8401 35105 8435 35139
rect 8435 35105 8444 35139
rect 8392 35096 8444 35105
rect 10968 35096 11020 35148
rect 8668 35071 8720 35080
rect 7932 35003 7984 35012
rect 7932 34969 7941 35003
rect 7941 34969 7975 35003
rect 7975 34969 7984 35003
rect 8668 35037 8677 35071
rect 8677 35037 8711 35071
rect 8711 35037 8720 35071
rect 8668 35028 8720 35037
rect 10784 35071 10836 35080
rect 10784 35037 10793 35071
rect 10793 35037 10827 35071
rect 10827 35037 10836 35071
rect 10784 35028 10836 35037
rect 7932 34960 7984 34969
rect 2044 34935 2096 34944
rect 2044 34901 2053 34935
rect 2053 34901 2087 34935
rect 2087 34901 2096 34935
rect 2044 34892 2096 34901
rect 3516 34935 3568 34944
rect 3516 34901 3525 34935
rect 3525 34901 3559 34935
rect 3559 34901 3568 34935
rect 3516 34892 3568 34901
rect 8024 34935 8076 34944
rect 8024 34901 8033 34935
rect 8033 34901 8067 34935
rect 8067 34901 8076 34935
rect 8024 34892 8076 34901
rect 8852 34892 8904 34944
rect 10416 34892 10468 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 4068 34688 4120 34740
rect 7380 34688 7432 34740
rect 10968 34688 11020 34740
rect 1860 34620 1912 34672
rect 2596 34620 2648 34672
rect 8484 34663 8536 34672
rect 8484 34629 8493 34663
rect 8493 34629 8527 34663
rect 8527 34629 8536 34663
rect 8484 34620 8536 34629
rect 8852 34620 8904 34672
rect 10784 34620 10836 34672
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 8024 34552 8076 34604
rect 8944 34595 8996 34604
rect 8944 34561 8953 34595
rect 8953 34561 8987 34595
rect 8987 34561 8996 34595
rect 8944 34552 8996 34561
rect 2044 34484 2096 34536
rect 2504 34527 2556 34536
rect 2504 34493 2513 34527
rect 2513 34493 2547 34527
rect 2547 34493 2556 34527
rect 2504 34484 2556 34493
rect 3516 34484 3568 34536
rect 4068 34484 4120 34536
rect 6184 34484 6236 34536
rect 8208 34484 8260 34536
rect 8852 34527 8904 34536
rect 3700 34459 3752 34468
rect 3700 34425 3734 34459
rect 3734 34425 3752 34459
rect 3700 34416 3752 34425
rect 8852 34493 8861 34527
rect 8861 34493 8895 34527
rect 8895 34493 8904 34527
rect 8852 34484 8904 34493
rect 9128 34552 9180 34604
rect 11428 34552 11480 34604
rect 10140 34484 10192 34536
rect 10416 34527 10468 34536
rect 10416 34493 10425 34527
rect 10425 34493 10459 34527
rect 10459 34493 10468 34527
rect 10416 34484 10468 34493
rect 10508 34527 10560 34536
rect 10508 34493 10517 34527
rect 10517 34493 10551 34527
rect 10551 34493 10560 34527
rect 10508 34484 10560 34493
rect 9956 34416 10008 34468
rect 4620 34348 4672 34400
rect 6920 34348 6972 34400
rect 7656 34348 7708 34400
rect 11428 34391 11480 34400
rect 11428 34357 11437 34391
rect 11437 34357 11471 34391
rect 11471 34357 11480 34391
rect 11428 34348 11480 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 1768 34144 1820 34196
rect 8944 34187 8996 34196
rect 1676 34119 1728 34128
rect 1676 34085 1685 34119
rect 1685 34085 1719 34119
rect 1719 34085 1728 34119
rect 1676 34076 1728 34085
rect 4620 34076 4672 34128
rect 8944 34153 8953 34187
rect 8953 34153 8987 34187
rect 8987 34153 8996 34187
rect 8944 34144 8996 34153
rect 11428 34144 11480 34196
rect 6736 34076 6788 34128
rect 8668 34119 8720 34128
rect 8668 34085 8677 34119
rect 8677 34085 8711 34119
rect 8711 34085 8720 34119
rect 8668 34076 8720 34085
rect 9128 34076 9180 34128
rect 10140 34119 10192 34128
rect 10140 34085 10174 34119
rect 10174 34085 10192 34119
rect 10140 34076 10192 34085
rect 10784 34076 10836 34128
rect 1492 34008 1544 34060
rect 2964 34008 3016 34060
rect 4068 34008 4120 34060
rect 5816 34008 5868 34060
rect 3700 33872 3752 33924
rect 4344 33804 4396 33856
rect 5816 33804 5868 33856
rect 9312 33940 9364 33992
rect 8024 33847 8076 33856
rect 8024 33813 8033 33847
rect 8033 33813 8067 33847
rect 8067 33813 8076 33847
rect 8024 33804 8076 33813
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 1400 33600 1452 33652
rect 5724 33600 5776 33652
rect 8668 33643 8720 33652
rect 8668 33609 8677 33643
rect 8677 33609 8711 33643
rect 8711 33609 8720 33643
rect 8668 33600 8720 33609
rect 9772 33600 9824 33652
rect 9956 33600 10008 33652
rect 1492 33532 1544 33584
rect 8576 33532 8628 33584
rect 2412 33507 2464 33516
rect 2412 33473 2421 33507
rect 2421 33473 2455 33507
rect 2455 33473 2464 33507
rect 2412 33464 2464 33473
rect 6736 33464 6788 33516
rect 4068 33396 4120 33448
rect 4804 33396 4856 33448
rect 11060 33464 11112 33516
rect 3056 33328 3108 33380
rect 2964 33260 3016 33312
rect 4344 33303 4396 33312
rect 4344 33269 4353 33303
rect 4353 33269 4387 33303
rect 4387 33269 4396 33303
rect 4344 33260 4396 33269
rect 4620 33260 4672 33312
rect 5816 33260 5868 33312
rect 6092 33260 6144 33312
rect 8208 33328 8260 33380
rect 9312 33328 9364 33380
rect 6644 33260 6696 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 4068 33056 4120 33108
rect 4988 33056 5040 33108
rect 6736 33099 6788 33108
rect 6736 33065 6745 33099
rect 6745 33065 6779 33099
rect 6779 33065 6788 33099
rect 6736 33056 6788 33065
rect 7288 33099 7340 33108
rect 7288 33065 7297 33099
rect 7297 33065 7331 33099
rect 7331 33065 7340 33099
rect 7288 33056 7340 33065
rect 10508 33056 10560 33108
rect 10784 32988 10836 33040
rect 4436 32920 4488 32972
rect 9496 32920 9548 32972
rect 10140 32920 10192 32972
rect 10232 32920 10284 32972
rect 6644 32852 6696 32904
rect 6276 32784 6328 32836
rect 8024 32852 8076 32904
rect 10876 32852 10928 32904
rect 3056 32759 3108 32768
rect 3056 32725 3065 32759
rect 3065 32725 3099 32759
rect 3099 32725 3108 32759
rect 3056 32716 3108 32725
rect 3424 32759 3476 32768
rect 3424 32725 3433 32759
rect 3433 32725 3467 32759
rect 3467 32725 3476 32759
rect 3424 32716 3476 32725
rect 4528 32759 4580 32768
rect 4528 32725 4537 32759
rect 4537 32725 4571 32759
rect 4571 32725 4580 32759
rect 4528 32716 4580 32725
rect 5264 32759 5316 32768
rect 5264 32725 5273 32759
rect 5273 32725 5307 32759
rect 5307 32725 5316 32759
rect 5264 32716 5316 32725
rect 5356 32716 5408 32768
rect 6920 32759 6972 32768
rect 6920 32725 6929 32759
rect 6929 32725 6963 32759
rect 6963 32725 6972 32759
rect 6920 32716 6972 32725
rect 9312 32759 9364 32768
rect 9312 32725 9321 32759
rect 9321 32725 9355 32759
rect 9355 32725 9364 32759
rect 9312 32716 9364 32725
rect 12532 32759 12584 32768
rect 12532 32725 12541 32759
rect 12541 32725 12575 32759
rect 12575 32725 12584 32759
rect 12532 32716 12584 32725
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 6276 32555 6328 32564
rect 6276 32521 6285 32555
rect 6285 32521 6319 32555
rect 6319 32521 6328 32555
rect 6276 32512 6328 32521
rect 7288 32512 7340 32564
rect 7472 32512 7524 32564
rect 8392 32512 8444 32564
rect 10876 32555 10928 32564
rect 10876 32521 10885 32555
rect 10885 32521 10919 32555
rect 10919 32521 10928 32555
rect 10876 32512 10928 32521
rect 1584 32419 1636 32428
rect 1584 32385 1593 32419
rect 1593 32385 1627 32419
rect 1627 32385 1636 32419
rect 1584 32376 1636 32385
rect 3424 32376 3476 32428
rect 4344 32444 4396 32496
rect 5264 32444 5316 32496
rect 5356 32419 5408 32428
rect 5356 32385 5365 32419
rect 5365 32385 5399 32419
rect 5399 32385 5408 32419
rect 5356 32376 5408 32385
rect 7564 32444 7616 32496
rect 10232 32487 10284 32496
rect 5540 32376 5592 32428
rect 4528 32308 4580 32360
rect 6828 32308 6880 32360
rect 4160 32240 4212 32292
rect 2228 32215 2280 32224
rect 2228 32181 2237 32215
rect 2237 32181 2271 32215
rect 2271 32181 2280 32215
rect 2228 32172 2280 32181
rect 3332 32215 3384 32224
rect 3332 32181 3341 32215
rect 3341 32181 3375 32215
rect 3375 32181 3384 32215
rect 3332 32172 3384 32181
rect 4436 32172 4488 32224
rect 4896 32215 4948 32224
rect 4896 32181 4905 32215
rect 4905 32181 4939 32215
rect 4939 32181 4948 32215
rect 4896 32172 4948 32181
rect 7288 32215 7340 32224
rect 7288 32181 7297 32215
rect 7297 32181 7331 32215
rect 7331 32181 7340 32215
rect 7288 32172 7340 32181
rect 8024 32376 8076 32428
rect 10232 32453 10241 32487
rect 10241 32453 10275 32487
rect 10275 32453 10284 32487
rect 10232 32444 10284 32453
rect 9496 32419 9548 32428
rect 9496 32385 9505 32419
rect 9505 32385 9539 32419
rect 9539 32385 9548 32419
rect 9496 32376 9548 32385
rect 10140 32376 10192 32428
rect 10784 32444 10836 32496
rect 12532 32376 12584 32428
rect 12900 32419 12952 32428
rect 12900 32385 12909 32419
rect 12909 32385 12943 32419
rect 12943 32385 12952 32419
rect 12900 32376 12952 32385
rect 13084 32419 13136 32428
rect 13084 32385 13093 32419
rect 13093 32385 13127 32419
rect 13127 32385 13136 32419
rect 13084 32376 13136 32385
rect 12164 32308 12216 32360
rect 7840 32240 7892 32292
rect 9404 32240 9456 32292
rect 12532 32240 12584 32292
rect 8668 32172 8720 32224
rect 8852 32172 8904 32224
rect 12440 32215 12492 32224
rect 12440 32181 12449 32215
rect 12449 32181 12483 32215
rect 12483 32181 12492 32215
rect 12440 32172 12492 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 2780 31968 2832 32020
rect 3332 31968 3384 32020
rect 5356 31968 5408 32020
rect 6644 31968 6696 32020
rect 6828 32011 6880 32020
rect 6828 31977 6837 32011
rect 6837 31977 6871 32011
rect 6871 31977 6880 32011
rect 6828 31968 6880 31977
rect 8576 31968 8628 32020
rect 9404 31968 9456 32020
rect 10508 32011 10560 32020
rect 10508 31977 10517 32011
rect 10517 31977 10551 32011
rect 10551 31977 10560 32011
rect 10508 31968 10560 31977
rect 13084 31968 13136 32020
rect 13820 31968 13872 32020
rect 6736 31900 6788 31952
rect 8484 31900 8536 31952
rect 8852 31943 8904 31952
rect 8852 31909 8861 31943
rect 8861 31909 8895 31943
rect 8895 31909 8904 31943
rect 8852 31900 8904 31909
rect 2872 31832 2924 31884
rect 4896 31832 4948 31884
rect 6184 31832 6236 31884
rect 6552 31832 6604 31884
rect 8208 31832 8260 31884
rect 9496 31832 9548 31884
rect 10876 31875 10928 31884
rect 10876 31841 10885 31875
rect 10885 31841 10919 31875
rect 10919 31841 10928 31875
rect 10876 31832 10928 31841
rect 12348 31875 12400 31884
rect 12348 31841 12382 31875
rect 12382 31841 12400 31875
rect 12348 31832 12400 31841
rect 5724 31807 5776 31816
rect 2688 31696 2740 31748
rect 5724 31773 5733 31807
rect 5733 31773 5767 31807
rect 5767 31773 5776 31807
rect 5724 31764 5776 31773
rect 4620 31696 4672 31748
rect 5540 31696 5592 31748
rect 6828 31764 6880 31816
rect 7288 31764 7340 31816
rect 10324 31764 10376 31816
rect 8208 31696 8260 31748
rect 10600 31764 10652 31816
rect 10784 31764 10836 31816
rect 12072 31807 12124 31816
rect 10508 31696 10560 31748
rect 12072 31773 12081 31807
rect 12081 31773 12115 31807
rect 12115 31773 12124 31807
rect 12072 31764 12124 31773
rect 11152 31696 11204 31748
rect 2412 31671 2464 31680
rect 2412 31637 2421 31671
rect 2421 31637 2455 31671
rect 2455 31637 2464 31671
rect 2412 31628 2464 31637
rect 4528 31671 4580 31680
rect 4528 31637 4537 31671
rect 4537 31637 4571 31671
rect 4571 31637 4580 31671
rect 4528 31628 4580 31637
rect 7380 31628 7432 31680
rect 7748 31628 7800 31680
rect 8024 31628 8076 31680
rect 8484 31671 8536 31680
rect 8484 31637 8493 31671
rect 8493 31637 8527 31671
rect 8527 31637 8536 31671
rect 8484 31628 8536 31637
rect 9864 31628 9916 31680
rect 10048 31628 10100 31680
rect 10416 31628 10468 31680
rect 11520 31671 11572 31680
rect 11520 31637 11529 31671
rect 11529 31637 11563 31671
rect 11563 31637 11572 31671
rect 11520 31628 11572 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 2688 31424 2740 31476
rect 3424 31424 3476 31476
rect 4160 31424 4212 31476
rect 6092 31424 6144 31476
rect 6736 31424 6788 31476
rect 7104 31424 7156 31476
rect 7748 31424 7800 31476
rect 8208 31467 8260 31476
rect 8208 31433 8217 31467
rect 8217 31433 8251 31467
rect 8251 31433 8260 31467
rect 8208 31424 8260 31433
rect 8392 31467 8444 31476
rect 8392 31433 8401 31467
rect 8401 31433 8435 31467
rect 8435 31433 8444 31467
rect 8392 31424 8444 31433
rect 9496 31424 9548 31476
rect 9864 31424 9916 31476
rect 12532 31467 12584 31476
rect 12532 31433 12541 31467
rect 12541 31433 12575 31467
rect 12575 31433 12584 31467
rect 12532 31424 12584 31433
rect 5632 31356 5684 31408
rect 6552 31356 6604 31408
rect 1584 31331 1636 31340
rect 1584 31297 1593 31331
rect 1593 31297 1627 31331
rect 1627 31297 1636 31331
rect 1584 31288 1636 31297
rect 3056 31288 3108 31340
rect 5540 31331 5592 31340
rect 5540 31297 5549 31331
rect 5549 31297 5583 31331
rect 5583 31297 5592 31331
rect 5540 31288 5592 31297
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 8484 31288 8536 31340
rect 10784 31288 10836 31340
rect 1676 31220 1728 31272
rect 2412 31220 2464 31272
rect 6828 31220 6880 31272
rect 3976 31152 4028 31204
rect 4528 31152 4580 31204
rect 3792 31127 3844 31136
rect 3792 31093 3801 31127
rect 3801 31093 3835 31127
rect 3835 31093 3844 31127
rect 3792 31084 3844 31093
rect 4436 31084 4488 31136
rect 5080 31084 5132 31136
rect 6184 31084 6236 31136
rect 6828 31127 6880 31136
rect 6828 31093 6837 31127
rect 6837 31093 6871 31127
rect 6871 31093 6880 31127
rect 6828 31084 6880 31093
rect 10968 31220 11020 31272
rect 12348 31220 12400 31272
rect 12808 31220 12860 31272
rect 8576 31152 8628 31204
rect 10324 31152 10376 31204
rect 11428 31152 11480 31204
rect 13084 31152 13136 31204
rect 7288 31127 7340 31136
rect 7288 31093 7297 31127
rect 7297 31093 7331 31127
rect 7331 31093 7340 31127
rect 8760 31127 8812 31136
rect 7288 31084 7340 31093
rect 8760 31093 8769 31127
rect 8769 31093 8803 31127
rect 8803 31093 8812 31127
rect 8760 31084 8812 31093
rect 11060 31084 11112 31136
rect 11520 31084 11572 31136
rect 12348 31084 12400 31136
rect 13268 31084 13320 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 1676 30923 1728 30932
rect 1676 30889 1685 30923
rect 1685 30889 1719 30923
rect 1719 30889 1728 30923
rect 1676 30880 1728 30889
rect 2688 30880 2740 30932
rect 2872 30923 2924 30932
rect 2872 30889 2881 30923
rect 2881 30889 2915 30923
rect 2915 30889 2924 30923
rect 2872 30880 2924 30889
rect 3516 30880 3568 30932
rect 3792 30880 3844 30932
rect 3976 30880 4028 30932
rect 5356 30923 5408 30932
rect 5356 30889 5365 30923
rect 5365 30889 5399 30923
rect 5399 30889 5408 30923
rect 5356 30880 5408 30889
rect 5632 30923 5684 30932
rect 5632 30889 5641 30923
rect 5641 30889 5675 30923
rect 5675 30889 5684 30923
rect 5632 30880 5684 30889
rect 6920 30880 6972 30932
rect 7288 30880 7340 30932
rect 8024 30923 8076 30932
rect 8024 30889 8033 30923
rect 8033 30889 8067 30923
rect 8067 30889 8076 30923
rect 8024 30880 8076 30889
rect 8392 30880 8444 30932
rect 8576 30923 8628 30932
rect 8576 30889 8585 30923
rect 8585 30889 8619 30923
rect 8619 30889 8628 30923
rect 8576 30880 8628 30889
rect 6736 30812 6788 30864
rect 12164 30812 12216 30864
rect 2044 30744 2096 30796
rect 4436 30787 4488 30796
rect 4436 30753 4445 30787
rect 4445 30753 4479 30787
rect 4479 30753 4488 30787
rect 4436 30744 4488 30753
rect 4988 30744 5040 30796
rect 6920 30787 6972 30796
rect 6920 30753 6954 30787
rect 6954 30753 6972 30787
rect 6920 30744 6972 30753
rect 7380 30744 7432 30796
rect 10876 30787 10928 30796
rect 10876 30753 10885 30787
rect 10885 30753 10919 30787
rect 10919 30753 10928 30787
rect 10876 30744 10928 30753
rect 12072 30787 12124 30796
rect 12072 30753 12081 30787
rect 12081 30753 12115 30787
rect 12115 30753 12124 30787
rect 12072 30744 12124 30753
rect 940 30608 992 30660
rect 4804 30676 4856 30728
rect 6552 30676 6604 30728
rect 10600 30676 10652 30728
rect 10968 30540 11020 30592
rect 12808 30540 12860 30592
rect 13452 30583 13504 30592
rect 13452 30549 13461 30583
rect 13461 30549 13495 30583
rect 13495 30549 13504 30583
rect 13452 30540 13504 30549
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 3516 30336 3568 30388
rect 6184 30336 6236 30388
rect 6736 30336 6788 30388
rect 10876 30336 10928 30388
rect 12440 30379 12492 30388
rect 12440 30345 12449 30379
rect 12449 30345 12483 30379
rect 12483 30345 12492 30379
rect 12440 30336 12492 30345
rect 9680 30311 9732 30320
rect 9680 30277 9689 30311
rect 9689 30277 9723 30311
rect 9723 30277 9732 30311
rect 9680 30268 9732 30277
rect 11520 30268 11572 30320
rect 11980 30268 12032 30320
rect 13820 30311 13872 30320
rect 4804 30200 4856 30252
rect 2044 30175 2096 30184
rect 2044 30141 2053 30175
rect 2053 30141 2087 30175
rect 2087 30141 2096 30175
rect 2044 30132 2096 30141
rect 4988 30132 5040 30184
rect 2596 29996 2648 30048
rect 5264 30064 5316 30116
rect 4160 30039 4212 30048
rect 4160 30005 4169 30039
rect 4169 30005 4203 30039
rect 4203 30005 4212 30039
rect 4160 29996 4212 30005
rect 4988 29996 5040 30048
rect 5816 30200 5868 30252
rect 6552 30200 6604 30252
rect 13820 30277 13829 30311
rect 13829 30277 13863 30311
rect 13863 30277 13872 30311
rect 13820 30268 13872 30277
rect 7288 30175 7340 30184
rect 7288 30141 7297 30175
rect 7297 30141 7331 30175
rect 7331 30141 7340 30175
rect 7288 30132 7340 30141
rect 13452 30200 13504 30252
rect 8024 30132 8076 30184
rect 9312 30132 9364 30184
rect 9680 30132 9732 30184
rect 10324 30132 10376 30184
rect 12348 30132 12400 30184
rect 5724 29996 5776 30048
rect 6644 30039 6696 30048
rect 6644 30005 6653 30039
rect 6653 30005 6687 30039
rect 6687 30005 6696 30039
rect 6644 29996 6696 30005
rect 6920 29996 6972 30048
rect 8668 30039 8720 30048
rect 8668 30005 8677 30039
rect 8677 30005 8711 30039
rect 8711 30005 8720 30039
rect 8668 29996 8720 30005
rect 11244 29996 11296 30048
rect 12256 29996 12308 30048
rect 13452 30039 13504 30048
rect 13452 30005 13461 30039
rect 13461 30005 13495 30039
rect 13495 30005 13504 30039
rect 13452 29996 13504 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 4436 29792 4488 29844
rect 5540 29792 5592 29844
rect 7932 29792 7984 29844
rect 4160 29724 4212 29776
rect 4804 29656 4856 29708
rect 7288 29724 7340 29776
rect 10876 29792 10928 29844
rect 8116 29656 8168 29708
rect 8392 29699 8444 29708
rect 8392 29665 8401 29699
rect 8401 29665 8435 29699
rect 8435 29665 8444 29699
rect 8392 29656 8444 29665
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 8576 29631 8628 29640
rect 8576 29597 8585 29631
rect 8585 29597 8619 29631
rect 8619 29597 8628 29631
rect 9772 29724 9824 29776
rect 11152 29724 11204 29776
rect 12072 29767 12124 29776
rect 12072 29733 12081 29767
rect 12081 29733 12115 29767
rect 12115 29733 12124 29767
rect 12072 29724 12124 29733
rect 12256 29724 12308 29776
rect 10324 29656 10376 29708
rect 12532 29699 12584 29708
rect 12532 29665 12541 29699
rect 12541 29665 12575 29699
rect 12575 29665 12584 29699
rect 12532 29656 12584 29665
rect 8576 29588 8628 29597
rect 11152 29520 11204 29572
rect 11244 29520 11296 29572
rect 13452 29588 13504 29640
rect 4988 29452 5040 29504
rect 6920 29495 6972 29504
rect 6920 29461 6929 29495
rect 6929 29461 6963 29495
rect 6963 29461 6972 29495
rect 6920 29452 6972 29461
rect 12808 29452 12860 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 3240 29248 3292 29300
rect 4528 29291 4580 29300
rect 4528 29257 4537 29291
rect 4537 29257 4571 29291
rect 4571 29257 4580 29291
rect 4528 29248 4580 29257
rect 6828 29291 6880 29300
rect 6828 29257 6837 29291
rect 6837 29257 6871 29291
rect 6871 29257 6880 29291
rect 6828 29248 6880 29257
rect 8484 29248 8536 29300
rect 9772 29248 9824 29300
rect 10048 29248 10100 29300
rect 10600 29291 10652 29300
rect 10600 29257 10609 29291
rect 10609 29257 10643 29291
rect 10643 29257 10652 29291
rect 10600 29248 10652 29257
rect 12900 29248 12952 29300
rect 13452 29248 13504 29300
rect 6644 29223 6696 29232
rect 6644 29189 6653 29223
rect 6653 29189 6687 29223
rect 6687 29189 6696 29223
rect 6644 29180 6696 29189
rect 4804 29112 4856 29164
rect 6920 29112 6972 29164
rect 7288 29155 7340 29164
rect 7288 29121 7297 29155
rect 7297 29121 7331 29155
rect 7331 29121 7340 29155
rect 7288 29112 7340 29121
rect 8208 29112 8260 29164
rect 8484 29155 8536 29164
rect 8484 29121 8493 29155
rect 8493 29121 8527 29155
rect 8527 29121 8536 29155
rect 8484 29112 8536 29121
rect 8668 29112 8720 29164
rect 9128 29112 9180 29164
rect 10324 29180 10376 29232
rect 10508 29180 10560 29232
rect 9864 29112 9916 29164
rect 10600 29112 10652 29164
rect 11244 29155 11296 29164
rect 11244 29121 11253 29155
rect 11253 29121 11287 29155
rect 11287 29121 11296 29155
rect 11244 29112 11296 29121
rect 11980 29180 12032 29232
rect 12256 29112 12308 29164
rect 12808 29112 12860 29164
rect 5172 29044 5224 29096
rect 6092 29044 6144 29096
rect 6644 29044 6696 29096
rect 7196 29019 7248 29028
rect 7196 28985 7205 29019
rect 7205 28985 7239 29019
rect 7239 28985 7248 29019
rect 7196 28976 7248 28985
rect 8392 28976 8444 29028
rect 10324 29044 10376 29096
rect 12900 29087 12952 29096
rect 12900 29053 12909 29087
rect 12909 29053 12943 29087
rect 12943 29053 12952 29087
rect 12900 29044 12952 29053
rect 9404 28976 9456 29028
rect 10876 28976 10928 29028
rect 13452 28976 13504 29028
rect 3332 28908 3384 28960
rect 8668 28908 8720 28960
rect 10416 28908 10468 28960
rect 10508 28908 10560 28960
rect 10600 28908 10652 28960
rect 12900 28908 12952 28960
rect 14188 28976 14240 29028
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 2964 28704 3016 28756
rect 4068 28704 4120 28756
rect 7196 28704 7248 28756
rect 8576 28704 8628 28756
rect 9128 28747 9180 28756
rect 9128 28713 9137 28747
rect 9137 28713 9171 28747
rect 9171 28713 9180 28747
rect 9128 28704 9180 28713
rect 10048 28704 10100 28756
rect 10324 28747 10376 28756
rect 10324 28713 10333 28747
rect 10333 28713 10367 28747
rect 10367 28713 10376 28747
rect 10324 28704 10376 28713
rect 10968 28704 11020 28756
rect 11980 28747 12032 28756
rect 11980 28713 11989 28747
rect 11989 28713 12023 28747
rect 12023 28713 12032 28747
rect 11980 28704 12032 28713
rect 12532 28704 12584 28756
rect 13084 28747 13136 28756
rect 13084 28713 13093 28747
rect 13093 28713 13127 28747
rect 13127 28713 13136 28747
rect 13084 28704 13136 28713
rect 7932 28636 7984 28688
rect 11152 28636 11204 28688
rect 8760 28568 8812 28620
rect 11244 28568 11296 28620
rect 7748 28543 7800 28552
rect 7748 28509 7757 28543
rect 7757 28509 7791 28543
rect 7791 28509 7800 28543
rect 7748 28500 7800 28509
rect 7840 28543 7892 28552
rect 7840 28509 7849 28543
rect 7849 28509 7883 28543
rect 7883 28509 7892 28543
rect 12164 28543 12216 28552
rect 7840 28500 7892 28509
rect 12164 28509 12173 28543
rect 12173 28509 12207 28543
rect 12207 28509 12216 28543
rect 12164 28500 12216 28509
rect 4344 28364 4396 28416
rect 5172 28432 5224 28484
rect 7104 28432 7156 28484
rect 10784 28432 10836 28484
rect 4988 28407 5040 28416
rect 4988 28373 4997 28407
rect 4997 28373 5031 28407
rect 5031 28373 5040 28407
rect 4988 28364 5040 28373
rect 6828 28364 6880 28416
rect 8116 28364 8168 28416
rect 8576 28364 8628 28416
rect 10600 28364 10652 28416
rect 10968 28364 11020 28416
rect 12532 28407 12584 28416
rect 12532 28373 12541 28407
rect 12541 28373 12575 28407
rect 12575 28373 12584 28407
rect 12532 28364 12584 28373
rect 12900 28364 12952 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 7748 28160 7800 28212
rect 8208 28203 8260 28212
rect 8208 28169 8217 28203
rect 8217 28169 8251 28203
rect 8251 28169 8260 28203
rect 8208 28160 8260 28169
rect 8760 28203 8812 28212
rect 8760 28169 8769 28203
rect 8769 28169 8803 28203
rect 8803 28169 8812 28203
rect 8760 28160 8812 28169
rect 11152 28203 11204 28212
rect 11152 28169 11161 28203
rect 11161 28169 11195 28203
rect 11195 28169 11204 28203
rect 11152 28160 11204 28169
rect 11980 28203 12032 28212
rect 11980 28169 11989 28203
rect 11989 28169 12023 28203
rect 12023 28169 12032 28203
rect 11980 28160 12032 28169
rect 12164 28092 12216 28144
rect 11152 28024 11204 28076
rect 11428 28024 11480 28076
rect 6828 27999 6880 28008
rect 6828 27965 6837 27999
rect 6837 27965 6871 27999
rect 6871 27965 6880 27999
rect 6828 27956 6880 27965
rect 6920 27888 6972 27940
rect 5356 27863 5408 27872
rect 5356 27829 5365 27863
rect 5365 27829 5399 27863
rect 5399 27829 5408 27863
rect 5356 27820 5408 27829
rect 7840 27888 7892 27940
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 5356 27616 5408 27668
rect 1676 27591 1728 27600
rect 1676 27557 1685 27591
rect 1685 27557 1719 27591
rect 1719 27557 1728 27591
rect 1676 27548 1728 27557
rect 8116 27616 8168 27668
rect 7748 27548 7800 27600
rect 8852 27548 8904 27600
rect 10324 27616 10376 27668
rect 12808 27659 12860 27668
rect 12808 27625 12817 27659
rect 12817 27625 12851 27659
rect 12851 27625 12860 27659
rect 12808 27616 12860 27625
rect 11244 27548 11296 27600
rect 6000 27523 6052 27532
rect 6000 27489 6009 27523
rect 6009 27489 6043 27523
rect 6043 27489 6052 27523
rect 6000 27480 6052 27489
rect 8116 27480 8168 27532
rect 9680 27480 9732 27532
rect 1676 27412 1728 27464
rect 6092 27455 6144 27464
rect 5724 27344 5776 27396
rect 6092 27421 6101 27455
rect 6101 27421 6135 27455
rect 6135 27421 6144 27455
rect 6092 27412 6144 27421
rect 7380 27412 7432 27464
rect 7840 27455 7892 27464
rect 7840 27421 7849 27455
rect 7849 27421 7883 27455
rect 7883 27421 7892 27455
rect 11428 27455 11480 27464
rect 7840 27412 7892 27421
rect 11428 27421 11437 27455
rect 11437 27421 11471 27455
rect 11471 27421 11480 27455
rect 11428 27412 11480 27421
rect 6828 27387 6880 27396
rect 6828 27353 6837 27387
rect 6837 27353 6871 27387
rect 6871 27353 6880 27387
rect 6828 27344 6880 27353
rect 7288 27387 7340 27396
rect 7288 27353 7297 27387
rect 7297 27353 7331 27387
rect 7331 27353 7340 27387
rect 7288 27344 7340 27353
rect 5172 27319 5224 27328
rect 5172 27285 5181 27319
rect 5181 27285 5215 27319
rect 5215 27285 5224 27319
rect 5172 27276 5224 27285
rect 5540 27276 5592 27328
rect 8760 27319 8812 27328
rect 8760 27285 8769 27319
rect 8769 27285 8803 27319
rect 8803 27285 8812 27319
rect 8760 27276 8812 27285
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 4804 27115 4856 27124
rect 4804 27081 4813 27115
rect 4813 27081 4847 27115
rect 4847 27081 4856 27115
rect 4804 27072 4856 27081
rect 6092 27115 6144 27124
rect 6092 27081 6101 27115
rect 6101 27081 6135 27115
rect 6135 27081 6144 27115
rect 6092 27072 6144 27081
rect 9680 27115 9732 27124
rect 9680 27081 9689 27115
rect 9689 27081 9723 27115
rect 9723 27081 9732 27115
rect 9680 27072 9732 27081
rect 11244 27072 11296 27124
rect 6000 27004 6052 27056
rect 10508 27004 10560 27056
rect 12072 27004 12124 27056
rect 6828 26936 6880 26988
rect 8760 26936 8812 26988
rect 3424 26911 3476 26920
rect 3424 26877 3433 26911
rect 3433 26877 3467 26911
rect 3467 26877 3476 26911
rect 3424 26868 3476 26877
rect 6920 26868 6972 26920
rect 8668 26868 8720 26920
rect 9036 26868 9088 26920
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 2964 26732 3016 26784
rect 7288 26843 7340 26852
rect 7288 26809 7297 26843
rect 7297 26809 7331 26843
rect 7331 26809 7340 26843
rect 7288 26800 7340 26809
rect 6828 26775 6880 26784
rect 6828 26741 6837 26775
rect 6837 26741 6871 26775
rect 6871 26741 6880 26775
rect 6828 26732 6880 26741
rect 7748 26732 7800 26784
rect 8208 26732 8260 26784
rect 8392 26732 8444 26784
rect 8668 26775 8720 26784
rect 8668 26741 8677 26775
rect 8677 26741 8711 26775
rect 8711 26741 8720 26775
rect 8668 26732 8720 26741
rect 9036 26775 9088 26784
rect 9036 26741 9045 26775
rect 9045 26741 9079 26775
rect 9079 26741 9088 26775
rect 9036 26732 9088 26741
rect 9772 26732 9824 26784
rect 10692 26732 10744 26784
rect 11244 26732 11296 26784
rect 11428 26732 11480 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 1676 26528 1728 26580
rect 3424 26571 3476 26580
rect 3424 26537 3433 26571
rect 3433 26537 3467 26571
rect 3467 26537 3476 26571
rect 3424 26528 3476 26537
rect 6920 26571 6972 26580
rect 6920 26537 6929 26571
rect 6929 26537 6963 26571
rect 6963 26537 6972 26571
rect 6920 26528 6972 26537
rect 7380 26571 7432 26580
rect 7380 26537 7389 26571
rect 7389 26537 7423 26571
rect 7423 26537 7432 26571
rect 7380 26528 7432 26537
rect 7840 26528 7892 26580
rect 2780 26503 2832 26512
rect 2780 26469 2789 26503
rect 2789 26469 2823 26503
rect 2823 26469 2832 26503
rect 2780 26460 2832 26469
rect 3976 26460 4028 26512
rect 2872 26435 2924 26444
rect 2872 26401 2881 26435
rect 2881 26401 2915 26435
rect 2915 26401 2924 26435
rect 4988 26460 5040 26512
rect 5632 26460 5684 26512
rect 10048 26460 10100 26512
rect 2872 26392 2924 26401
rect 5172 26435 5224 26444
rect 5172 26401 5206 26435
rect 5206 26401 5224 26435
rect 5172 26392 5224 26401
rect 2964 26367 3016 26376
rect 2964 26333 2973 26367
rect 2973 26333 3007 26367
rect 3007 26333 3016 26367
rect 2964 26324 3016 26333
rect 5908 26256 5960 26308
rect 8392 26188 8444 26240
rect 9036 26256 9088 26308
rect 9312 26188 9364 26240
rect 11428 26299 11480 26308
rect 11428 26265 11437 26299
rect 11437 26265 11471 26299
rect 11471 26265 11480 26299
rect 11428 26256 11480 26265
rect 10324 26188 10376 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 2596 25984 2648 26036
rect 3976 25984 4028 26036
rect 5632 25984 5684 26036
rect 8760 26027 8812 26036
rect 8760 25993 8769 26027
rect 8769 25993 8803 26027
rect 8803 25993 8812 26027
rect 8760 25984 8812 25993
rect 5172 25916 5224 25968
rect 5540 25891 5592 25900
rect 5540 25857 5549 25891
rect 5549 25857 5583 25891
rect 5583 25857 5592 25891
rect 5540 25848 5592 25857
rect 5908 25848 5960 25900
rect 9312 25984 9364 26036
rect 3424 25780 3476 25832
rect 6828 25780 6880 25832
rect 8852 25780 8904 25832
rect 2780 25712 2832 25764
rect 5540 25712 5592 25764
rect 8760 25712 8812 25764
rect 9404 25755 9456 25764
rect 9404 25721 9416 25755
rect 9416 25721 9456 25755
rect 9404 25712 9456 25721
rect 2136 25687 2188 25696
rect 2136 25653 2145 25687
rect 2145 25653 2179 25687
rect 2179 25653 2188 25687
rect 2136 25644 2188 25653
rect 2964 25644 3016 25696
rect 5264 25644 5316 25696
rect 8484 25644 8536 25696
rect 10784 25644 10836 25696
rect 11244 25644 11296 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 2136 25440 2188 25492
rect 2872 25440 2924 25492
rect 5172 25483 5224 25492
rect 5172 25449 5181 25483
rect 5181 25449 5215 25483
rect 5215 25449 5224 25483
rect 5172 25440 5224 25449
rect 5540 25483 5592 25492
rect 5540 25449 5549 25483
rect 5549 25449 5583 25483
rect 5583 25449 5592 25483
rect 5540 25440 5592 25449
rect 8484 25483 8536 25492
rect 8484 25449 8493 25483
rect 8493 25449 8527 25483
rect 8527 25449 8536 25483
rect 8484 25440 8536 25449
rect 8852 25440 8904 25492
rect 2780 25372 2832 25424
rect 3424 25304 3476 25356
rect 4436 25347 4488 25356
rect 4436 25313 4445 25347
rect 4445 25313 4479 25347
rect 4479 25313 4488 25347
rect 4436 25304 4488 25313
rect 8668 25372 8720 25424
rect 5724 25304 5776 25356
rect 6092 25304 6144 25356
rect 8208 25304 8260 25356
rect 8760 25304 8812 25356
rect 4528 25279 4580 25288
rect 4528 25245 4537 25279
rect 4537 25245 4571 25279
rect 4571 25245 4580 25279
rect 4528 25236 4580 25245
rect 4620 25236 4672 25288
rect 5172 25236 5224 25288
rect 8668 25279 8720 25288
rect 8668 25245 8677 25279
rect 8677 25245 8711 25279
rect 8711 25245 8720 25279
rect 8668 25236 8720 25245
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 11244 25372 11296 25424
rect 10600 25347 10652 25356
rect 10600 25313 10634 25347
rect 10634 25313 10652 25347
rect 10600 25304 10652 25313
rect 10324 25236 10376 25245
rect 6184 25168 6236 25220
rect 7656 25168 7708 25220
rect 7288 25100 7340 25152
rect 9680 25100 9732 25152
rect 9864 25100 9916 25152
rect 10048 25143 10100 25152
rect 10048 25109 10057 25143
rect 10057 25109 10091 25143
rect 10091 25109 10100 25143
rect 10048 25100 10100 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4436 24896 4488 24948
rect 6092 24939 6144 24948
rect 6092 24905 6101 24939
rect 6101 24905 6135 24939
rect 6135 24905 6144 24939
rect 6092 24896 6144 24905
rect 8484 24896 8536 24948
rect 4620 24828 4672 24880
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 4528 24692 4580 24744
rect 8392 24760 8444 24812
rect 9404 24803 9456 24812
rect 9404 24769 9413 24803
rect 9413 24769 9447 24803
rect 9447 24769 9456 24803
rect 9404 24760 9456 24769
rect 9864 24760 9916 24812
rect 11428 24760 11480 24812
rect 4252 24624 4304 24676
rect 5448 24624 5500 24676
rect 2412 24556 2464 24608
rect 5172 24599 5224 24608
rect 5172 24565 5181 24599
rect 5181 24565 5215 24599
rect 5215 24565 5224 24599
rect 5172 24556 5224 24565
rect 6920 24556 6972 24608
rect 10416 24624 10468 24676
rect 11336 24624 11388 24676
rect 7196 24599 7248 24608
rect 7196 24565 7205 24599
rect 7205 24565 7239 24599
rect 7239 24565 7248 24599
rect 7196 24556 7248 24565
rect 7288 24556 7340 24608
rect 7656 24556 7708 24608
rect 8576 24556 8628 24608
rect 9496 24556 9548 24608
rect 10324 24599 10376 24608
rect 10324 24565 10333 24599
rect 10333 24565 10367 24599
rect 10367 24565 10376 24599
rect 10324 24556 10376 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 4436 24352 4488 24404
rect 4528 24352 4580 24404
rect 9404 24352 9456 24404
rect 9680 24395 9732 24404
rect 9680 24361 9689 24395
rect 9689 24361 9723 24395
rect 9723 24361 9732 24395
rect 9680 24352 9732 24361
rect 10600 24352 10652 24404
rect 3976 24216 4028 24268
rect 5540 24216 5592 24268
rect 6828 24216 6880 24268
rect 8668 24216 8720 24268
rect 9680 24216 9732 24268
rect 4252 24148 4304 24200
rect 5264 24191 5316 24200
rect 5264 24157 5273 24191
rect 5273 24157 5307 24191
rect 5307 24157 5316 24191
rect 5264 24148 5316 24157
rect 6184 24148 6236 24200
rect 5080 24080 5132 24132
rect 10324 24216 10376 24268
rect 10876 24216 10928 24268
rect 10784 24148 10836 24200
rect 10324 24080 10376 24132
rect 6920 24055 6972 24064
rect 6920 24021 6929 24055
rect 6929 24021 6963 24055
rect 6963 24021 6972 24055
rect 6920 24012 6972 24021
rect 11244 24012 11296 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 3976 23808 4028 23860
rect 4252 23851 4304 23860
rect 4252 23817 4261 23851
rect 4261 23817 4295 23851
rect 4295 23817 4304 23851
rect 4252 23808 4304 23817
rect 4804 23808 4856 23860
rect 5172 23808 5224 23860
rect 6184 23851 6236 23860
rect 6184 23817 6193 23851
rect 6193 23817 6227 23851
rect 6227 23817 6236 23851
rect 6184 23808 6236 23817
rect 5356 23740 5408 23792
rect 4804 23672 4856 23724
rect 6828 23808 6880 23860
rect 9864 23808 9916 23860
rect 10876 23808 10928 23860
rect 8024 23740 8076 23792
rect 8392 23672 8444 23724
rect 8668 23672 8720 23724
rect 9864 23672 9916 23724
rect 10784 23672 10836 23724
rect 6000 23604 6052 23656
rect 9680 23647 9732 23656
rect 9680 23613 9689 23647
rect 9689 23613 9723 23647
rect 9723 23613 9732 23647
rect 9680 23604 9732 23613
rect 10232 23604 10284 23656
rect 6920 23536 6972 23588
rect 7656 23536 7708 23588
rect 5172 23468 5224 23520
rect 7472 23468 7524 23520
rect 9588 23536 9640 23588
rect 10784 23536 10836 23588
rect 11060 23536 11112 23588
rect 8116 23468 8168 23520
rect 9312 23468 9364 23520
rect 10324 23511 10376 23520
rect 10324 23477 10333 23511
rect 10333 23477 10367 23511
rect 10367 23477 10376 23511
rect 10324 23468 10376 23477
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 5264 23264 5316 23316
rect 7196 23264 7248 23316
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 5172 23239 5224 23248
rect 5172 23205 5181 23239
rect 5181 23205 5215 23239
rect 5215 23205 5224 23239
rect 5172 23196 5224 23205
rect 5356 23196 5408 23248
rect 11336 23196 11388 23248
rect 4160 23060 4212 23112
rect 6184 23128 6236 23180
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 11244 23128 11296 23180
rect 8116 23060 8168 23112
rect 7840 22967 7892 22976
rect 7840 22933 7849 22967
rect 7849 22933 7883 22967
rect 7883 22933 7892 22967
rect 7840 22924 7892 22933
rect 8852 22924 8904 22976
rect 9312 22967 9364 22976
rect 9312 22933 9321 22967
rect 9321 22933 9355 22967
rect 9355 22933 9364 22967
rect 9312 22924 9364 22933
rect 10232 22967 10284 22976
rect 10232 22933 10241 22967
rect 10241 22933 10275 22967
rect 10275 22933 10284 22967
rect 10232 22924 10284 22933
rect 10600 22924 10652 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 5356 22720 5408 22772
rect 5540 22720 5592 22772
rect 7196 22720 7248 22772
rect 7472 22720 7524 22772
rect 8300 22763 8352 22772
rect 8300 22729 8309 22763
rect 8309 22729 8343 22763
rect 8343 22729 8352 22763
rect 8300 22720 8352 22729
rect 5724 22652 5776 22704
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 10048 22584 10100 22636
rect 3700 22516 3752 22568
rect 4160 22516 4212 22568
rect 7288 22516 7340 22568
rect 10232 22559 10284 22568
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 1676 22491 1728 22500
rect 1676 22457 1685 22491
rect 1685 22457 1719 22491
rect 1719 22457 1728 22491
rect 1676 22448 1728 22457
rect 3424 22423 3476 22432
rect 3424 22389 3433 22423
rect 3433 22389 3467 22423
rect 3467 22389 3476 22423
rect 3424 22380 3476 22389
rect 7012 22380 7064 22432
rect 7840 22423 7892 22432
rect 7840 22389 7849 22423
rect 7849 22389 7883 22423
rect 7883 22389 7892 22423
rect 7840 22380 7892 22389
rect 8116 22380 8168 22432
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 8668 22380 8720 22389
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 9864 22423 9916 22432
rect 9864 22389 9873 22423
rect 9873 22389 9907 22423
rect 9907 22389 9916 22423
rect 9864 22380 9916 22389
rect 11336 22380 11388 22432
rect 13360 22584 13412 22636
rect 12164 22448 12216 22500
rect 13084 22448 13136 22500
rect 11980 22380 12032 22432
rect 12808 22423 12860 22432
rect 12808 22389 12817 22423
rect 12817 22389 12851 22423
rect 12851 22389 12860 22423
rect 12808 22380 12860 22389
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 2412 22219 2464 22228
rect 2412 22185 2421 22219
rect 2421 22185 2455 22219
rect 2455 22185 2464 22219
rect 2412 22176 2464 22185
rect 5080 22219 5132 22228
rect 5080 22185 5089 22219
rect 5089 22185 5123 22219
rect 5123 22185 5132 22219
rect 5080 22176 5132 22185
rect 7288 22176 7340 22228
rect 8024 22219 8076 22228
rect 8024 22185 8033 22219
rect 8033 22185 8067 22219
rect 8067 22185 8076 22219
rect 8024 22176 8076 22185
rect 9404 22176 9456 22228
rect 10232 22176 10284 22228
rect 11980 22176 12032 22228
rect 12992 22176 13044 22228
rect 3700 22151 3752 22160
rect 2504 22040 2556 22092
rect 3700 22117 3709 22151
rect 3709 22117 3743 22151
rect 3743 22117 3752 22151
rect 3700 22108 3752 22117
rect 5540 22108 5592 22160
rect 7012 22108 7064 22160
rect 7564 22108 7616 22160
rect 10140 22108 10192 22160
rect 2688 22040 2740 22092
rect 3424 22040 3476 22092
rect 6184 22083 6236 22092
rect 6184 22049 6193 22083
rect 6193 22049 6227 22083
rect 6227 22049 6236 22083
rect 6184 22040 6236 22049
rect 8484 22040 8536 22092
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 2412 21904 2464 21956
rect 3240 21972 3292 22024
rect 11888 22108 11940 22160
rect 12808 22108 12860 22160
rect 5172 21972 5224 22024
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 10140 22015 10192 22024
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 10232 21972 10284 22024
rect 10600 21972 10652 22024
rect 10692 21972 10744 22024
rect 10876 21972 10928 22024
rect 12624 22040 12676 22092
rect 12900 22040 12952 22092
rect 12256 21972 12308 22024
rect 12440 21972 12492 22024
rect 13176 21972 13228 22024
rect 13360 21972 13412 22024
rect 13636 21972 13688 22024
rect 8208 21904 8260 21956
rect 11888 21904 11940 21956
rect 13084 21904 13136 21956
rect 1400 21836 1452 21888
rect 9864 21836 9916 21888
rect 10692 21879 10744 21888
rect 10692 21845 10701 21879
rect 10701 21845 10735 21879
rect 10735 21845 10744 21879
rect 10692 21836 10744 21845
rect 11244 21836 11296 21888
rect 13360 21836 13412 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 2412 21675 2464 21684
rect 2412 21641 2421 21675
rect 2421 21641 2455 21675
rect 2455 21641 2464 21675
rect 2412 21632 2464 21641
rect 3240 21632 3292 21684
rect 5724 21632 5776 21684
rect 7656 21675 7708 21684
rect 7656 21641 7665 21675
rect 7665 21641 7699 21675
rect 7699 21641 7708 21675
rect 7656 21632 7708 21641
rect 8116 21632 8168 21684
rect 8484 21675 8536 21684
rect 8484 21641 8493 21675
rect 8493 21641 8527 21675
rect 8527 21641 8536 21675
rect 8484 21632 8536 21641
rect 10048 21632 10100 21684
rect 10600 21632 10652 21684
rect 11980 21675 12032 21684
rect 11980 21641 11989 21675
rect 11989 21641 12023 21675
rect 12023 21641 12032 21675
rect 11980 21632 12032 21641
rect 12072 21632 12124 21684
rect 12348 21632 12400 21684
rect 12992 21675 13044 21684
rect 12992 21641 13001 21675
rect 13001 21641 13035 21675
rect 13035 21641 13044 21675
rect 12992 21632 13044 21641
rect 13176 21632 13228 21684
rect 13636 21675 13688 21684
rect 13636 21641 13645 21675
rect 13645 21641 13679 21675
rect 13679 21641 13688 21675
rect 13636 21632 13688 21641
rect 8024 21564 8076 21616
rect 9956 21564 10008 21616
rect 11888 21564 11940 21616
rect 2504 21539 2556 21548
rect 2504 21505 2513 21539
rect 2513 21505 2547 21539
rect 2547 21505 2556 21539
rect 2504 21496 2556 21505
rect 8392 21496 8444 21548
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 11336 21496 11388 21548
rect 12808 21496 12860 21548
rect 8668 21428 8720 21480
rect 2228 21360 2280 21412
rect 3148 21360 3200 21412
rect 10048 21360 10100 21412
rect 10600 21403 10652 21412
rect 10600 21369 10609 21403
rect 10609 21369 10643 21403
rect 10643 21369 10652 21403
rect 10600 21360 10652 21369
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 5172 21335 5224 21344
rect 5172 21301 5181 21335
rect 5181 21301 5215 21335
rect 5215 21301 5224 21335
rect 5172 21292 5224 21301
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 6092 21292 6144 21344
rect 9312 21292 9364 21344
rect 9864 21292 9916 21344
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 1676 21088 1728 21140
rect 2872 21088 2924 21140
rect 8668 21088 8720 21140
rect 10140 21088 10192 21140
rect 10692 21088 10744 21140
rect 12348 21131 12400 21140
rect 12348 21097 12357 21131
rect 12357 21097 12391 21131
rect 12391 21097 12400 21131
rect 12348 21088 12400 21097
rect 2964 21020 3016 21072
rect 4712 21020 4764 21072
rect 5448 21020 5500 21072
rect 9956 21063 10008 21072
rect 9956 21029 9965 21063
rect 9965 21029 9999 21063
rect 9999 21029 10008 21063
rect 9956 21020 10008 21029
rect 3056 20952 3108 21004
rect 4528 20995 4580 21004
rect 4528 20961 4537 20995
rect 4537 20961 4571 20995
rect 4571 20961 4580 20995
rect 4528 20952 4580 20961
rect 6184 20952 6236 21004
rect 6552 20952 6604 21004
rect 7840 20952 7892 21004
rect 9772 20952 9824 21004
rect 10416 20952 10468 21004
rect 10508 20952 10560 21004
rect 12072 20952 12124 21004
rect 4620 20927 4672 20936
rect 4620 20893 4629 20927
rect 4629 20893 4663 20927
rect 4663 20893 4672 20927
rect 4620 20884 4672 20893
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 10876 20927 10928 20936
rect 10876 20893 10885 20927
rect 10885 20893 10919 20927
rect 10919 20893 10928 20927
rect 10876 20884 10928 20893
rect 3148 20816 3200 20868
rect 11612 20816 11664 20868
rect 2688 20748 2740 20800
rect 7840 20791 7892 20800
rect 7840 20757 7849 20791
rect 7849 20757 7883 20791
rect 7883 20757 7892 20791
rect 7840 20748 7892 20757
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 2964 20544 3016 20596
rect 4528 20544 4580 20596
rect 5540 20544 5592 20596
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 11612 20587 11664 20596
rect 11612 20553 11621 20587
rect 11621 20553 11655 20587
rect 11655 20553 11664 20587
rect 11612 20544 11664 20553
rect 12348 20544 12400 20596
rect 2228 20519 2280 20528
rect 2228 20485 2237 20519
rect 2237 20485 2271 20519
rect 2271 20485 2280 20519
rect 2228 20476 2280 20485
rect 4620 20519 4672 20528
rect 4620 20485 4629 20519
rect 4629 20485 4663 20519
rect 4663 20485 4672 20519
rect 4620 20476 4672 20485
rect 6184 20476 6236 20528
rect 2504 20408 2556 20460
rect 11428 20408 11480 20460
rect 12072 20476 12124 20528
rect 8116 20340 8168 20392
rect 2872 20272 2924 20324
rect 8484 20272 8536 20324
rect 10048 20272 10100 20324
rect 4988 20204 5040 20256
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 10140 20204 10192 20256
rect 10508 20247 10560 20256
rect 10508 20213 10517 20247
rect 10517 20213 10551 20247
rect 10551 20213 10560 20247
rect 10508 20204 10560 20213
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 2504 20000 2556 20052
rect 4528 20043 4580 20052
rect 4528 20009 4537 20043
rect 4537 20009 4571 20043
rect 4571 20009 4580 20043
rect 4528 20000 4580 20009
rect 4896 20043 4948 20052
rect 4896 20009 4905 20043
rect 4905 20009 4939 20043
rect 4939 20009 4948 20043
rect 4896 20000 4948 20009
rect 6184 20000 6236 20052
rect 2872 19932 2924 19984
rect 3516 19932 3568 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 7288 19864 7340 19916
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 4252 19796 4304 19848
rect 5080 19839 5132 19848
rect 5080 19805 5089 19839
rect 5089 19805 5123 19839
rect 5123 19805 5132 19839
rect 5080 19796 5132 19805
rect 7104 19796 7156 19848
rect 7840 20000 7892 20052
rect 10416 20000 10468 20052
rect 10784 20000 10836 20052
rect 10876 20000 10928 20052
rect 10508 19932 10560 19984
rect 11428 19975 11480 19984
rect 11428 19941 11462 19975
rect 11462 19941 11480 19975
rect 11428 19932 11480 19941
rect 11244 19864 11296 19916
rect 10140 19796 10192 19848
rect 10876 19796 10928 19848
rect 5724 19728 5776 19780
rect 2688 19660 2740 19712
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 1400 19456 1452 19508
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 11060 19456 11112 19508
rect 11428 19456 11480 19508
rect 5448 19388 5500 19440
rect 10876 19388 10928 19440
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 5080 19320 5132 19372
rect 6184 19320 6236 19372
rect 3056 19252 3108 19304
rect 3332 19295 3384 19304
rect 3332 19261 3341 19295
rect 3341 19261 3375 19295
rect 3375 19261 3384 19295
rect 3332 19252 3384 19261
rect 4988 19295 5040 19304
rect 4988 19261 4997 19295
rect 4997 19261 5031 19295
rect 5031 19261 5040 19295
rect 4988 19252 5040 19261
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 7104 19295 7156 19304
rect 7104 19261 7138 19295
rect 7138 19261 7156 19295
rect 7104 19252 7156 19261
rect 9220 19252 9272 19304
rect 4896 19184 4948 19236
rect 6092 19184 6144 19236
rect 6828 19184 6880 19236
rect 3332 19116 3384 19168
rect 4252 19116 4304 19168
rect 4712 19116 4764 19168
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 5540 19116 5592 19168
rect 8208 19159 8260 19168
rect 8208 19125 8217 19159
rect 8217 19125 8251 19159
rect 8251 19125 8260 19159
rect 8208 19116 8260 19125
rect 8392 19116 8444 19168
rect 9404 19184 9456 19236
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 4988 18955 5040 18964
rect 4988 18921 4997 18955
rect 4997 18921 5031 18955
rect 5031 18921 5040 18955
rect 4988 18912 5040 18921
rect 5724 18955 5776 18964
rect 5724 18921 5733 18955
rect 5733 18921 5767 18955
rect 5767 18921 5776 18955
rect 5724 18912 5776 18921
rect 7104 18912 7156 18964
rect 9220 18912 9272 18964
rect 10416 18955 10468 18964
rect 10416 18921 10425 18955
rect 10425 18921 10459 18955
rect 10459 18921 10468 18955
rect 10416 18912 10468 18921
rect 10692 18912 10744 18964
rect 5080 18844 5132 18896
rect 5540 18776 5592 18828
rect 6092 18776 6144 18828
rect 10876 18776 10928 18828
rect 4712 18708 4764 18760
rect 7288 18708 7340 18760
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 3332 18572 3384 18624
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 7840 18572 7892 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 2780 18368 2832 18420
rect 4712 18411 4764 18420
rect 4712 18377 4721 18411
rect 4721 18377 4755 18411
rect 4755 18377 4764 18411
rect 4712 18368 4764 18377
rect 4988 18368 5040 18420
rect 6000 18368 6052 18420
rect 5540 18300 5592 18352
rect 6828 18300 6880 18352
rect 3148 18232 3200 18284
rect 3516 18232 3568 18284
rect 5264 18232 5316 18284
rect 3700 18164 3752 18216
rect 10692 18368 10744 18420
rect 11060 18368 11112 18420
rect 7288 18232 7340 18284
rect 8208 18232 8260 18284
rect 5632 18096 5684 18148
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 4528 18028 4580 18080
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 6092 18028 6144 18080
rect 7104 18028 7156 18080
rect 8024 18028 8076 18080
rect 8300 18028 8352 18080
rect 9312 18028 9364 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 5448 17867 5500 17876
rect 5448 17833 5457 17867
rect 5457 17833 5491 17867
rect 5491 17833 5500 17867
rect 5448 17824 5500 17833
rect 5724 17824 5776 17876
rect 7288 17867 7340 17876
rect 7288 17833 7297 17867
rect 7297 17833 7331 17867
rect 7331 17833 7340 17867
rect 7288 17824 7340 17833
rect 8300 17756 8352 17808
rect 10232 17756 10284 17808
rect 4344 17731 4396 17740
rect 4344 17697 4378 17731
rect 4378 17697 4396 17731
rect 4344 17688 4396 17697
rect 9680 17688 9732 17740
rect 10416 17688 10468 17740
rect 3240 17620 3292 17672
rect 8484 17620 8536 17672
rect 9956 17620 10008 17672
rect 7104 17484 7156 17536
rect 7748 17484 7800 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 3516 17280 3568 17332
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 5632 17323 5684 17332
rect 5632 17289 5641 17323
rect 5641 17289 5675 17323
rect 5675 17289 5684 17323
rect 5632 17280 5684 17289
rect 8300 17280 8352 17332
rect 9680 17280 9732 17332
rect 10508 17280 10560 17332
rect 11152 17212 11204 17264
rect 11980 17212 12032 17264
rect 3976 17144 4028 17196
rect 4344 17187 4396 17196
rect 4344 17153 4353 17187
rect 4353 17153 4387 17187
rect 4387 17153 4396 17187
rect 4344 17144 4396 17153
rect 3976 17008 4028 17060
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 8392 17144 8444 17196
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 8300 17076 8352 17128
rect 9956 17144 10008 17196
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 7564 17008 7616 17060
rect 5448 16940 5500 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 9404 16983 9456 16992
rect 9404 16949 9413 16983
rect 9413 16949 9447 16983
rect 9447 16949 9456 16983
rect 9404 16940 9456 16949
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 3976 16736 4028 16788
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 5540 16736 5592 16788
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 8484 16736 8536 16788
rect 9312 16736 9364 16788
rect 1676 16711 1728 16720
rect 1676 16677 1685 16711
rect 1685 16677 1719 16711
rect 1719 16677 1728 16711
rect 1676 16668 1728 16677
rect 2872 16668 2924 16720
rect 7748 16668 7800 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 5080 16643 5132 16652
rect 5080 16609 5089 16643
rect 5089 16609 5123 16643
rect 5123 16609 5132 16643
rect 5080 16600 5132 16609
rect 6828 16600 6880 16652
rect 7932 16643 7984 16652
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 8024 16643 8076 16652
rect 8024 16609 8033 16643
rect 8033 16609 8067 16643
rect 8067 16609 8076 16643
rect 8024 16600 8076 16609
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 11612 16600 11664 16652
rect 8484 16532 8536 16584
rect 9588 16532 9640 16584
rect 2780 16464 2832 16516
rect 9956 16507 10008 16516
rect 9956 16473 9965 16507
rect 9965 16473 9999 16507
rect 9999 16473 10008 16507
rect 9956 16464 10008 16473
rect 10324 16464 10376 16516
rect 4528 16396 4580 16448
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 1400 16192 1452 16244
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 2780 16192 2832 16201
rect 5540 16192 5592 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 9312 16192 9364 16244
rect 9496 16192 9548 16244
rect 10692 16192 10744 16244
rect 11152 16192 11204 16244
rect 3240 15988 3292 16040
rect 3976 15988 4028 16040
rect 6828 15988 6880 16040
rect 8760 15988 8812 16040
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 9864 16031 9916 16040
rect 9864 15997 9898 16031
rect 9898 15997 9916 16031
rect 9864 15988 9916 15997
rect 4528 15963 4580 15972
rect 4528 15929 4562 15963
rect 4562 15929 4580 15963
rect 4528 15920 4580 15929
rect 7380 15963 7432 15972
rect 7380 15929 7414 15963
rect 7414 15929 7432 15963
rect 7380 15920 7432 15929
rect 11612 15963 11664 15972
rect 11612 15929 11621 15963
rect 11621 15929 11655 15963
rect 11655 15929 11664 15963
rect 11612 15920 11664 15929
rect 12256 15920 12308 15972
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 4160 15895 4212 15904
rect 4160 15861 4169 15895
rect 4169 15861 4203 15895
rect 4203 15861 4212 15895
rect 4160 15852 4212 15861
rect 5264 15852 5316 15904
rect 7932 15852 7984 15904
rect 9496 15852 9548 15904
rect 11060 15852 11112 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 7288 15648 7340 15700
rect 7932 15648 7984 15700
rect 8300 15648 8352 15700
rect 8668 15648 8720 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10048 15648 10100 15700
rect 11060 15648 11112 15700
rect 7472 15580 7524 15632
rect 4160 15512 4212 15564
rect 7380 15512 7432 15564
rect 9680 15512 9732 15564
rect 3976 15444 4028 15496
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 9588 15444 9640 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11520 15512 11572 15564
rect 8760 15308 8812 15360
rect 12256 15308 12308 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 5080 15104 5132 15156
rect 7472 15104 7524 15156
rect 7656 15104 7708 15156
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 10324 15104 10376 15156
rect 11520 15147 11572 15156
rect 11520 15113 11529 15147
rect 11529 15113 11563 15147
rect 11563 15113 11572 15147
rect 11520 15104 11572 15113
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 4528 14968 4580 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 12900 15036 12952 15088
rect 13084 15036 13136 15088
rect 7288 14968 7340 15020
rect 12716 14968 12768 15020
rect 6552 14900 6604 14952
rect 8300 14900 8352 14952
rect 8760 14900 8812 14952
rect 12164 14900 12216 14952
rect 9036 14875 9088 14884
rect 9036 14841 9045 14875
rect 9045 14841 9079 14875
rect 9079 14841 9088 14875
rect 9036 14832 9088 14841
rect 9496 14832 9548 14884
rect 12808 14875 12860 14884
rect 12808 14841 12817 14875
rect 12817 14841 12851 14875
rect 12851 14841 12860 14875
rect 12808 14832 12860 14841
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 5264 14764 5316 14816
rect 5724 14764 5776 14816
rect 9220 14764 9272 14816
rect 12164 14764 12216 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 5816 14560 5868 14612
rect 8208 14560 8260 14612
rect 9036 14560 9088 14612
rect 9588 14560 9640 14612
rect 12164 14560 12216 14612
rect 12716 14603 12768 14612
rect 12716 14569 12725 14603
rect 12725 14569 12759 14603
rect 12759 14569 12768 14603
rect 12716 14560 12768 14569
rect 12808 14560 12860 14612
rect 1676 14535 1728 14544
rect 1676 14501 1685 14535
rect 1685 14501 1719 14535
rect 1719 14501 1728 14535
rect 1676 14492 1728 14501
rect 6184 14467 6236 14476
rect 6184 14433 6218 14467
rect 6218 14433 6236 14467
rect 6184 14424 6236 14433
rect 7288 14424 7340 14476
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 1676 14356 1728 14408
rect 5540 14356 5592 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 9680 14288 9732 14340
rect 10324 14288 10376 14340
rect 10508 14288 10560 14340
rect 5264 14263 5316 14272
rect 5264 14229 5273 14263
rect 5273 14229 5307 14263
rect 5307 14229 5316 14263
rect 5264 14220 5316 14229
rect 10140 14263 10192 14272
rect 10140 14229 10149 14263
rect 10149 14229 10183 14263
rect 10183 14229 10192 14263
rect 10140 14220 10192 14229
rect 11060 14220 11112 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 5264 14016 5316 14068
rect 7472 14016 7524 14068
rect 8116 14016 8168 14068
rect 1676 13991 1728 14000
rect 1676 13957 1685 13991
rect 1685 13957 1719 13991
rect 1719 13957 1728 13991
rect 1676 13948 1728 13957
rect 5632 13948 5684 14000
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 7196 13880 7248 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 9588 14016 9640 14068
rect 10600 14059 10652 14068
rect 10600 14025 10609 14059
rect 10609 14025 10643 14059
rect 10643 14025 10652 14059
rect 10600 14016 10652 14025
rect 10692 14016 10744 14068
rect 11520 14016 11572 14068
rect 8668 13948 8720 14000
rect 9128 13948 9180 14000
rect 7380 13880 7432 13889
rect 9496 13880 9548 13932
rect 10692 13880 10744 13932
rect 12164 14016 12216 14068
rect 12716 13880 12768 13932
rect 9312 13744 9364 13796
rect 11060 13812 11112 13864
rect 13084 13812 13136 13864
rect 10876 13676 10928 13728
rect 12992 13744 13044 13796
rect 13820 13744 13872 13796
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 7196 13472 7248 13524
rect 8668 13472 8720 13524
rect 9312 13472 9364 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 11060 13472 11112 13524
rect 11428 13472 11480 13524
rect 12992 13472 13044 13524
rect 13360 13472 13412 13524
rect 10600 13404 10652 13456
rect 12256 13404 12308 13456
rect 12808 13404 12860 13456
rect 13084 13404 13136 13456
rect 11244 13268 11296 13320
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 3424 13132 3476 13184
rect 4068 13132 4120 13184
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 8300 13132 8352 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 10508 12928 10560 12980
rect 11428 12928 11480 12980
rect 11520 12928 11572 12980
rect 12256 12860 12308 12912
rect 10324 12792 10376 12844
rect 10508 12792 10560 12844
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8208 12699 8260 12708
rect 8208 12665 8220 12699
rect 8220 12665 8260 12699
rect 8208 12656 8260 12665
rect 11244 12656 11296 12708
rect 11428 12656 11480 12708
rect 9496 12588 9548 12640
rect 11520 12588 11572 12640
rect 12624 12588 12676 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 5632 12384 5684 12436
rect 5816 12384 5868 12436
rect 9772 12384 9824 12436
rect 9864 12384 9916 12436
rect 8300 12316 8352 12368
rect 8668 12316 8720 12368
rect 10232 12316 10284 12368
rect 10692 12316 10744 12368
rect 11152 12316 11204 12368
rect 4620 12291 4672 12300
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 9588 12248 9640 12300
rect 9864 12248 9916 12300
rect 11244 12248 11296 12300
rect 4252 12180 4304 12232
rect 4344 12180 4396 12232
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 5724 12180 5776 12232
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 8208 12112 8260 12164
rect 8760 12180 8812 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 11152 12223 11204 12232
rect 10048 12155 10100 12164
rect 10048 12121 10057 12155
rect 10057 12121 10091 12155
rect 10091 12121 10100 12155
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 10048 12112 10100 12121
rect 4068 12044 4120 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 12624 12044 12676 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 4896 11840 4948 11892
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 7932 11840 7984 11892
rect 8576 11840 8628 11892
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 9956 11815 10008 11824
rect 9956 11781 9965 11815
rect 9965 11781 9999 11815
rect 9999 11781 10008 11815
rect 9956 11772 10008 11781
rect 4252 11679 4304 11688
rect 4252 11645 4261 11679
rect 4261 11645 4295 11679
rect 4295 11645 4304 11679
rect 4252 11636 4304 11645
rect 12164 11747 12216 11756
rect 4528 11679 4580 11688
rect 4528 11645 4551 11679
rect 4551 11645 4580 11679
rect 4528 11636 4580 11645
rect 10508 11636 10560 11688
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 12624 11704 12676 11756
rect 12532 11636 12584 11688
rect 13084 11636 13136 11688
rect 2228 11611 2280 11620
rect 2228 11577 2237 11611
rect 2237 11577 2271 11611
rect 2271 11577 2280 11611
rect 2228 11568 2280 11577
rect 4344 11568 4396 11620
rect 5724 11500 5776 11552
rect 10048 11568 10100 11620
rect 8760 11500 8812 11552
rect 9956 11500 10008 11552
rect 11060 11500 11112 11552
rect 12164 11500 12216 11552
rect 13728 11500 13780 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 4252 11296 4304 11348
rect 7748 11339 7800 11348
rect 4620 11228 4672 11280
rect 7748 11305 7757 11339
rect 7757 11305 7791 11339
rect 7791 11305 7800 11339
rect 7748 11296 7800 11305
rect 8024 11296 8076 11348
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 5448 11228 5500 11280
rect 6828 11228 6880 11280
rect 7932 11228 7984 11280
rect 8484 11296 8536 11348
rect 9496 11296 9548 11348
rect 9956 11296 10008 11348
rect 11244 11296 11296 11348
rect 12624 11296 12676 11348
rect 8576 11228 8628 11280
rect 5724 11160 5776 11212
rect 8208 11135 8260 11144
rect 3332 10956 3384 11008
rect 3976 10956 4028 11008
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 7932 11024 7984 11076
rect 9588 11092 9640 11144
rect 11152 11228 11204 11280
rect 9956 11203 10008 11212
rect 9956 11169 9990 11203
rect 9990 11169 10008 11203
rect 9956 11160 10008 11169
rect 6460 10999 6512 11008
rect 6460 10965 6469 10999
rect 6469 10965 6503 10999
rect 6503 10965 6512 10999
rect 6460 10956 6512 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 4620 10752 4672 10804
rect 5540 10752 5592 10804
rect 8576 10752 8628 10804
rect 9588 10752 9640 10804
rect 10968 10752 11020 10804
rect 6460 10684 6512 10736
rect 4528 10616 4580 10668
rect 7932 10684 7984 10736
rect 9956 10684 10008 10736
rect 10692 10684 10744 10736
rect 3056 10548 3108 10600
rect 4068 10548 4120 10600
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 10784 10616 10836 10668
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 5080 10480 5132 10532
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 4896 10412 4948 10421
rect 5724 10412 5776 10464
rect 7564 10412 7616 10464
rect 9588 10412 9640 10464
rect 10600 10412 10652 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 3332 10208 3384 10260
rect 6000 10208 6052 10260
rect 6644 10208 6696 10260
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 7380 10140 7432 10192
rect 8116 10140 8168 10192
rect 9680 10208 9732 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 10232 10208 10284 10260
rect 10784 10251 10836 10260
rect 10784 10217 10793 10251
rect 10793 10217 10827 10251
rect 10827 10217 10836 10251
rect 10784 10208 10836 10217
rect 9864 10140 9916 10192
rect 3148 10072 3200 10124
rect 3332 10072 3384 10124
rect 4988 10072 5040 10124
rect 8576 10072 8628 10124
rect 4160 10004 4212 10056
rect 5080 10004 5132 10056
rect 5172 10004 5224 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 10508 10004 10560 10056
rect 9772 9936 9824 9988
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 4528 9664 4580 9716
rect 5724 9664 5776 9716
rect 8300 9664 8352 9716
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 3332 9596 3384 9648
rect 5448 9596 5500 9648
rect 9772 9639 9824 9648
rect 9772 9605 9781 9639
rect 9781 9605 9815 9639
rect 9815 9605 9824 9639
rect 9772 9596 9824 9605
rect 10232 9596 10284 9648
rect 4528 9528 4580 9580
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 7104 9528 7156 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 8760 9528 8812 9580
rect 4712 9503 4764 9512
rect 4712 9469 4721 9503
rect 4721 9469 4755 9503
rect 4755 9469 4764 9503
rect 4712 9460 4764 9469
rect 6828 9460 6880 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 8392 9460 8444 9512
rect 8668 9460 8720 9512
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 6920 9392 6972 9444
rect 5816 9324 5868 9376
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 7104 9324 7156 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 7932 9324 7984 9376
rect 8668 9324 8720 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 5172 9120 5224 9172
rect 7472 9120 7524 9172
rect 8576 9120 8628 9172
rect 5540 9052 5592 9104
rect 6644 9052 6696 9104
rect 7104 9052 7156 9104
rect 7564 9052 7616 9104
rect 4436 8984 4488 9036
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 6736 8959 6788 8968
rect 4528 8848 4580 8900
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 3976 8780 4028 8832
rect 8116 8823 8168 8832
rect 8116 8789 8125 8823
rect 8125 8789 8159 8823
rect 8159 8789 8168 8823
rect 8116 8780 8168 8789
rect 8300 8780 8352 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 10416 8780 10468 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 4988 8576 5040 8628
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 6184 8483 6236 8492
rect 5724 8440 5776 8449
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7012 8440 7064 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8116 8440 8168 8492
rect 2504 8372 2556 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 6644 8415 6696 8424
rect 5632 8372 5684 8381
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 7288 8415 7340 8424
rect 6644 8372 6696 8381
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 9404 8576 9456 8628
rect 10600 8483 10652 8492
rect 9864 8372 9916 8424
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10968 8372 11020 8424
rect 2596 8304 2648 8356
rect 10416 8347 10468 8356
rect 10416 8313 10425 8347
rect 10425 8313 10459 8347
rect 10459 8313 10468 8347
rect 10416 8304 10468 8313
rect 3516 8236 3568 8288
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 8484 8236 8536 8288
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 9036 8236 9088 8288
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 4528 8032 4580 8084
rect 4804 8075 4856 8084
rect 4804 8041 4813 8075
rect 4813 8041 4847 8075
rect 4847 8041 4856 8075
rect 4804 8032 4856 8041
rect 6184 8032 6236 8084
rect 7104 8032 7156 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8300 8032 8352 8084
rect 9036 8075 9088 8084
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 10140 8032 10192 8084
rect 10600 8032 10652 8084
rect 1676 8007 1728 8016
rect 1676 7973 1685 8007
rect 1685 7973 1719 8007
rect 1719 7973 1728 8007
rect 1676 7964 1728 7973
rect 7564 7964 7616 8016
rect 9864 7964 9916 8016
rect 2412 7896 2464 7948
rect 5264 7939 5316 7948
rect 5264 7905 5298 7939
rect 5298 7905 5316 7939
rect 5264 7896 5316 7905
rect 7840 7896 7892 7948
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 11796 7896 11848 7948
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8300 7760 8352 7812
rect 9588 7828 9640 7880
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 3424 7692 3476 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 3056 7488 3108 7540
rect 3516 7488 3568 7540
rect 7840 7488 7892 7540
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 12440 7488 12492 7540
rect 5632 7420 5684 7472
rect 7380 7463 7432 7472
rect 3516 7327 3568 7336
rect 3516 7293 3550 7327
rect 3550 7293 3568 7327
rect 3516 7284 3568 7293
rect 7380 7429 7389 7463
rect 7389 7429 7423 7463
rect 7423 7429 7432 7463
rect 7380 7420 7432 7429
rect 6736 7284 6788 7336
rect 9404 7352 9456 7404
rect 3424 7216 3476 7268
rect 4988 7216 5040 7268
rect 5908 7216 5960 7268
rect 9588 7284 9640 7336
rect 10140 7327 10192 7336
rect 10140 7293 10174 7327
rect 10174 7293 10192 7327
rect 1400 7148 1452 7200
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 5264 7148 5316 7200
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 8024 7148 8076 7200
rect 10140 7284 10192 7293
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 10968 7148 11020 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 4804 6944 4856 6996
rect 5080 6944 5132 6996
rect 6828 6944 6880 6996
rect 8484 6944 8536 6996
rect 9588 6944 9640 6996
rect 11980 6944 12032 6996
rect 6736 6876 6788 6928
rect 8300 6876 8352 6928
rect 8392 6919 8444 6928
rect 8392 6885 8401 6919
rect 8401 6885 8435 6919
rect 8435 6885 8444 6919
rect 8392 6876 8444 6885
rect 8944 6876 8996 6928
rect 12624 6919 12676 6928
rect 12624 6885 12633 6919
rect 12633 6885 12667 6919
rect 12667 6885 12676 6919
rect 12624 6876 12676 6885
rect 1584 6808 1636 6860
rect 3976 6808 4028 6860
rect 5448 6808 5500 6860
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 2596 6740 2648 6792
rect 4896 6740 4948 6792
rect 4620 6672 4672 6724
rect 6644 6740 6696 6792
rect 8208 6740 8260 6792
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 9404 6808 9456 6860
rect 9956 6851 10008 6860
rect 9956 6817 9990 6851
rect 9990 6817 10008 6851
rect 9956 6808 10008 6817
rect 10968 6808 11020 6860
rect 9588 6740 9640 6792
rect 11060 6740 11112 6792
rect 12716 6783 12768 6792
rect 5448 6672 5500 6724
rect 8944 6672 8996 6724
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 13360 6740 13412 6792
rect 12440 6672 12492 6724
rect 940 6604 992 6656
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 3424 6604 3476 6656
rect 7748 6604 7800 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12808 6604 12860 6656
rect 13636 6604 13688 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2044 6400 2096 6452
rect 5080 6400 5132 6452
rect 5448 6443 5500 6452
rect 5448 6409 5457 6443
rect 5457 6409 5491 6443
rect 5491 6409 5500 6443
rect 5448 6400 5500 6409
rect 6736 6400 6788 6452
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 1492 6264 1544 6316
rect 2412 6196 2464 6248
rect 5264 6332 5316 6384
rect 5540 6332 5592 6384
rect 8760 6332 8812 6384
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 7564 6264 7616 6316
rect 9956 6400 10008 6452
rect 11244 6400 11296 6452
rect 13360 6400 13412 6452
rect 5172 6196 5224 6248
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 7840 6196 7892 6248
rect 8484 6196 8536 6248
rect 9496 6196 9548 6248
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 12532 6196 12584 6248
rect 12808 6196 12860 6248
rect 1584 6128 1636 6180
rect 2320 6128 2372 6180
rect 2412 6060 2464 6112
rect 2596 6060 2648 6112
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 4988 6128 5040 6180
rect 7748 6128 7800 6180
rect 9312 6128 9364 6180
rect 9588 6128 9640 6180
rect 11060 6128 11112 6180
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 9680 6060 9732 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 12624 6128 12676 6180
rect 12532 6060 12584 6112
rect 13360 6060 13412 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 2780 5856 2832 5908
rect 4344 5856 4396 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 5264 5856 5316 5908
rect 2964 5788 3016 5840
rect 6092 5788 6144 5840
rect 6644 5856 6696 5908
rect 6920 5856 6972 5908
rect 8392 5856 8444 5908
rect 9312 5856 9364 5908
rect 11336 5856 11388 5908
rect 12164 5856 12216 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 2872 5720 2924 5772
rect 4068 5763 4120 5772
rect 4068 5729 4077 5763
rect 4077 5729 4111 5763
rect 4111 5729 4120 5763
rect 4068 5720 4120 5729
rect 5540 5763 5592 5772
rect 5540 5729 5549 5763
rect 5549 5729 5583 5763
rect 5583 5729 5592 5763
rect 5540 5720 5592 5729
rect 5908 5720 5960 5772
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 8392 5720 8444 5772
rect 8852 5720 8904 5772
rect 9772 5720 9824 5772
rect 13268 5763 13320 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 7288 5695 7340 5704
rect 3148 5584 3200 5636
rect 5080 5584 5132 5636
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 11796 5652 11848 5704
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 10048 5584 10100 5636
rect 11980 5584 12032 5636
rect 2136 5516 2188 5568
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 10600 5559 10652 5568
rect 10600 5525 10609 5559
rect 10609 5525 10643 5559
rect 10643 5525 10652 5559
rect 10600 5516 10652 5525
rect 11336 5516 11388 5568
rect 12808 5652 12860 5704
rect 12808 5516 12860 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 2872 5312 2924 5364
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 5908 5287 5960 5296
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 5908 5253 5917 5287
rect 5917 5253 5951 5287
rect 5951 5253 5960 5287
rect 5908 5244 5960 5253
rect 3056 5176 3108 5228
rect 3424 5176 3476 5228
rect 2688 5108 2740 5160
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 5080 5040 5132 5092
rect 7288 5176 7340 5228
rect 9404 5312 9456 5364
rect 9588 5312 9640 5364
rect 9772 5312 9824 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 12900 5312 12952 5364
rect 13268 5312 13320 5364
rect 11336 5176 11388 5228
rect 12900 5108 12952 5160
rect 7564 5040 7616 5092
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 10508 5015 10560 5024
rect 10508 4981 10517 5015
rect 10517 4981 10551 5015
rect 10551 4981 10560 5015
rect 10508 4972 10560 4981
rect 10600 5015 10652 5024
rect 10600 4981 10609 5015
rect 10609 4981 10643 5015
rect 10643 4981 10652 5015
rect 11336 5015 11388 5024
rect 10600 4972 10652 4981
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 4160 4768 4212 4820
rect 4988 4768 5040 4820
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 6736 4768 6788 4820
rect 6920 4768 6972 4820
rect 7656 4768 7708 4820
rect 8116 4768 8168 4820
rect 10140 4768 10192 4820
rect 11060 4811 11112 4820
rect 11060 4777 11069 4811
rect 11069 4777 11103 4811
rect 11103 4777 11112 4811
rect 11060 4768 11112 4777
rect 2504 4700 2556 4752
rect 4896 4743 4948 4752
rect 4896 4709 4905 4743
rect 4905 4709 4939 4743
rect 4939 4709 4948 4743
rect 4896 4700 4948 4709
rect 5448 4700 5500 4752
rect 7104 4700 7156 4752
rect 8392 4700 8444 4752
rect 3148 4632 3200 4684
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 4804 4632 4856 4641
rect 5724 4632 5776 4684
rect 7012 4632 7064 4684
rect 8208 4632 8260 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 11336 4632 11388 4684
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 5080 4607 5132 4616
rect 2504 4496 2556 4548
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 9680 4564 9732 4616
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11060 4564 11112 4616
rect 7564 4539 7616 4548
rect 7564 4505 7573 4539
rect 7573 4505 7607 4539
rect 7607 4505 7616 4539
rect 7564 4496 7616 4505
rect 3516 4471 3568 4480
rect 3516 4437 3525 4471
rect 3525 4437 3559 4471
rect 3559 4437 3568 4471
rect 3516 4428 3568 4437
rect 4068 4428 4120 4480
rect 7472 4428 7524 4480
rect 10508 4428 10560 4480
rect 10692 4428 10744 4480
rect 12716 4428 12768 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2320 4267 2372 4276
rect 2320 4233 2329 4267
rect 2329 4233 2363 4267
rect 2363 4233 2372 4267
rect 2320 4224 2372 4233
rect 2872 4224 2924 4276
rect 5080 4224 5132 4276
rect 6552 4224 6604 4276
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 10324 4224 10376 4276
rect 11060 4224 11112 4276
rect 3516 4156 3568 4208
rect 3608 4156 3660 4208
rect 4068 4156 4120 4208
rect 4896 4156 4948 4208
rect 3056 4088 3108 4140
rect 6920 4156 6972 4208
rect 8116 4156 8168 4208
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 12992 4131 13044 4140
rect 1952 4020 2004 4072
rect 3516 4020 3568 4072
rect 8484 4020 8536 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 10140 4020 10192 4072
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 1676 3995 1728 4004
rect 1676 3961 1685 3995
rect 1685 3961 1719 3995
rect 1719 3961 1728 3995
rect 1676 3952 1728 3961
rect 2320 3952 2372 4004
rect 3884 3995 3936 4004
rect 3884 3961 3893 3995
rect 3893 3961 3927 3995
rect 3927 3961 3936 3995
rect 3884 3952 3936 3961
rect 3332 3884 3384 3936
rect 6092 3884 6144 3936
rect 8392 3952 8444 4004
rect 9588 3952 9640 4004
rect 10416 3884 10468 3936
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 3608 3680 3660 3732
rect 4068 3680 4120 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6736 3680 6788 3732
rect 7288 3680 7340 3732
rect 9588 3680 9640 3732
rect 10508 3680 10560 3732
rect 10692 3680 10744 3732
rect 11336 3680 11388 3732
rect 572 3612 624 3664
rect 1308 3612 1360 3664
rect 2780 3655 2832 3664
rect 2780 3621 2789 3655
rect 2789 3621 2823 3655
rect 2823 3621 2832 3655
rect 2780 3612 2832 3621
rect 5816 3612 5868 3664
rect 6368 3612 6420 3664
rect 6920 3612 6972 3664
rect 3516 3544 3568 3596
rect 5264 3544 5316 3596
rect 9588 3544 9640 3596
rect 10232 3544 10284 3596
rect 11060 3587 11112 3596
rect 11060 3553 11069 3587
rect 11069 3553 11103 3587
rect 11103 3553 11112 3587
rect 11060 3544 11112 3553
rect 11152 3544 11204 3596
rect 12532 3544 12584 3596
rect 13176 3544 13228 3596
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 12716 3476 12768 3528
rect 1860 3408 1912 3460
rect 2596 3408 2648 3460
rect 8300 3451 8352 3460
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 9404 3408 9456 3460
rect 9772 3408 9824 3460
rect 10232 3408 10284 3460
rect 3056 3340 3108 3392
rect 4252 3340 4304 3392
rect 8484 3340 8536 3392
rect 10140 3340 10192 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2872 3136 2924 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 5080 3136 5132 3188
rect 5448 3179 5500 3188
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 7196 3136 7248 3188
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 9588 3179 9640 3188
rect 2596 3068 2648 3120
rect 3240 3068 3292 3120
rect 4068 3068 4120 3120
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3424 3000 3476 3052
rect 9588 3145 9597 3179
rect 9597 3145 9631 3179
rect 9631 3145 9640 3179
rect 9588 3136 9640 3145
rect 11428 3136 11480 3188
rect 12440 3179 12492 3188
rect 11152 3068 11204 3120
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 12716 3068 12768 3120
rect 3976 2932 4028 2984
rect 6276 2932 6328 2984
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 7288 2932 7340 2984
rect 13452 3000 13504 3052
rect 13820 3000 13872 3052
rect 14924 3000 14976 3052
rect 4620 2864 4672 2916
rect 5080 2864 5132 2916
rect 12716 2932 12768 2984
rect 11060 2864 11112 2916
rect 11428 2864 11480 2916
rect 13728 2932 13780 2984
rect 204 2796 256 2848
rect 1768 2796 1820 2848
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13452 2796 13504 2805
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 3056 2592 3108 2644
rect 3976 2592 4028 2644
rect 4712 2592 4764 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 7196 2635 7248 2644
rect 7196 2601 7205 2635
rect 7205 2601 7239 2635
rect 7239 2601 7248 2635
rect 8484 2635 8536 2644
rect 7196 2592 7248 2601
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 8576 2592 8628 2644
rect 9680 2592 9732 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 4252 2524 4304 2576
rect 9496 2524 9548 2576
rect 10140 2524 10192 2576
rect 10784 2524 10836 2576
rect 12164 2524 12216 2576
rect 1400 2456 1452 2508
rect 1768 2499 1820 2508
rect 1768 2465 1791 2499
rect 1791 2465 1820 2499
rect 1768 2456 1820 2465
rect 5448 2388 5500 2440
rect 8024 2499 8076 2508
rect 8024 2465 8033 2499
rect 8033 2465 8067 2499
rect 8067 2465 8076 2499
rect 8024 2456 8076 2465
rect 9772 2456 9824 2508
rect 11888 2456 11940 2508
rect 9956 2388 10008 2440
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 11152 2388 11204 2440
rect 13452 2388 13504 2440
rect 3148 2320 3200 2372
rect 6276 2363 6328 2372
rect 6276 2329 6285 2363
rect 6285 2329 6319 2363
rect 6319 2329 6328 2363
rect 6276 2320 6328 2329
rect 9772 2320 9824 2372
rect 10232 2320 10284 2372
rect 3424 2252 3476 2304
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 7656 2295 7708 2304
rect 7656 2261 7665 2295
rect 7665 2261 7699 2295
rect 7699 2261 7708 2295
rect 7656 2252 7708 2261
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 5724 1232 5776 1284
rect 7840 1232 7892 1284
rect 6920 552 6972 604
rect 7104 552 7156 604
rect 9956 552 10008 604
rect 10140 552 10192 604
rect 10600 552 10652 604
rect 10876 552 10928 604
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39520 10654 40000
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39520 14242 40000
rect 14554 39520 14610 40000
rect 14922 39522 14978 40000
rect 14922 39520 15056 39522
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 35290 244 39520
rect 584 35834 612 39520
rect 572 35828 624 35834
rect 572 35770 624 35776
rect 204 35284 256 35290
rect 204 35226 256 35232
rect 952 30666 980 39520
rect 1412 33658 1440 39520
rect 1582 38720 1638 38729
rect 1582 38655 1638 38664
rect 1490 34640 1546 34649
rect 1596 34610 1624 38655
rect 1674 36408 1730 36417
rect 1674 36343 1730 36352
rect 1490 34575 1546 34584
rect 1584 34604 1636 34610
rect 1504 34066 1532 34575
rect 1584 34546 1636 34552
rect 1688 34134 1716 36343
rect 1780 34202 1808 39520
rect 2148 35290 2176 39520
rect 2608 35834 2636 39520
rect 2596 35828 2648 35834
rect 2596 35770 2648 35776
rect 2976 35601 3004 39520
rect 3344 35737 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4016 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3988 35834 4016 37182
rect 3976 35828 4028 35834
rect 3976 35770 4028 35776
rect 3330 35728 3386 35737
rect 3330 35663 3386 35672
rect 3240 35624 3292 35630
rect 2962 35592 3018 35601
rect 3240 35566 3292 35572
rect 2962 35527 3018 35536
rect 2228 35488 2280 35494
rect 2228 35430 2280 35436
rect 2136 35284 2188 35290
rect 2136 35226 2188 35232
rect 1860 35148 1912 35154
rect 1860 35090 1912 35096
rect 1872 34678 1900 35090
rect 2044 34944 2096 34950
rect 2044 34886 2096 34892
rect 1860 34672 1912 34678
rect 1860 34614 1912 34620
rect 2056 34542 2084 34886
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 1768 34196 1820 34202
rect 1768 34138 1820 34144
rect 1676 34128 1728 34134
rect 1582 34096 1638 34105
rect 1492 34060 1544 34066
rect 1676 34070 1728 34076
rect 1582 34031 1638 34040
rect 1492 34002 1544 34008
rect 1400 33652 1452 33658
rect 1400 33594 1452 33600
rect 1504 33590 1532 34002
rect 1492 33584 1544 33590
rect 1492 33526 1544 33532
rect 1596 32434 1624 34031
rect 2056 32473 2084 34478
rect 2240 33289 2268 35430
rect 2504 35148 2556 35154
rect 2504 35090 2556 35096
rect 2516 34542 2544 35090
rect 2596 34672 2648 34678
rect 2596 34614 2648 34620
rect 2504 34536 2556 34542
rect 2504 34478 2556 34484
rect 2410 33552 2466 33561
rect 2410 33487 2412 33496
rect 2464 33487 2466 33496
rect 2412 33458 2464 33464
rect 2226 33280 2282 33289
rect 2226 33215 2282 33224
rect 2042 32464 2098 32473
rect 1584 32428 1636 32434
rect 2042 32399 2098 32408
rect 1584 32370 1636 32376
rect 2228 32224 2280 32230
rect 2228 32166 2280 32172
rect 2240 31929 2268 32166
rect 2226 31920 2282 31929
rect 2226 31855 2282 31864
rect 2412 31680 2464 31686
rect 1582 31648 1638 31657
rect 2412 31622 2464 31628
rect 1582 31583 1638 31592
rect 1596 31346 1624 31583
rect 1584 31340 1636 31346
rect 1584 31282 1636 31288
rect 2424 31278 2452 31622
rect 1676 31272 1728 31278
rect 1676 31214 1728 31220
rect 2412 31272 2464 31278
rect 2412 31214 2464 31220
rect 1688 30938 1716 31214
rect 1676 30932 1728 30938
rect 1676 30874 1728 30880
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 940 30660 992 30666
rect 940 30602 992 30608
rect 2056 30190 2084 30738
rect 2044 30184 2096 30190
rect 2042 30152 2044 30161
rect 2096 30152 2098 30161
rect 2042 30087 2098 30096
rect 1674 29336 1730 29345
rect 1674 29271 1730 29280
rect 1688 27606 1716 29271
rect 1676 27600 1728 27606
rect 1676 27542 1728 27548
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 1582 27024 1638 27033
rect 1582 26959 1638 26968
rect 1596 24818 1624 26959
rect 1688 26790 1716 27406
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26586 1716 26726
rect 1676 26580 1728 26586
rect 1676 26522 1728 26528
rect 2136 25696 2188 25702
rect 2136 25638 2188 25644
rect 2148 25498 2176 25638
rect 2136 25492 2188 25498
rect 2136 25434 2188 25440
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2226 22672 2282 22681
rect 2226 22607 2228 22616
rect 2280 22607 2282 22616
rect 2228 22578 2280 22584
rect 1676 22500 1728 22506
rect 1676 22442 1728 22448
rect 1688 22273 1716 22442
rect 1674 22264 1730 22273
rect 2424 22234 2452 24550
rect 2516 24177 2544 34478
rect 2608 30054 2636 34614
rect 2964 34060 3016 34066
rect 2964 34002 3016 34008
rect 2976 33318 3004 34002
rect 3056 33380 3108 33386
rect 3056 33322 3108 33328
rect 2964 33312 3016 33318
rect 2964 33254 3016 33260
rect 2780 32020 2832 32026
rect 2780 31962 2832 31968
rect 2688 31748 2740 31754
rect 2688 31690 2740 31696
rect 2700 31482 2728 31690
rect 2688 31476 2740 31482
rect 2688 31418 2740 31424
rect 2688 30932 2740 30938
rect 2792 30920 2820 31962
rect 2872 31884 2924 31890
rect 2872 31826 2924 31832
rect 2884 30938 2912 31826
rect 2740 30892 2820 30920
rect 2872 30932 2924 30938
rect 2688 30874 2740 30880
rect 2872 30874 2924 30880
rect 2596 30048 2648 30054
rect 2596 29990 2648 29996
rect 2976 28762 3004 33254
rect 3068 32774 3096 33322
rect 3056 32768 3108 32774
rect 3056 32710 3108 32716
rect 3068 31346 3096 32710
rect 3056 31340 3108 31346
rect 3056 31282 3108 31288
rect 3252 29306 3280 35566
rect 4172 35290 4200 39520
rect 4540 36378 4568 39520
rect 4528 36372 4580 36378
rect 4528 36314 4580 36320
rect 4252 36236 4304 36242
rect 4252 36178 4304 36184
rect 4264 35494 4292 36178
rect 4252 35488 4304 35494
rect 4252 35430 4304 35436
rect 4160 35284 4212 35290
rect 4160 35226 4212 35232
rect 4068 35148 4120 35154
rect 4068 35090 4120 35096
rect 3516 34944 3568 34950
rect 3516 34886 3568 34892
rect 3528 34542 3556 34886
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 4080 34785 4108 35090
rect 4066 34776 4122 34785
rect 4066 34711 4068 34720
rect 4120 34711 4122 34720
rect 4068 34682 4120 34688
rect 4080 34651 4108 34682
rect 3516 34536 3568 34542
rect 3516 34478 3568 34484
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 3700 34468 3752 34474
rect 3700 34410 3752 34416
rect 3712 33930 3740 34410
rect 4080 34066 4108 34478
rect 4068 34060 4120 34066
rect 4068 34002 4120 34008
rect 3700 33924 3752 33930
rect 3700 33866 3752 33872
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 4080 33454 4108 34002
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4080 33114 4108 33390
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3424 32768 3476 32774
rect 3424 32710 3476 32716
rect 3436 32434 3464 32710
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3424 32428 3476 32434
rect 3424 32370 3476 32376
rect 3332 32224 3384 32230
rect 3332 32166 3384 32172
rect 3344 32026 3372 32166
rect 3332 32020 3384 32026
rect 3332 31962 3384 31968
rect 3436 31482 3464 32370
rect 4160 32292 4212 32298
rect 4160 32234 4212 32240
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 4172 31482 4200 32234
rect 3424 31476 3476 31482
rect 3424 31418 3476 31424
rect 4160 31476 4212 31482
rect 4160 31418 4212 31424
rect 3976 31204 4028 31210
rect 3976 31146 4028 31152
rect 3792 31136 3844 31142
rect 3792 31078 3844 31084
rect 3804 30938 3832 31078
rect 3988 30938 4016 31146
rect 3516 30932 3568 30938
rect 3516 30874 3568 30880
rect 3792 30932 3844 30938
rect 3792 30874 3844 30880
rect 3976 30932 4028 30938
rect 3976 30874 4028 30880
rect 3528 30394 3556 30874
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3516 30388 3568 30394
rect 3516 30330 3568 30336
rect 4160 30048 4212 30054
rect 4160 29990 4212 29996
rect 4172 29782 4200 29990
rect 4160 29776 4212 29782
rect 4160 29718 4212 29724
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3240 29300 3292 29306
rect 3240 29242 3292 29248
rect 3332 28960 3384 28966
rect 3332 28902 3384 28908
rect 2964 28756 3016 28762
rect 2964 28698 3016 28704
rect 2964 26784 3016 26790
rect 2964 26726 3016 26732
rect 2780 26512 2832 26518
rect 2780 26454 2832 26460
rect 2792 26058 2820 26454
rect 2872 26444 2924 26450
rect 2872 26386 2924 26392
rect 2608 26042 2820 26058
rect 2596 26036 2820 26042
rect 2648 26030 2820 26036
rect 2596 25978 2648 25984
rect 2780 25764 2832 25770
rect 2780 25706 2832 25712
rect 2792 25430 2820 25706
rect 2884 25498 2912 26386
rect 2976 26382 3004 26726
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 2976 25702 3004 26318
rect 2964 25696 3016 25702
rect 2964 25638 3016 25644
rect 2872 25492 2924 25498
rect 2872 25434 2924 25440
rect 2780 25424 2832 25430
rect 2780 25366 2832 25372
rect 2778 24576 2834 24585
rect 2778 24511 2834 24520
rect 2502 24168 2558 24177
rect 2502 24103 2558 24112
rect 1674 22199 1730 22208
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2412 21956 2464 21962
rect 2412 21898 2464 21904
rect 1400 21888 1452 21894
rect 1400 21830 1452 21836
rect 1412 19922 1440 21830
rect 2424 21690 2452 21898
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2516 21554 2544 22034
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21146 1716 21286
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 2240 20534 2268 21354
rect 2228 20528 2280 20534
rect 2228 20470 2280 20476
rect 2516 20466 2544 21490
rect 2700 20806 2728 22034
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2516 20058 2544 20402
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 1582 19952 1638 19961
rect 1400 19916 1452 19922
rect 1582 19887 1638 19896
rect 1400 19858 1452 19864
rect 1412 19514 1440 19858
rect 1596 19854 1624 19887
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 2792 19802 2820 24511
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 2884 21146 2912 21966
rect 3252 21690 3280 21966
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3148 21412 3200 21418
rect 3148 21354 3200 21360
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 2976 20602 3004 21014
rect 3056 21004 3108 21010
rect 3056 20946 3108 20952
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2884 19990 2912 20266
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2792 19774 2912 19802
rect 2688 19712 2740 19718
rect 2740 19689 2820 19700
rect 2740 19680 2834 19689
rect 2740 19672 2778 19680
rect 2688 19654 2740 19660
rect 2778 19615 2834 19624
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 2792 18426 2820 19615
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 1674 17640 1730 17649
rect 1674 17575 1730 17584
rect 1688 16726 1716 17575
rect 2884 16726 2912 19774
rect 2976 19514 3004 20538
rect 3068 19689 3096 20946
rect 3160 20874 3188 21354
rect 3148 20868 3200 20874
rect 3148 20810 3200 20816
rect 3054 19680 3110 19689
rect 3054 19615 3110 19624
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 3344 19310 3372 28902
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3424 26920 3476 26926
rect 3424 26862 3476 26868
rect 3436 26586 3464 26862
rect 3424 26580 3476 26586
rect 3424 26522 3476 26528
rect 3436 25838 3464 26522
rect 3976 26512 4028 26518
rect 3976 26454 4028 26460
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3988 26042 4016 26454
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3424 25832 3476 25838
rect 3424 25774 3476 25780
rect 3436 25362 3464 25774
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3988 23866 4016 24210
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 3436 22098 3464 22374
rect 3712 22166 3740 22510
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3516 19984 3568 19990
rect 3516 19926 3568 19932
rect 3528 19378 3556 19926
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 1412 16697 1440 16723
rect 1676 16720 1728 16726
rect 1398 16688 1454 16697
rect 1676 16662 1728 16668
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 1398 16623 1400 16632
rect 1452 16623 1454 16632
rect 1400 16594 1452 16600
rect 1412 16250 1440 16594
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2792 16250 2820 16458
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 1688 14550 1716 15127
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 14006 1716 14350
rect 1676 14000 1728 14006
rect 1674 13968 1676 13977
rect 1728 13968 1730 13977
rect 1674 13903 1730 13912
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1596 11762 1624 12815
rect 3068 12220 3096 19246
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18630 3372 19110
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3160 17882 3188 18226
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3252 16998 3280 17614
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16046 3280 16934
rect 3344 16561 3372 18566
rect 3528 18290 3556 19314
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3700 18216 3752 18222
rect 3698 18184 3700 18193
rect 3752 18184 3754 18193
rect 3698 18119 3754 18128
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3528 17338 3556 18022
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3974 17232 4030 17241
rect 3974 17167 3976 17176
rect 4028 17167 4030 17176
rect 3976 17138 4028 17144
rect 3974 17096 4030 17105
rect 3974 17031 3976 17040
rect 4028 17031 4030 17040
rect 3976 17002 4028 17008
rect 3988 16794 4016 17002
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3330 16552 3386 16561
rect 3330 16487 3386 16496
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3792 15904 3844 15910
rect 3790 15872 3792 15881
rect 3844 15872 3846 15881
rect 3790 15807 3846 15816
rect 3988 15502 4016 15982
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3792 14816 3844 14822
rect 3790 14784 3792 14793
rect 3988 14804 4016 15438
rect 3844 14784 4016 14804
rect 3846 14776 4016 14784
rect 3790 14719 3846 14728
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 4080 13190 4108 28698
rect 4264 24682 4292 35430
rect 4620 34400 4672 34406
rect 4620 34342 4672 34348
rect 4632 34134 4660 34342
rect 4620 34128 4672 34134
rect 4620 34070 4672 34076
rect 4344 33856 4396 33862
rect 4344 33798 4396 33804
rect 4356 33318 4384 33798
rect 4632 33318 4660 34070
rect 4804 33448 4856 33454
rect 4804 33390 4856 33396
rect 4344 33312 4396 33318
rect 4344 33254 4396 33260
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4356 32502 4384 33254
rect 4436 32972 4488 32978
rect 4436 32914 4488 32920
rect 4344 32496 4396 32502
rect 4344 32438 4396 32444
rect 4448 32230 4476 32914
rect 4528 32768 4580 32774
rect 4528 32710 4580 32716
rect 4540 32366 4568 32710
rect 4528 32360 4580 32366
rect 4528 32302 4580 32308
rect 4436 32224 4488 32230
rect 4436 32166 4488 32172
rect 4448 31142 4476 32166
rect 4632 31754 4660 33254
rect 4620 31748 4672 31754
rect 4620 31690 4672 31696
rect 4528 31680 4580 31686
rect 4816 31668 4844 33390
rect 5000 33114 5028 39520
rect 5368 37210 5396 39520
rect 5368 37182 5580 37210
rect 5552 36378 5580 37182
rect 5540 36372 5592 36378
rect 5540 36314 5592 36320
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 5460 35494 5488 36178
rect 5540 35556 5592 35562
rect 5540 35498 5592 35504
rect 5448 35488 5500 35494
rect 5448 35430 5500 35436
rect 4988 33108 5040 33114
rect 4988 33050 5040 33056
rect 5264 32768 5316 32774
rect 5264 32710 5316 32716
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5276 32502 5304 32710
rect 5264 32496 5316 32502
rect 5264 32438 5316 32444
rect 5368 32434 5396 32710
rect 5356 32428 5408 32434
rect 5356 32370 5408 32376
rect 4896 32224 4948 32230
rect 4896 32166 4948 32172
rect 4908 31890 4936 32166
rect 5368 32026 5396 32370
rect 5356 32020 5408 32026
rect 5356 31962 5408 31968
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 4816 31640 4936 31668
rect 4528 31622 4580 31628
rect 4540 31210 4568 31622
rect 4528 31204 4580 31210
rect 4528 31146 4580 31152
rect 4436 31136 4488 31142
rect 4436 31078 4488 31084
rect 4436 30796 4488 30802
rect 4436 30738 4488 30744
rect 4448 30297 4476 30738
rect 4434 30288 4490 30297
rect 4434 30223 4490 30232
rect 4448 29850 4476 30223
rect 4436 29844 4488 29850
rect 4436 29786 4488 29792
rect 4540 29306 4568 31146
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4816 30258 4844 30670
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4816 29714 4844 30194
rect 4804 29708 4856 29714
rect 4804 29650 4856 29656
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4816 29170 4844 29650
rect 4804 29164 4856 29170
rect 4804 29106 4856 29112
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4252 24676 4304 24682
rect 4252 24618 4304 24624
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4264 23866 4292 24142
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4172 22574 4200 23054
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4252 19848 4304 19854
rect 4356 19836 4384 28358
rect 4816 27130 4844 29106
rect 4804 27124 4856 27130
rect 4804 27066 4856 27072
rect 4436 25356 4488 25362
rect 4436 25298 4488 25304
rect 4448 24954 4476 25298
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4448 24410 4476 24890
rect 4540 24750 4568 25230
rect 4632 24886 4660 25230
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4528 24744 4580 24750
rect 4528 24686 4580 24692
rect 4540 24410 4568 24686
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4528 24404 4580 24410
rect 4528 24346 4580 24352
rect 4802 24168 4858 24177
rect 4802 24103 4858 24112
rect 4816 23866 4844 24103
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4816 23730 4844 23802
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 4528 21004 4580 21010
rect 4528 20946 4580 20952
rect 4540 20602 4568 20946
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4540 20058 4568 20538
rect 4632 20534 4660 20878
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4304 19808 4384 19836
rect 4252 19790 4304 19796
rect 4264 19174 4292 19790
rect 4724 19174 4752 21014
rect 4908 20856 4936 31640
rect 5354 31376 5410 31385
rect 5354 31311 5410 31320
rect 5080 31136 5132 31142
rect 5080 31078 5132 31084
rect 4988 30796 5040 30802
rect 4988 30738 5040 30744
rect 5000 30190 5028 30738
rect 4988 30184 5040 30190
rect 4986 30152 4988 30161
rect 5040 30152 5042 30161
rect 4986 30087 5042 30096
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 5000 29510 5028 29990
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 5000 28422 5028 29446
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 5000 26518 5028 28358
rect 4988 26512 5040 26518
rect 4988 26454 5040 26460
rect 5092 24313 5120 31078
rect 5368 30938 5396 31311
rect 5356 30932 5408 30938
rect 5356 30874 5408 30880
rect 5264 30116 5316 30122
rect 5264 30058 5316 30064
rect 5170 29744 5226 29753
rect 5170 29679 5226 29688
rect 5184 29102 5212 29679
rect 5276 29209 5304 30058
rect 5262 29200 5318 29209
rect 5262 29135 5318 29144
rect 5172 29096 5224 29102
rect 5172 29038 5224 29044
rect 5184 28490 5212 29038
rect 5172 28484 5224 28490
rect 5172 28426 5224 28432
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 5368 27674 5396 27814
rect 5356 27668 5408 27674
rect 5356 27610 5408 27616
rect 5172 27328 5224 27334
rect 5172 27270 5224 27276
rect 5184 26450 5212 27270
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 5184 26330 5212 26386
rect 5184 26302 5304 26330
rect 5172 25968 5224 25974
rect 5172 25910 5224 25916
rect 5184 25498 5212 25910
rect 5276 25702 5304 26302
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5172 25492 5224 25498
rect 5172 25434 5224 25440
rect 5184 25294 5212 25434
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5276 24818 5304 25638
rect 5264 24812 5316 24818
rect 5460 24800 5488 35430
rect 5552 32434 5580 35498
rect 5736 33658 5764 39520
rect 6196 35834 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6184 35828 6236 35834
rect 6184 35770 6236 35776
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 5828 33862 5856 34002
rect 5816 33856 5868 33862
rect 5816 33798 5868 33804
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 5828 33318 5856 33798
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 5540 31748 5592 31754
rect 5540 31690 5592 31696
rect 5552 31346 5580 31690
rect 5632 31408 5684 31414
rect 5736 31385 5764 31758
rect 5632 31350 5684 31356
rect 5722 31376 5778 31385
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 5552 29850 5580 31282
rect 5644 30938 5672 31350
rect 5722 31311 5778 31320
rect 5632 30932 5684 30938
rect 5632 30874 5684 30880
rect 5828 30258 5856 33254
rect 6012 30705 6040 35430
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6656 35290 6684 37726
rect 6932 35834 6960 39520
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 6644 35284 6696 35290
rect 6644 35226 6696 35232
rect 6184 35148 6236 35154
rect 6184 35090 6236 35096
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 6196 34542 6224 35090
rect 6184 34536 6236 34542
rect 6184 34478 6236 34484
rect 6092 33312 6144 33318
rect 6090 33280 6092 33289
rect 6144 33280 6146 33289
rect 6090 33215 6146 33224
rect 6196 31890 6224 34478
rect 6932 34406 6960 35090
rect 7392 34746 7420 39520
rect 7472 35488 7524 35494
rect 7470 35456 7472 35465
rect 7524 35456 7526 35465
rect 7470 35391 7526 35400
rect 7760 35290 7788 39520
rect 8024 35760 8076 35766
rect 8022 35728 8024 35737
rect 8076 35728 8078 35737
rect 8022 35663 8078 35672
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 7932 35012 7984 35018
rect 7932 34954 7984 34960
rect 7562 34776 7618 34785
rect 7380 34740 7432 34746
rect 7562 34711 7618 34720
rect 7380 34682 7432 34688
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6736 34128 6788 34134
rect 6736 34070 6788 34076
rect 6748 33522 6776 34070
rect 7286 33552 7342 33561
rect 6736 33516 6788 33522
rect 7286 33487 7342 33496
rect 6736 33458 6788 33464
rect 6644 33312 6696 33318
rect 6644 33254 6696 33260
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6656 32910 6684 33254
rect 6748 33114 6776 33458
rect 7300 33114 7328 33487
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 6644 32904 6696 32910
rect 6644 32846 6696 32852
rect 6276 32836 6328 32842
rect 6276 32778 6328 32784
rect 6288 32570 6316 32778
rect 6276 32564 6328 32570
rect 6276 32506 6328 32512
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6656 32026 6684 32846
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6828 32360 6880 32366
rect 6828 32302 6880 32308
rect 6840 32026 6868 32302
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 6736 31952 6788 31958
rect 6736 31894 6788 31900
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 6552 31884 6604 31890
rect 6552 31826 6604 31832
rect 6092 31476 6144 31482
rect 6092 31418 6144 31424
rect 5998 30696 6054 30705
rect 5998 30631 6054 30640
rect 5816 30252 5868 30258
rect 5816 30194 5868 30200
rect 5724 30048 5776 30054
rect 5724 29990 5776 29996
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 5736 27402 5764 29990
rect 6012 27538 6040 30631
rect 6104 29102 6132 31418
rect 6196 31142 6224 31826
rect 6564 31414 6592 31826
rect 6748 31482 6776 31894
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6552 31408 6604 31414
rect 6552 31350 6604 31356
rect 6840 31278 6868 31758
rect 6828 31272 6880 31278
rect 6748 31232 6828 31260
rect 6184 31136 6236 31142
rect 6184 31078 6236 31084
rect 6196 30394 6224 31078
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6748 30870 6776 31232
rect 6828 31214 6880 31220
rect 6828 31136 6880 31142
rect 6828 31078 6880 31084
rect 6840 30977 6868 31078
rect 6826 30968 6882 30977
rect 6932 30938 6960 32710
rect 7300 32570 7328 33050
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7300 31822 7328 32166
rect 7288 31816 7340 31822
rect 7288 31758 7340 31764
rect 7380 31680 7432 31686
rect 7380 31622 7432 31628
rect 7104 31476 7156 31482
rect 7104 31418 7156 31424
rect 6826 30903 6882 30912
rect 6920 30932 6972 30938
rect 6920 30874 6972 30880
rect 6736 30864 6788 30870
rect 6736 30806 6788 30812
rect 6826 30832 6882 30841
rect 6826 30767 6882 30776
rect 6920 30796 6972 30802
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6564 30258 6592 30670
rect 6736 30388 6788 30394
rect 6736 30330 6788 30336
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29238 6684 29990
rect 6644 29232 6696 29238
rect 6644 29174 6696 29180
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6090 27568 6146 27577
rect 6000 27532 6052 27538
rect 6090 27503 6146 27512
rect 6000 27474 6052 27480
rect 5724 27396 5776 27402
rect 5724 27338 5776 27344
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5552 25906 5580 27270
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 5644 26042 5672 26454
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5540 25764 5592 25770
rect 5540 25706 5592 25712
rect 5552 25498 5580 25706
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5736 25362 5764 27338
rect 6012 27062 6040 27474
rect 6104 27470 6132 27503
rect 6092 27464 6144 27470
rect 6092 27406 6144 27412
rect 6104 27130 6132 27406
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6000 27056 6052 27062
rect 6000 26998 6052 27004
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 5908 26308 5960 26314
rect 5908 26250 5960 26256
rect 5920 25906 5948 26250
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 6104 24954 6132 25298
rect 6184 25220 6236 25226
rect 6184 25162 6236 25168
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 5460 24772 5672 24800
rect 5264 24754 5316 24760
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5078 24304 5134 24313
rect 5078 24239 5134 24248
rect 5080 24132 5132 24138
rect 5080 24074 5132 24080
rect 5092 22234 5120 24074
rect 5184 23866 5212 24550
rect 5276 24206 5304 24754
rect 5448 24676 5500 24682
rect 5448 24618 5500 24624
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5184 23254 5212 23462
rect 5276 23322 5304 24142
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5368 23254 5396 23734
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5368 22778 5396 23190
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5184 21350 5212 21966
rect 5460 21457 5488 24618
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 22778 5580 24210
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5446 21448 5502 21457
rect 5446 21383 5502 21392
rect 5552 21350 5580 22102
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 4908 20828 5028 20856
rect 5000 20516 5028 20828
rect 4908 20488 5028 20516
rect 4908 20058 4936 20488
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4908 19242 4936 19994
rect 5000 19310 5028 20198
rect 5080 19848 5132 19854
rect 5184 19825 5212 21286
rect 5644 21162 5672 24772
rect 6196 24206 6224 25162
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 6196 23866 6224 24142
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5736 22030 5764 22646
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5736 21690 5764 21966
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5368 21134 5672 21162
rect 5080 19790 5132 19796
rect 5170 19816 5226 19825
rect 5092 19378 5120 19790
rect 5170 19751 5226 19760
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15570 4200 15846
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4172 15162 4200 15506
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 15042 4292 19110
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4724 18426 4752 18702
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4356 17202 4384 17682
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4540 16454 4568 18022
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4540 15978 4568 16390
rect 4528 15972 4580 15978
rect 4528 15914 4580 15920
rect 4172 15014 4292 15042
rect 4540 15026 4568 15914
rect 4528 15020 4580 15026
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3068 12192 3188 12220
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 2226 11656 2282 11665
rect 2226 11591 2228 11600
rect 2280 11591 2282 11600
rect 2228 11562 2280 11568
rect 3056 10600 3108 10606
rect 1674 10568 1730 10577
rect 3056 10542 3108 10548
rect 1674 10503 1730 10512
rect 1490 8120 1546 8129
rect 1490 8055 1546 8064
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 940 6656 992 6662
rect 940 6598 992 6604
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 480 244 2790
rect 584 480 612 3606
rect 952 480 980 6598
rect 1412 5658 1440 7142
rect 1504 6322 1532 8055
rect 1688 8022 1716 10503
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2870 8392 2926 8401
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 2410 7984 2466 7993
rect 2410 7919 2412 7928
rect 2464 7919 2466 7928
rect 2412 7890 2464 7896
rect 2424 7546 2452 7890
rect 2516 7750 2544 8366
rect 2596 8356 2648 8362
rect 2870 8327 2926 8336
rect 2596 8298 2648 8304
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1596 6186 1624 6802
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1584 6180 1636 6186
rect 1584 6122 1636 6128
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 1596 5710 1624 5743
rect 1320 5630 1440 5658
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1320 3670 1348 5630
rect 1964 5370 1992 6598
rect 2056 6458 2084 7142
rect 2608 6798 2636 8298
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2424 6361 2452 6598
rect 2410 6352 2466 6361
rect 2410 6287 2466 6296
rect 2424 6254 2452 6287
rect 2412 6248 2464 6254
rect 2608 6202 2636 6734
rect 2412 6190 2464 6196
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2516 6174 2636 6202
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1308 3664 1360 3670
rect 1308 3606 1360 3612
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 1465 1440 2450
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 1504 1306 1532 4111
rect 1964 4078 1992 5306
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1688 3505 1716 3946
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1780 2514 1808 2790
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 1872 2394 1900 3402
rect 1412 1278 1532 1306
rect 1780 2366 1900 2394
rect 1412 480 1440 1278
rect 1780 480 1808 2366
rect 2148 480 2176 5510
rect 2332 4282 2360 6122
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5234 2452 6054
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2424 4826 2452 5170
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2516 4758 2544 6174
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2516 4554 2544 4694
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2332 4010 2360 4218
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2608 3466 2636 6054
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2792 5250 2820 5850
rect 2884 5778 2912 8327
rect 2976 5846 3004 10406
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3160 10130 3188 12192
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10470 3372 10950
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10266 3372 10406
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3344 9654 3372 10066
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3436 7834 3464 13126
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3988 10470 4016 10950
rect 4080 10606 4108 12038
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3988 8838 4016 10406
rect 4172 10146 4200 15014
rect 4528 14962 4580 14968
rect 4908 12345 4936 19178
rect 5000 18970 5028 19246
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 5092 18902 5120 19110
rect 5080 18896 5132 18902
rect 5078 18864 5080 18873
rect 5132 18864 5134 18873
rect 5078 18799 5134 18808
rect 5092 18773 5120 18799
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4894 12336 4950 12345
rect 4620 12300 4672 12306
rect 4894 12271 4950 12280
rect 4620 12242 4672 12248
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4264 11694 4292 12174
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4264 11354 4292 11630
rect 4356 11626 4384 12174
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4172 10118 4292 10146
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3252 7806 3464 7834
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2884 5370 2912 5714
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2700 5222 2820 5250
rect 3068 5234 3096 7482
rect 3252 6225 3280 7806
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7274 3464 7686
rect 3528 7546 3556 8230
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 7342 3556 7482
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3436 6662 3464 7210
rect 3988 6866 4016 8774
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3238 6216 3294 6225
rect 3238 6151 3294 6160
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 5228 3108 5234
rect 2700 5166 2728 5222
rect 3056 5170 3108 5176
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 3160 4690 3188 5578
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2872 4616 2924 4622
rect 2778 4584 2834 4593
rect 2872 4558 2924 4564
rect 2778 4519 2834 4528
rect 2792 3924 2820 4519
rect 2884 4282 2912 4558
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2792 3896 2912 3924
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2608 480 2636 3062
rect 2792 3058 2820 3606
rect 2884 3534 2912 3896
rect 3068 3534 3096 4082
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2884 3194 2912 3470
rect 3068 3398 3096 3470
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 3068 2650 3096 3334
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3160 2378 3188 4626
rect 3252 3126 3280 6151
rect 3436 5234 3464 6598
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 4172 6100 4200 9998
rect 4080 6072 4200 6100
rect 4080 5778 4108 6072
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5658 4108 5714
rect 4264 5658 4292 10118
rect 4356 9178 4384 11562
rect 4540 11218 4568 11630
rect 4632 11286 4660 12242
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 11898 4936 12174
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4540 10674 4568 11154
rect 4632 10810 4660 11222
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 9722 4568 10610
rect 4896 10464 4948 10470
rect 5000 10452 5028 18362
rect 5276 18290 5304 18566
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 16794 5212 18022
rect 5276 17338 5304 18226
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5092 15881 5120 16594
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 15910 5304 16526
rect 5264 15904 5316 15910
rect 5078 15872 5134 15881
rect 5264 15846 5316 15852
rect 5078 15807 5134 15816
rect 5092 15162 5120 15807
rect 5368 15178 5396 21134
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5460 20618 5488 21014
rect 5460 20602 5580 20618
rect 5460 20596 5592 20602
rect 5460 20590 5540 20596
rect 5540 20538 5592 20544
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5460 19122 5488 19382
rect 5540 19168 5592 19174
rect 5460 19116 5540 19122
rect 5460 19110 5592 19116
rect 5460 19094 5580 19110
rect 5460 17882 5488 19094
rect 5736 18970 5764 19722
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5552 18358 5580 18770
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5644 17338 5672 18090
rect 5736 17882 5764 18906
rect 6012 18426 6040 23598
rect 6196 23186 6224 23802
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 6196 22098 6224 23122
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6104 19242 6132 21286
rect 6196 21010 6224 22034
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6196 20534 6224 20946
rect 6564 20602 6592 20946
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 6196 20058 6224 20470
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6196 19378 6224 19994
rect 6550 19816 6606 19825
rect 6550 19751 6606 19760
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6564 19310 6592 19751
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6104 18086 6132 18770
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 15706 5488 16934
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5552 16250 5580 16730
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5080 15156 5132 15162
rect 5368 15150 5672 15178
rect 5080 15098 5132 15104
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5538 14784 5594 14793
rect 5276 14278 5304 14758
rect 5538 14719 5594 14728
rect 5552 14414 5580 14719
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 14074 5304 14214
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5552 13870 5580 14350
rect 5644 14006 5672 15150
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5540 13864 5592 13870
rect 5460 13812 5540 13818
rect 5460 13806 5592 13812
rect 5460 13790 5580 13806
rect 5078 12744 5134 12753
rect 5078 12679 5134 12688
rect 5092 10538 5120 12679
rect 5460 11286 5488 13790
rect 5644 12442 5672 13942
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5736 12322 5764 14758
rect 5828 14618 5856 14962
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5644 12294 5764 12322
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5460 11098 5488 11222
rect 5460 11070 5580 11098
rect 5552 10810 5580 11070
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 4948 10424 5028 10452
rect 4896 10406 4948 10412
rect 4908 9761 4936 10406
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5000 9926 5028 10066
rect 5092 10062 5120 10474
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4894 9752 4950 9761
rect 4528 9716 4580 9722
rect 4894 9687 4950 9696
rect 4528 9658 4580 9664
rect 4434 9616 4490 9625
rect 4540 9586 4568 9658
rect 4434 9551 4490 9560
rect 4528 9580 4580 9586
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4448 9042 4476 9551
rect 4528 9522 4580 9528
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4448 8634 4476 8978
rect 4540 8906 4568 9522
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4540 8090 4568 8842
rect 4724 8401 4752 9454
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4710 8392 4766 8401
rect 4710 8327 4766 8336
rect 4816 8090 4844 8910
rect 5000 8634 5028 9862
rect 5184 9382 5212 9998
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5184 9178 5212 9318
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4632 6730 4660 7142
rect 4816 7002 4844 8026
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5078 7848 5134 7857
rect 5000 7274 5028 7822
rect 5078 7783 5134 7792
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 5092 7002 5120 7783
rect 5276 7206 5304 7890
rect 5354 7304 5410 7313
rect 5354 7239 5410 7248
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5914 4384 6054
rect 4632 5914 4660 6666
rect 4908 6322 4936 6734
rect 5092 6458 5120 6938
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4080 5630 4200 5658
rect 4264 5630 4384 5658
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3777 3372 3878
rect 3330 3768 3386 3777
rect 3330 3703 3386 3712
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3436 3058 3464 5170
rect 4172 4826 4200 5630
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3528 4214 3556 4422
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 4080 4214 4108 4422
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 4068 4208 4120 4214
rect 4264 4185 4292 5510
rect 4068 4150 4120 4156
rect 4250 4176 4306 4185
rect 3528 4078 3556 4150
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3620 3738 3648 4150
rect 4250 4111 4306 4120
rect 3882 4040 3938 4049
rect 4356 4026 4384 5630
rect 4908 5370 4936 6258
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 5000 5574 5028 6122
rect 5184 5914 5212 6190
rect 5276 5914 5304 6326
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 5000 4826 5028 5510
rect 5092 5098 5120 5578
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4526 4312 4582 4321
rect 4526 4247 4582 4256
rect 3882 3975 3884 3984
rect 3936 3975 3938 3984
rect 3988 3998 4384 4026
rect 3884 3946 3936 3952
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3528 3194 3556 3538
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 3436 2310 3464 2994
rect 3988 2990 4016 3998
rect 4356 3913 4384 3998
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4080 3126 4108 3674
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4158 2952 4214 2961
rect 3988 2650 4016 2926
rect 4158 2887 4214 2896
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3330 1728 3386 1737
rect 3330 1663 3386 1672
rect 2962 1592 3018 1601
rect 2962 1527 3018 1536
rect 2976 480 3004 1527
rect 3344 480 3372 1663
rect 3790 1456 3846 1465
rect 3790 1391 3846 1400
rect 3804 480 3832 1391
rect 4172 480 4200 2887
rect 4264 2582 4292 3334
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4540 480 4568 4247
rect 4816 4049 4844 4626
rect 4908 4214 4936 4694
rect 5092 4622 5120 5034
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5092 4282 5120 4558
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4986 4176 5042 4185
rect 4986 4111 5042 4120
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4710 3496 4766 3505
rect 4632 2922 4660 3470
rect 4710 3431 4766 3440
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4724 2650 4752 3431
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5000 480 5028 4111
rect 5092 3738 5120 4218
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5092 3194 5120 3674
rect 5276 3602 5304 5850
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5092 2650 5120 2858
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5368 480 5396 7239
rect 5460 6984 5488 9590
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5552 8430 5580 9046
rect 5644 8430 5672 12294
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5736 11558 5764 12174
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11218 5764 11494
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10470 5764 11154
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10062 5764 10406
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5736 9722 5764 9998
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 8498 5764 9522
rect 5828 9382 5856 12378
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5632 8424 5684 8430
rect 5828 8378 5856 9318
rect 5632 8366 5684 8372
rect 5644 7478 5672 8366
rect 5736 8350 5856 8378
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5460 6956 5580 6984
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5460 6730 5488 6802
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6458 5488 6666
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5552 6390 5580 6956
rect 5630 6488 5686 6497
rect 5630 6423 5686 6432
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5166 5580 5714
rect 5540 5160 5592 5166
rect 5538 5128 5540 5137
rect 5592 5128 5594 5137
rect 5538 5063 5594 5072
rect 5448 4752 5500 4758
rect 5644 4740 5672 6423
rect 5736 4865 5764 8350
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 5896 5948 7210
rect 6012 6497 6040 10202
rect 6104 10033 6132 18022
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6564 14958 6592 15438
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6196 13938 6224 14418
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10742 6500 10950
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6656 10266 6684 29038
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6748 10146 6776 30330
rect 6840 29306 6868 30767
rect 6920 30738 6972 30744
rect 6932 30054 6960 30738
rect 6920 30048 6972 30054
rect 6920 29990 6972 29996
rect 7010 29880 7066 29889
rect 7010 29815 7066 29824
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 6932 29170 6960 29446
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 28014 6868 28358
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 6920 27940 6972 27946
rect 6920 27882 6972 27888
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6840 26994 6868 27338
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6932 26926 6960 27882
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6840 25838 6868 26726
rect 6932 26586 6960 26862
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6840 23866 6868 24210
rect 6932 24070 6960 24550
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6932 23594 6960 24006
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 7024 22438 7052 29815
rect 7116 28490 7144 31418
rect 7392 31346 7420 31622
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7288 31136 7340 31142
rect 7288 31078 7340 31084
rect 7300 30938 7328 31078
rect 7288 30932 7340 30938
rect 7288 30874 7340 30880
rect 7392 30802 7420 31282
rect 7380 30796 7432 30802
rect 7380 30738 7432 30744
rect 7288 30184 7340 30190
rect 7288 30126 7340 30132
rect 7300 29782 7328 30126
rect 7484 29889 7512 32506
rect 7576 32502 7604 34711
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7564 32496 7616 32502
rect 7564 32438 7616 32444
rect 7470 29880 7526 29889
rect 7470 29815 7526 29824
rect 7288 29776 7340 29782
rect 7288 29718 7340 29724
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7208 28762 7236 28970
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7104 28484 7156 28490
rect 7104 28426 7156 28432
rect 7300 27402 7328 29106
rect 7470 28656 7526 28665
rect 7470 28591 7526 28600
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 7286 26888 7342 26897
rect 7286 26823 7288 26832
rect 7340 26823 7342 26832
rect 7288 26794 7340 26800
rect 7392 26586 7420 27406
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7392 26489 7420 26522
rect 7378 26480 7434 26489
rect 7378 26415 7434 26424
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7102 24712 7158 24721
rect 7102 24647 7158 24656
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7024 22166 7052 22374
rect 7012 22160 7064 22166
rect 7012 22102 7064 22108
rect 7116 19938 7144 24647
rect 7300 24614 7328 25094
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7208 23322 7236 24550
rect 7484 24426 7512 28591
rect 7300 24398 7512 24426
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 7024 19910 7144 19938
rect 6932 19281 6960 19858
rect 6918 19272 6974 19281
rect 6840 19242 6918 19258
rect 6828 19236 6918 19242
rect 6880 19230 6918 19236
rect 6918 19207 6974 19216
rect 6828 19178 6880 19184
rect 6826 18728 6882 18737
rect 6826 18663 6882 18672
rect 6840 18358 6868 18663
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6840 18170 6868 18294
rect 6840 18142 6960 18170
rect 6932 17082 6960 18142
rect 7024 17241 7052 19910
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19310 7144 19790
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18970 7144 19246
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17542 7144 18022
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7010 17232 7066 17241
rect 7010 17167 7066 17176
rect 6932 17054 7052 17082
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 16046 6868 16594
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6840 10606 6868 11222
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6564 10118 6776 10146
rect 6090 10024 6146 10033
rect 6090 9959 6146 9968
rect 6564 9874 6592 10118
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6104 9846 6592 9874
rect 5998 6488 6054 6497
rect 5998 6423 6054 6432
rect 5998 6352 6054 6361
rect 5998 6287 6054 6296
rect 5828 5868 5948 5896
rect 5722 4856 5778 4865
rect 5722 4791 5778 4800
rect 5500 4712 5672 4740
rect 5448 4694 5500 4700
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5736 3738 5764 4626
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5828 3670 5856 5868
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 5302 5948 5714
rect 5908 5296 5960 5302
rect 5906 5264 5908 5273
rect 5960 5264 5962 5273
rect 5906 5199 5962 5208
rect 6012 4826 6040 6287
rect 6104 5846 6132 9846
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6656 9110 6684 9998
rect 6932 9602 6960 13466
rect 7024 11801 7052 17054
rect 7116 12753 7144 17478
rect 7208 13938 7236 22714
rect 7300 22574 7328 24398
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7484 22778 7512 23462
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7300 22234 7328 22510
rect 7576 22386 7604 32438
rect 7668 29753 7696 34342
rect 7840 32292 7892 32298
rect 7840 32234 7892 32240
rect 7748 31680 7800 31686
rect 7748 31622 7800 31628
rect 7760 31482 7788 31622
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 7654 29744 7710 29753
rect 7654 29679 7710 29688
rect 7654 29472 7710 29481
rect 7654 29407 7710 29416
rect 7668 27690 7696 29407
rect 7852 28665 7880 32234
rect 7944 29850 7972 34954
rect 8024 34944 8076 34950
rect 8220 34898 8248 39520
rect 8300 35488 8352 35494
rect 8300 35430 8352 35436
rect 8024 34886 8076 34892
rect 8036 34610 8064 34886
rect 8128 34870 8248 34898
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 8024 33856 8076 33862
rect 8024 33798 8076 33804
rect 8036 32910 8064 33798
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 8036 32434 8064 32846
rect 8024 32428 8076 32434
rect 8024 32370 8076 32376
rect 8036 31686 8064 32370
rect 8024 31680 8076 31686
rect 8024 31622 8076 31628
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 8036 30190 8064 30874
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 8128 29714 8156 34870
rect 8206 34776 8262 34785
rect 8206 34711 8262 34720
rect 8220 34542 8248 34711
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 8208 33380 8260 33386
rect 8208 33322 8260 33328
rect 8220 31890 8248 33322
rect 8208 31884 8260 31890
rect 8208 31826 8260 31832
rect 8208 31748 8260 31754
rect 8208 31690 8260 31696
rect 8220 31482 8248 31690
rect 8208 31476 8260 31482
rect 8208 31418 8260 31424
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 8128 29073 8156 29650
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 8114 29064 8170 29073
rect 8114 28999 8170 29008
rect 7932 28688 7984 28694
rect 7838 28656 7894 28665
rect 7932 28630 7984 28636
rect 7838 28591 7894 28600
rect 7748 28552 7800 28558
rect 7746 28520 7748 28529
rect 7840 28552 7892 28558
rect 7800 28520 7802 28529
rect 7840 28494 7892 28500
rect 7746 28455 7802 28464
rect 7760 28218 7788 28455
rect 7748 28212 7800 28218
rect 7748 28154 7800 28160
rect 7852 27946 7880 28494
rect 7840 27940 7892 27946
rect 7840 27882 7892 27888
rect 7668 27662 7788 27690
rect 7760 27606 7788 27662
rect 7748 27600 7800 27606
rect 7748 27542 7800 27548
rect 7760 26790 7788 27542
rect 7852 27470 7880 27882
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7748 26784 7800 26790
rect 7748 26726 7800 26732
rect 7656 25220 7708 25226
rect 7656 25162 7708 25168
rect 7668 24818 7696 25162
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7656 24608 7708 24614
rect 7654 24576 7656 24585
rect 7708 24576 7710 24585
rect 7654 24511 7710 24520
rect 7656 23588 7708 23594
rect 7656 23530 7708 23536
rect 7484 22358 7604 22386
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7300 20097 7328 22170
rect 7286 20088 7342 20097
rect 7286 20023 7342 20032
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7300 19825 7328 19858
rect 7286 19816 7342 19825
rect 7286 19751 7342 19760
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7300 18290 7328 18702
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7300 17882 7328 18226
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7300 15706 7328 17818
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16697 7420 16934
rect 7378 16688 7434 16697
rect 7378 16623 7434 16632
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7300 15026 7328 15642
rect 7392 15570 7420 15914
rect 7484 15638 7512 22358
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7576 20233 7604 22102
rect 7668 21690 7696 23530
rect 7760 22545 7788 26726
rect 7852 26586 7880 27406
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22681 7880 22918
rect 7838 22672 7894 22681
rect 7838 22607 7894 22616
rect 7746 22536 7802 22545
rect 7746 22471 7802 22480
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7852 21010 7880 22374
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7562 20224 7618 20233
rect 7562 20159 7618 20168
rect 7576 18737 7604 20159
rect 7852 20058 7880 20742
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7562 18728 7618 18737
rect 7944 18714 7972 28630
rect 8116 28416 8168 28422
rect 8116 28358 8168 28364
rect 8128 27674 8156 28358
rect 8220 28218 8248 29106
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 8128 27538 8156 27610
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 8220 25362 8248 26726
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 8312 24857 8340 35430
rect 8392 35148 8444 35154
rect 8392 35090 8444 35096
rect 8404 32570 8432 35090
rect 8484 34672 8536 34678
rect 8482 34640 8484 34649
rect 8536 34640 8538 34649
rect 8482 34575 8538 34584
rect 8588 33590 8616 39520
rect 8956 37210 8984 39520
rect 8772 37182 8984 37210
rect 8668 35080 8720 35086
rect 8668 35022 8720 35028
rect 8680 34134 8708 35022
rect 8668 34128 8720 34134
rect 8668 34070 8720 34076
rect 8680 33658 8708 34070
rect 8772 33810 8800 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9218 35592 9274 35601
rect 9218 35527 9274 35536
rect 9232 35494 9260 35527
rect 9220 35488 9272 35494
rect 9220 35430 9272 35436
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 8864 34678 8892 34886
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8852 34672 8904 34678
rect 8852 34614 8904 34620
rect 8864 34542 8892 34614
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 9128 34604 9180 34610
rect 9128 34546 9180 34552
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8956 34202 8984 34546
rect 8944 34196 8996 34202
rect 8944 34138 8996 34144
rect 9140 34134 9168 34546
rect 9128 34128 9180 34134
rect 9128 34070 9180 34076
rect 9312 33992 9364 33998
rect 9312 33934 9364 33940
rect 8772 33782 8892 33810
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8576 33584 8628 33590
rect 8576 33526 8628 33532
rect 8392 32564 8444 32570
rect 8392 32506 8444 32512
rect 8482 32328 8538 32337
rect 8482 32263 8538 32272
rect 8496 31958 8524 32263
rect 8588 32026 8616 33526
rect 8864 32230 8892 33782
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9324 33386 9352 33934
rect 9312 33380 9364 33386
rect 9312 33322 9364 33328
rect 9324 32774 9352 33322
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8852 32224 8904 32230
rect 8852 32166 8904 32172
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8484 31952 8536 31958
rect 8390 31920 8446 31929
rect 8484 31894 8536 31900
rect 8390 31855 8446 31864
rect 8404 31482 8432 31855
rect 8680 31793 8708 32166
rect 8864 31958 8892 32166
rect 8852 31952 8904 31958
rect 8852 31894 8904 31900
rect 8666 31784 8722 31793
rect 8666 31719 8722 31728
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8392 31476 8444 31482
rect 8392 31418 8444 31424
rect 8496 31346 8524 31622
rect 8484 31340 8536 31346
rect 8484 31282 8536 31288
rect 8392 30932 8444 30938
rect 8496 30920 8524 31282
rect 8576 31204 8628 31210
rect 8576 31146 8628 31152
rect 8588 30977 8616 31146
rect 8760 31136 8812 31142
rect 8760 31078 8812 31084
rect 8444 30892 8524 30920
rect 8574 30968 8630 30977
rect 8574 30903 8576 30912
rect 8392 30874 8444 30880
rect 8628 30903 8630 30912
rect 8576 30874 8628 30880
rect 8772 30841 8800 31078
rect 8758 30832 8814 30841
rect 8758 30767 8814 30776
rect 8864 30297 8892 31894
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8850 30288 8906 30297
rect 8850 30223 8906 30232
rect 8390 30152 8446 30161
rect 8390 30087 8446 30096
rect 8404 29714 8432 30087
rect 8668 30048 8720 30054
rect 8668 29990 8720 29996
rect 8392 29708 8444 29714
rect 8392 29650 8444 29656
rect 8404 29034 8432 29650
rect 8484 29640 8536 29646
rect 8576 29640 8628 29646
rect 8484 29582 8536 29588
rect 8574 29608 8576 29617
rect 8628 29608 8630 29617
rect 8496 29306 8524 29582
rect 8574 29543 8630 29552
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 8482 29200 8538 29209
rect 8482 29135 8484 29144
rect 8536 29135 8538 29144
rect 8484 29106 8536 29112
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 8404 26790 8432 28970
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8392 26240 8444 26246
rect 8390 26208 8392 26217
rect 8444 26208 8446 26217
rect 8390 26143 8446 26152
rect 8496 25786 8524 29106
rect 8588 28762 8616 29543
rect 8680 29170 8708 29990
rect 8668 29164 8720 29170
rect 8668 29106 8720 29112
rect 8666 29064 8722 29073
rect 8666 28999 8722 29008
rect 8680 28966 8708 28999
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8576 28756 8628 28762
rect 8576 28698 8628 28704
rect 8576 28416 8628 28422
rect 8680 28404 8708 28902
rect 8760 28620 8812 28626
rect 8760 28562 8812 28568
rect 8628 28376 8708 28404
rect 8576 28358 8628 28364
rect 8404 25758 8524 25786
rect 8298 24848 8354 24857
rect 8404 24818 8432 25758
rect 8484 25696 8536 25702
rect 8484 25638 8536 25644
rect 8496 25498 8524 25638
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8496 24954 8524 25434
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8482 24848 8538 24857
rect 8298 24783 8354 24792
rect 8392 24812 8444 24818
rect 8482 24783 8538 24792
rect 8392 24754 8444 24760
rect 8404 24721 8432 24754
rect 8390 24712 8446 24721
rect 8390 24647 8446 24656
rect 8496 24392 8524 24783
rect 8588 24614 8616 28358
rect 8772 28218 8800 28562
rect 8760 28212 8812 28218
rect 8760 28154 8812 28160
rect 8864 27690 8892 30223
rect 9324 30190 9352 32710
rect 9416 32298 9444 39520
rect 9784 33833 9812 39520
rect 10152 35714 10180 39520
rect 9876 35686 10180 35714
rect 9770 33824 9826 33833
rect 9770 33759 9826 33768
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 9496 32972 9548 32978
rect 9496 32914 9548 32920
rect 9508 32434 9536 32914
rect 9496 32428 9548 32434
rect 9548 32388 9628 32416
rect 9496 32370 9548 32376
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 9128 29164 9180 29170
rect 9128 29106 9180 29112
rect 9140 28762 9168 29106
rect 9416 29034 9444 31962
rect 9496 31884 9548 31890
rect 9496 31826 9548 31832
rect 9508 31482 9536 31826
rect 9496 31476 9548 31482
rect 9496 31418 9548 31424
rect 9494 31376 9550 31385
rect 9494 31311 9550 31320
rect 9404 29028 9456 29034
rect 9404 28970 9456 28976
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8680 27662 8892 27690
rect 8680 26926 8708 27662
rect 8852 27600 8904 27606
rect 8852 27542 8904 27548
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8772 26994 8800 27270
rect 8760 26988 8812 26994
rect 8760 26930 8812 26936
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8668 26784 8720 26790
rect 8668 26726 8720 26732
rect 8680 25430 8708 26726
rect 8772 26042 8800 26930
rect 8760 26036 8812 26042
rect 8760 25978 8812 25984
rect 8772 25770 8800 25978
rect 8864 25838 8892 27542
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9508 27010 9536 31311
rect 9600 29617 9628 32388
rect 9784 30433 9812 33594
rect 9876 31686 9904 35686
rect 10324 35624 10376 35630
rect 10324 35566 10376 35572
rect 10140 35284 10192 35290
rect 10140 35226 10192 35232
rect 10152 34542 10180 35226
rect 10230 34640 10286 34649
rect 10230 34575 10286 34584
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 9956 34468 10008 34474
rect 9956 34410 10008 34416
rect 9968 33658 9996 34410
rect 10152 34218 10180 34478
rect 10060 34190 10180 34218
rect 9956 33652 10008 33658
rect 9956 33594 10008 33600
rect 10060 33130 10088 34190
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 9968 33102 10088 33130
rect 9968 31770 9996 33102
rect 10152 32978 10180 34070
rect 10244 32978 10272 34575
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10244 32502 10272 32914
rect 10232 32496 10284 32502
rect 10232 32438 10284 32444
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 9948 31742 9996 31770
rect 9864 31680 9916 31686
rect 9948 31668 9976 31742
rect 10048 31680 10100 31686
rect 9948 31640 9996 31668
rect 9864 31622 9916 31628
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9770 30424 9826 30433
rect 9770 30359 9826 30368
rect 9680 30320 9732 30326
rect 9784 30308 9812 30359
rect 9732 30280 9812 30308
rect 9680 30262 9732 30268
rect 9680 30184 9732 30190
rect 9678 30152 9680 30161
rect 9732 30152 9734 30161
rect 9678 30087 9734 30096
rect 9772 29776 9824 29782
rect 9772 29718 9824 29724
rect 9586 29608 9642 29617
rect 9586 29543 9642 29552
rect 9678 29472 9734 29481
rect 9678 29407 9734 29416
rect 9692 27690 9720 29407
rect 9784 29306 9812 29718
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9876 29170 9904 31418
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9862 29064 9918 29073
rect 9862 28999 9918 29008
rect 9692 27662 9812 27690
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9692 27130 9720 27474
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9508 26982 9720 27010
rect 9036 26920 9088 26926
rect 9036 26862 9088 26868
rect 9048 26790 9076 26862
rect 9036 26784 9088 26790
rect 9036 26726 9088 26732
rect 9048 26314 9076 26726
rect 9036 26308 9088 26314
rect 9036 26250 9088 26256
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9324 26042 9352 26182
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 8852 25832 8904 25838
rect 8852 25774 8904 25780
rect 8760 25764 8812 25770
rect 8760 25706 8812 25712
rect 8864 25498 8892 25774
rect 9404 25764 9456 25770
rect 9404 25706 9456 25712
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8668 25424 8720 25430
rect 8668 25366 8720 25372
rect 8760 25356 8812 25362
rect 8760 25298 8812 25304
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8496 24364 8616 24392
rect 8024 23792 8076 23798
rect 8024 23734 8076 23740
rect 8036 22234 8064 23734
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8128 23118 8156 23462
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8128 22438 8156 23054
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 8036 21622 8064 22170
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 21690 8156 21966
rect 8220 21962 8248 23122
rect 8312 22778 8340 23258
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 8404 21554 8432 23666
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8496 21690 8524 22034
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8022 20088 8078 20097
rect 8022 20023 8078 20032
rect 7562 18663 7618 18672
rect 7852 18686 7972 18714
rect 7852 18630 7880 18686
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 17134 7788 17478
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 16794 7604 17002
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7760 16726 7788 17070
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7484 15162 7512 15574
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14482 7328 14962
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7196 13932 7248 13938
rect 7300 13920 7328 14418
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7380 13932 7432 13938
rect 7300 13892 7380 13920
rect 7196 13874 7248 13880
rect 7380 13874 7432 13880
rect 7208 13530 7236 13874
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7102 12744 7158 12753
rect 7102 12679 7158 12688
rect 7010 11792 7066 11801
rect 7010 11727 7066 11736
rect 7024 9625 7052 11727
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 6840 9574 6960 9602
rect 7010 9616 7066 9625
rect 6840 9518 6868 9574
rect 7010 9551 7066 9560
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6932 9330 6960 9386
rect 7116 9382 7144 9522
rect 7392 9518 7420 10134
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 6840 9302 6960 9330
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6196 8090 6224 8434
rect 6644 8424 6696 8430
rect 6748 8401 6776 8910
rect 6644 8366 6696 8372
rect 6734 8392 6790 8401
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6656 6882 6684 8366
rect 6734 8327 6790 8336
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 7041 6776 7278
rect 6734 7032 6790 7041
rect 6840 7002 6868 9302
rect 7024 8498 7052 9318
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6734 6967 6790 6976
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6196 6854 6684 6882
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6092 3936 6144 3942
rect 6090 3904 6092 3913
rect 6144 3904 6146 3913
rect 6090 3839 6146 3848
rect 6090 3768 6146 3777
rect 6196 3754 6224 6854
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6656 5914 6684 6734
rect 6748 6458 6776 6870
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6769 6868 6802
rect 6826 6760 6882 6769
rect 6826 6695 6882 6704
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6932 5914 6960 8230
rect 7116 8090 7144 9046
rect 7286 8936 7342 8945
rect 7286 8871 7342 8880
rect 7300 8430 7328 8871
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7392 7478 7420 9454
rect 7484 9382 7512 14010
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 10266 7604 10406
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7576 9586 7604 10202
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7484 8090 7512 9114
rect 7576 9110 7604 9522
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7576 8022 7604 8434
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 7024 7206 7052 7239
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7378 6896 7434 6905
rect 7378 6831 7434 6840
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6826 5808 6882 5817
rect 6826 5743 6882 5752
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6748 4826 6776 5510
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6564 3924 6592 4218
rect 6564 3896 6684 3924
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6146 3726 6224 3754
rect 6090 3703 6146 3712
rect 5816 3664 5868 3670
rect 6368 3664 6420 3670
rect 5816 3606 5868 3612
rect 6182 3632 6238 3641
rect 6368 3606 6420 3612
rect 6182 3567 6238 3576
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5460 2650 5488 3130
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5460 2446 5488 2586
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 1465 5856 2246
rect 5814 1456 5870 1465
rect 5814 1391 5870 1400
rect 5724 1284 5776 1290
rect 5724 1226 5776 1232
rect 5736 480 5764 1226
rect 6196 480 6224 3567
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 2990 6316 3470
rect 6380 3194 6408 3606
rect 6656 3233 6684 3896
rect 6748 3738 6776 4762
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6642 3224 6698 3233
rect 6368 3188 6420 3194
rect 6642 3159 6698 3168
rect 6368 3130 6420 3136
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6274 2408 6330 2417
rect 6274 2343 6276 2352
rect 6328 2343 6330 2352
rect 6276 2314 6328 2320
rect 6840 1306 6868 5743
rect 6932 4826 6960 5850
rect 7116 5778 7144 6054
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7024 4690 7052 4966
rect 7116 4758 7144 5714
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5234 7328 5646
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7102 4584 7158 4593
rect 7102 4519 7158 4528
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6932 3670 6960 4150
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6564 1278 6868 1306
rect 6564 480 6592 1278
rect 7116 610 7144 4519
rect 7300 3738 7328 5170
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7196 3188 7248 3194
rect 7300 3176 7328 3674
rect 7248 3148 7328 3176
rect 7196 3130 7248 3136
rect 7300 2990 7328 3148
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7208 2650 7236 2926
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 6920 604 6972 610
rect 6920 546 6972 552
rect 7104 604 7156 610
rect 7104 546 7156 552
rect 6932 480 6960 546
rect 7392 480 7420 6831
rect 7576 6322 7604 7958
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 6089 7512 6190
rect 7470 6080 7526 6089
rect 7470 6015 7526 6024
rect 7576 5216 7604 6258
rect 7668 5284 7696 15098
rect 7746 11656 7802 11665
rect 7746 11591 7802 11600
rect 7760 11354 7788 11591
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7852 7954 7880 18566
rect 8036 18086 8064 20023
rect 8128 19718 8156 20334
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8128 19417 8156 19654
rect 8114 19408 8170 19417
rect 8114 19343 8170 19352
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8220 18290 8248 19110
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17814 8340 18022
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8312 17338 8340 17750
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8114 17232 8170 17241
rect 8404 17202 8432 19110
rect 8496 17678 8524 20266
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8114 17167 8170 17176
rect 8392 17196 8444 17202
rect 8022 16688 8078 16697
rect 7932 16652 7984 16658
rect 8022 16623 8024 16632
rect 7932 16594 7984 16600
rect 8076 16623 8078 16632
rect 8024 16594 8076 16600
rect 7944 15910 7972 16594
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7944 15706 7972 15846
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 8128 14074 8156 17167
rect 8392 17138 8444 17144
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 15858 8340 17070
rect 8496 16794 8524 17614
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8496 16590 8524 16730
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8496 16250 8524 16526
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8220 15830 8340 15858
rect 8220 15502 8248 15830
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 14618 8248 15438
rect 8312 15162 8340 15642
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8312 13190 8340 14894
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 7944 12782 7972 13126
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7944 11898 7972 12718
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8220 12170 8248 12650
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8390 12336 8446 12345
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7944 11393 7972 11834
rect 7930 11384 7986 11393
rect 8036 11354 8064 12038
rect 7930 11319 7986 11328
rect 8024 11348 8076 11354
rect 7944 11286 7972 11319
rect 8024 11290 8076 11296
rect 7932 11280 7984 11286
rect 8312 11234 8340 12310
rect 8390 12271 8446 12280
rect 7932 11222 7984 11228
rect 8128 11206 8340 11234
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7944 10742 7972 11018
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7944 10266 7972 10678
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8128 10198 8156 11206
rect 8208 11144 8260 11150
rect 8260 11092 8340 11098
rect 8208 11086 8340 11092
rect 8220 11070 8340 11086
rect 8312 10266 8340 11070
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8312 9722 8340 10202
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8404 9602 8432 12271
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8496 11880 8524 12174
rect 8588 12050 8616 24364
rect 8680 24274 8708 25230
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8680 23730 8708 24210
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8680 21486 8708 22374
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8680 21146 8708 21422
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8666 21040 8722 21049
rect 8666 20975 8722 20984
rect 8680 16561 8708 20975
rect 8772 18057 8800 25298
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9416 24818 9444 25706
rect 9692 25242 9720 26982
rect 9784 26790 9812 27662
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9692 25214 9812 25242
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 9416 24410 9444 24754
rect 9692 24698 9720 25094
rect 9600 24670 9720 24698
rect 9784 24698 9812 25214
rect 9876 25158 9904 28999
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9862 24848 9918 24857
rect 9862 24783 9864 24792
rect 9916 24783 9918 24792
rect 9864 24754 9916 24760
rect 9784 24670 9904 24698
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9312 23520 9364 23526
rect 9312 23462 9364 23468
rect 9324 22982 9352 23462
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 8758 18048 8814 18057
rect 8758 17983 8814 17992
rect 8666 16552 8722 16561
rect 8666 16487 8722 16496
rect 8680 15706 8708 16487
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8680 14006 8708 15642
rect 8772 15366 8800 15982
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 14958 8800 15302
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8680 12374 8708 13466
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8588 12022 8708 12050
rect 8576 11892 8628 11898
rect 8496 11852 8576 11880
rect 8496 11354 8524 11852
rect 8576 11834 8628 11840
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8588 10810 8616 11222
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8404 9574 8524 9602
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7932 9376 7984 9382
rect 7984 9324 8064 9330
rect 7932 9318 8064 9324
rect 7944 9302 8064 9318
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7852 7546 7880 7890
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8036 7206 8064 9302
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8128 8498 8156 8774
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8312 8090 8340 8774
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 7954 8432 9454
rect 8496 8412 8524 9574
rect 8588 9178 8616 10066
rect 8680 9518 8708 12022
rect 8772 11558 8800 12174
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 9586 8800 11494
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8680 8838 8708 9318
rect 8758 8936 8814 8945
rect 8758 8871 8814 8880
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8496 8384 8616 8412
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8312 7290 8340 7754
rect 8220 7262 8340 7290
rect 7840 7200 7892 7206
rect 7838 7168 7840 7177
rect 8024 7200 8076 7206
rect 7892 7168 7894 7177
rect 8024 7142 8076 7148
rect 7838 7103 7894 7112
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6186 7788 6598
rect 7840 6248 7892 6254
rect 7838 6216 7840 6225
rect 7892 6216 7894 6225
rect 7748 6180 7800 6186
rect 7838 6151 7894 6160
rect 7748 6122 7800 6128
rect 7838 5672 7894 5681
rect 7838 5607 7894 5616
rect 7668 5256 7788 5284
rect 7576 5188 7696 5216
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4486 7512 4966
rect 7576 4554 7604 5034
rect 7668 4826 7696 5188
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4282 7512 4422
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7760 3505 7788 5256
rect 7746 3496 7802 3505
rect 7746 3431 7802 3440
rect 7746 3088 7802 3097
rect 7746 3023 7802 3032
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7668 1601 7696 2246
rect 7654 1592 7710 1601
rect 7654 1527 7710 1536
rect 7760 480 7788 3023
rect 7852 1290 7880 5607
rect 8036 4457 8064 7142
rect 8220 6798 8248 7262
rect 8300 7200 8352 7206
rect 8404 7177 8432 7890
rect 8496 7886 8524 8230
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8300 7142 8352 7148
rect 8390 7168 8446 7177
rect 8312 6934 8340 7142
rect 8390 7103 8446 7112
rect 8496 7002 8524 7822
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6361 8248 6734
rect 8206 6352 8262 6361
rect 8206 6287 8262 6296
rect 8404 5914 8432 6870
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 6254 8524 6734
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8404 5370 8432 5714
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8128 4622 8156 4762
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8220 4570 8248 4626
rect 8022 4448 8078 4457
rect 8022 4383 8078 4392
rect 8128 4214 8156 4558
rect 8220 4542 8340 4570
rect 8206 4448 8262 4457
rect 8206 4383 8262 4392
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8022 2544 8078 2553
rect 8022 2479 8024 2488
rect 8076 2479 8078 2488
rect 8024 2450 8076 2456
rect 7840 1284 7892 1290
rect 7840 1226 7892 1232
rect 8220 480 8248 4383
rect 8312 3466 8340 4542
rect 8404 4010 8432 4694
rect 8496 4185 8524 5510
rect 8482 4176 8538 4185
rect 8482 4111 8538 4120
rect 8484 4072 8536 4078
rect 8588 4060 8616 8384
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 6905 8708 8230
rect 8666 6896 8722 6905
rect 8666 6831 8722 6840
rect 8666 6760 8722 6769
rect 8666 6695 8722 6704
rect 8680 6458 8708 6695
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8772 6390 8800 8871
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8772 5658 8800 6326
rect 8864 5778 8892 22918
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22234 9444 22374
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 9312 21344 9364 21350
rect 9312 21286 9364 21292
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9218 19408 9274 19417
rect 9218 19343 9274 19352
rect 9232 19310 9260 19343
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 18970 9260 19246
rect 9324 19122 9352 21286
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19242 9444 20198
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9324 19094 9444 19122
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9324 17134 9352 18022
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9324 16794 9352 17070
rect 9416 16998 9444 19094
rect 9508 17105 9536 24550
rect 9600 23594 9628 24670
rect 9678 24576 9734 24585
rect 9678 24511 9734 24520
rect 9692 24410 9720 24511
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9678 24304 9734 24313
rect 9678 24239 9680 24248
rect 9732 24239 9734 24248
rect 9680 24210 9732 24216
rect 9876 23866 9904 24670
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9692 22137 9720 23598
rect 9876 23322 9904 23666
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9678 22128 9734 22137
rect 9678 22063 9734 22072
rect 9876 21894 9904 22374
rect 9864 21888 9916 21894
rect 9678 21856 9734 21865
rect 9864 21830 9916 21836
rect 9678 21791 9734 21800
rect 9692 17746 9720 21791
rect 9968 21706 9996 31640
rect 10048 31622 10100 31628
rect 10060 29481 10088 31622
rect 10046 29472 10102 29481
rect 10046 29407 10102 29416
rect 10048 29300 10100 29306
rect 10048 29242 10100 29248
rect 10060 28762 10088 29242
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 10048 26512 10100 26518
rect 10048 26454 10100 26460
rect 10060 25158 10088 26454
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10060 22642 10088 25094
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10152 22166 10180 32370
rect 10244 23662 10272 32438
rect 10336 31822 10364 35566
rect 10416 34944 10468 34950
rect 10416 34886 10468 34892
rect 10428 34542 10456 34886
rect 10416 34536 10468 34542
rect 10416 34478 10468 34484
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10520 33114 10548 34478
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 10506 32464 10562 32473
rect 10506 32399 10562 32408
rect 10520 32026 10548 32399
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10612 31822 10640 39520
rect 10980 35714 11008 39520
rect 10704 35686 11008 35714
rect 10324 31816 10376 31822
rect 10324 31758 10376 31764
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10508 31748 10560 31754
rect 10508 31690 10560 31696
rect 10416 31680 10468 31686
rect 10416 31622 10468 31628
rect 10324 31204 10376 31210
rect 10324 31146 10376 31152
rect 10336 30705 10364 31146
rect 10322 30696 10378 30705
rect 10322 30631 10378 30640
rect 10322 30424 10378 30433
rect 10322 30359 10378 30368
rect 10336 30190 10364 30359
rect 10324 30184 10376 30190
rect 10324 30126 10376 30132
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10336 29238 10364 29650
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10336 28762 10364 29038
rect 10428 28966 10456 31622
rect 10520 30025 10548 31690
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10506 30016 10562 30025
rect 10506 29951 10562 29960
rect 10506 29880 10562 29889
rect 10506 29815 10562 29824
rect 10520 29238 10548 29815
rect 10612 29306 10640 30670
rect 10600 29300 10652 29306
rect 10600 29242 10652 29248
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10612 28966 10640 29106
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10324 28756 10376 28762
rect 10324 28698 10376 28704
rect 10336 27674 10364 28698
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10520 27062 10548 28902
rect 10612 28422 10640 28902
rect 10600 28416 10652 28422
rect 10600 28358 10652 28364
rect 10508 27056 10560 27062
rect 10508 26998 10560 27004
rect 10704 26874 10732 35686
rect 10968 35148 11020 35154
rect 11020 35108 11100 35136
rect 10968 35090 11020 35096
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10796 34678 10824 35022
rect 11072 34762 11100 35108
rect 10980 34746 11100 34762
rect 10968 34740 11100 34746
rect 11020 34734 11100 34740
rect 10968 34682 11020 34688
rect 10784 34672 10836 34678
rect 10784 34614 10836 34620
rect 10796 34134 10824 34614
rect 10784 34128 10836 34134
rect 10784 34070 10836 34076
rect 11072 33522 11100 34734
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10784 33040 10836 33046
rect 10782 33008 10784 33017
rect 10836 33008 10838 33017
rect 10782 32943 10838 32952
rect 10796 32502 10824 32943
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10888 32570 10916 32846
rect 10876 32564 10928 32570
rect 10876 32506 10928 32512
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 10874 31920 10930 31929
rect 10874 31855 10876 31864
rect 10928 31855 10930 31864
rect 10876 31826 10928 31832
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 10796 31346 10824 31758
rect 11152 31748 11204 31754
rect 11152 31690 11204 31696
rect 10784 31340 10836 31346
rect 10784 31282 10836 31288
rect 10796 28490 10824 31282
rect 10968 31272 11020 31278
rect 11164 31260 11192 31690
rect 11020 31232 11192 31260
rect 10968 31214 11020 31220
rect 11060 31136 11112 31142
rect 11060 31078 11112 31084
rect 10876 30796 10928 30802
rect 10876 30738 10928 30744
rect 10888 30394 10916 30738
rect 10968 30592 11020 30598
rect 10968 30534 11020 30540
rect 10876 30388 10928 30394
rect 10876 30330 10928 30336
rect 10888 29850 10916 30330
rect 10876 29844 10928 29850
rect 10876 29786 10928 29792
rect 10876 29028 10928 29034
rect 10876 28970 10928 28976
rect 10888 28540 10916 28970
rect 10980 28762 11008 30534
rect 11072 29186 11100 31078
rect 11164 30433 11192 31232
rect 11150 30424 11206 30433
rect 11150 30359 11206 30368
rect 11150 30152 11206 30161
rect 11150 30087 11206 30096
rect 11164 29782 11192 30087
rect 11244 30048 11296 30054
rect 11244 29990 11296 29996
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 11150 29608 11206 29617
rect 11256 29578 11284 29990
rect 11150 29543 11152 29552
rect 11204 29543 11206 29552
rect 11244 29572 11296 29578
rect 11152 29514 11204 29520
rect 11244 29514 11296 29520
rect 11072 29158 11192 29186
rect 11256 29170 11284 29514
rect 10968 28756 11020 28762
rect 10968 28698 11020 28704
rect 11164 28694 11192 29158
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 10888 28512 11100 28540
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10520 26846 10732 26874
rect 10324 26240 10376 26246
rect 10324 26182 10376 26188
rect 10336 25294 10364 26182
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10416 24676 10468 24682
rect 10416 24618 10468 24624
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 10336 24274 10364 24550
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10324 24132 10376 24138
rect 10324 24074 10376 24080
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 10336 23526 10364 24074
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10244 22574 10272 22918
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10244 22234 10272 22510
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9876 21678 9996 21706
rect 10060 21690 10088 22034
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10048 21684 10100 21690
rect 9876 21350 9904 21678
rect 10048 21626 10100 21632
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9968 21078 9996 21558
rect 10046 21448 10102 21457
rect 10046 21383 10048 21392
rect 10100 21383 10102 21392
rect 10048 21354 10100 21360
rect 10152 21146 10180 21966
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17338 9720 17682
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9218 15056 9274 15065
rect 9218 14991 9274 15000
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 9048 14618 9076 14826
rect 9232 14822 9260 14991
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9140 13410 9168 13942
rect 9324 13802 9352 16186
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9324 13530 9352 13738
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9140 13382 9352 13410
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 9034 8392 9090 8401
rect 9034 8327 9090 8336
rect 9048 8294 9076 8327
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8090 9076 8230
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8942 7304 8998 7313
rect 8942 7239 8998 7248
rect 8956 6934 8984 7239
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8942 6760 8998 6769
rect 8942 6695 8944 6704
rect 8996 6695 8998 6704
rect 8944 6666 8996 6672
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6186 9352 13382
rect 9416 8634 9444 16934
rect 9508 16250 9536 17031
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9600 16046 9628 16526
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9508 14890 9536 15846
rect 9692 15706 9720 16623
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9508 13938 9536 14826
rect 9600 14618 9628 15438
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9600 14074 9628 14554
rect 9692 14346 9720 15506
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 11354 9536 12582
rect 9784 12442 9812 20946
rect 10048 20324 10100 20330
rect 10048 20266 10100 20272
rect 10060 20074 10088 20266
rect 10140 20256 10192 20262
rect 10138 20224 10140 20233
rect 10192 20224 10194 20233
rect 10138 20159 10194 20168
rect 10138 20088 10194 20097
rect 10060 20046 10138 20074
rect 10138 20023 10194 20032
rect 10152 19854 10180 20023
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 9862 18864 9918 18873
rect 9862 18799 9918 18808
rect 9876 16402 9904 18799
rect 10046 18048 10102 18057
rect 10046 17983 10102 17992
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9968 17202 9996 17614
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9968 16522 9996 17138
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9876 16374 9996 16402
rect 9862 16144 9918 16153
rect 9862 16079 9918 16088
rect 9876 16046 9904 16079
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9968 15858 9996 16374
rect 9876 15830 9996 15858
rect 9876 12442 9904 15830
rect 10060 15706 10088 17983
rect 10244 17814 10272 21966
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10336 16640 10364 23462
rect 10428 21010 10456 24618
rect 10520 21593 10548 26846
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10612 24410 10640 25298
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10612 22982 10640 24346
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 22030 10640 22918
rect 10704 22030 10732 26726
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10796 24206 10824 25638
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10796 23730 10824 24142
rect 10888 23866 10916 24210
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10784 23588 10836 23594
rect 10784 23530 10836 23536
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10612 21690 10640 21966
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10506 21584 10562 21593
rect 10506 21519 10562 21528
rect 10600 21412 10652 21418
rect 10600 21354 10652 21360
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 20262 10548 20946
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10428 18970 10456 19994
rect 10520 19990 10548 20198
rect 10508 19984 10560 19990
rect 10508 19926 10560 19932
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10612 17785 10640 21354
rect 10704 21350 10732 21830
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10704 21146 10732 21286
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10796 21026 10824 23530
rect 10980 22080 11008 28358
rect 11072 23594 11100 28512
rect 11164 28218 11192 28630
rect 11256 28626 11284 29106
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11152 28212 11204 28218
rect 11152 28154 11204 28160
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10980 22052 11100 22080
rect 10876 22024 10928 22030
rect 10928 21984 11008 22012
rect 10876 21966 10928 21972
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10704 20998 10824 21026
rect 10704 19938 10732 20998
rect 10888 20942 10916 21490
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10796 20058 10824 20878
rect 10888 20058 10916 20878
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10704 19910 10824 19938
rect 10690 19816 10746 19825
rect 10690 19751 10746 19760
rect 10704 18970 10732 19751
rect 10796 19281 10824 19910
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10888 19446 10916 19790
rect 10876 19440 10928 19446
rect 10874 19408 10876 19417
rect 10928 19408 10930 19417
rect 10874 19343 10930 19352
rect 10782 19272 10838 19281
rect 10782 19207 10838 19216
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10704 18426 10732 18906
rect 10796 18816 10824 19207
rect 10876 18828 10928 18834
rect 10796 18788 10876 18816
rect 10876 18770 10928 18776
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10598 17776 10654 17785
rect 10416 17740 10468 17746
rect 10598 17711 10654 17720
rect 10416 17682 10468 17688
rect 10428 16998 10456 17682
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10244 16612 10364 16640
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 13977 10180 14214
rect 10138 13968 10194 13977
rect 10138 13903 10194 13912
rect 10244 13852 10272 16612
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10336 15502 10364 16458
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 15162 10364 15438
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10152 13824 10272 13852
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9954 12336 10010 12345
rect 9600 12306 9812 12322
rect 9588 12300 9812 12306
rect 9640 12294 9812 12300
rect 9588 12242 9640 12248
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9586 11384 9642 11393
rect 9496 11348 9548 11354
rect 9586 11319 9642 11328
rect 9496 11290 9548 11296
rect 9600 11150 9628 11319
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9600 10810 9628 11086
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10146 9628 10406
rect 9692 10266 9720 12174
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9600 10118 9720 10146
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7886 9628 8230
rect 9588 7880 9640 7886
rect 9692 7857 9720 10118
rect 9784 9994 9812 12294
rect 9864 12300 9916 12306
rect 9954 12271 10010 12280
rect 9864 12242 9916 12248
rect 9876 10198 9904 12242
rect 9968 11830 9996 12271
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9968 11558 9996 11766
rect 10060 11626 10088 12106
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9968 11218 9996 11290
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9968 10742 9996 11154
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10060 10554 10088 11562
rect 9968 10526 10088 10554
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9588 7822 9640 7828
rect 9678 7848 9734 7857
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 7206 9444 7346
rect 9600 7342 9628 7822
rect 9678 7783 9734 7792
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 6866 9444 7142
rect 9600 7002 9628 7278
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9600 6798 9628 6938
rect 9588 6792 9640 6798
rect 9402 6760 9458 6769
rect 9588 6734 9640 6740
rect 9402 6695 9458 6704
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9324 5914 9352 6122
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8772 5630 8892 5658
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4321 8800 4966
rect 8758 4312 8814 4321
rect 8758 4247 8814 4256
rect 8536 4032 8708 4060
rect 8484 4014 8536 4020
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8496 2650 8524 3334
rect 8574 3224 8630 3233
rect 8574 3159 8576 3168
rect 8628 3159 8630 3168
rect 8576 3130 8628 3136
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8588 480 8616 2586
rect 8680 2009 8708 4032
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8666 2000 8722 2009
rect 8666 1935 8722 1944
rect 8772 1737 8800 2246
rect 8758 1728 8814 1737
rect 8758 1663 8814 1672
rect 8864 1442 8892 5630
rect 9416 5522 9444 6695
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5658 9536 6190
rect 9600 6186 9628 6734
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5817 9720 6054
rect 9678 5808 9734 5817
rect 9784 5778 9812 9590
rect 9876 8430 9904 10134
rect 9968 9602 9996 10526
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10060 9722 10088 10202
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9968 9574 10088 9602
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9876 8022 9904 8366
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9864 8016 9916 8022
rect 9968 7993 9996 8230
rect 9864 7958 9916 7964
rect 9954 7984 10010 7993
rect 9954 7919 10010 7928
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9968 6458 9996 6802
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10060 6338 10088 9574
rect 10152 9489 10180 13824
rect 10336 12850 10364 14282
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10232 12368 10284 12374
rect 10428 12322 10456 16934
rect 10520 16697 10548 17274
rect 10506 16688 10562 16697
rect 10506 16623 10562 16632
rect 10704 16250 10732 18362
rect 10888 18086 10916 18770
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10690 16144 10746 16153
rect 10690 16079 10746 16088
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10520 14346 10548 14418
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10520 12986 10548 14282
rect 10612 14074 10640 14418
rect 10704 14414 10732 16079
rect 10888 15314 10916 18022
rect 10796 15286 10916 15314
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 14074 10732 14350
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10612 13462 10640 14010
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10704 13530 10732 13874
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10796 13308 10824 15286
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10612 13280 10824 13308
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10232 12310 10284 12316
rect 10244 10266 10272 12310
rect 10336 12294 10456 12322
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10244 9654 10272 10202
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10138 9480 10194 9489
rect 10138 9415 10194 9424
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10152 7342 10180 8026
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9968 6310 10088 6338
rect 9678 5743 9734 5752
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9508 5630 9720 5658
rect 9416 5494 9536 5522
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9402 5400 9458 5409
rect 9402 5335 9404 5344
rect 9456 5335 9458 5344
rect 9404 5306 9456 5312
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9036 4072 9088 4078
rect 9034 4040 9036 4049
rect 9088 4040 9090 4049
rect 9034 3975 9090 3984
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9416 3369 9444 3402
rect 9402 3360 9458 3369
rect 8956 3292 9252 3312
rect 9402 3295 9458 3304
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 9402 2816 9458 2825
rect 9402 2751 9458 2760
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8864 1414 8984 1442
rect 8956 480 8984 1414
rect 9416 480 9444 2751
rect 9508 2582 9536 5494
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9600 4010 9628 5306
rect 9692 5250 9720 5630
rect 9784 5370 9812 5714
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9692 5222 9812 5250
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9692 3754 9720 4558
rect 9600 3738 9720 3754
rect 9588 3732 9720 3738
rect 9640 3726 9720 3732
rect 9588 3674 9640 3680
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9600 3194 9628 3538
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9692 2650 9720 3726
rect 9784 3466 9812 5222
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9770 2680 9826 2689
rect 9680 2644 9732 2650
rect 9770 2615 9826 2624
rect 9680 2586 9732 2592
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9784 2514 9812 2615
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9968 2446 9996 6310
rect 10232 6248 10284 6254
rect 10230 6216 10232 6225
rect 10284 6216 10286 6225
rect 10230 6151 10286 6160
rect 10046 5672 10102 5681
rect 10046 5607 10048 5616
rect 10100 5607 10102 5616
rect 10048 5578 10100 5584
rect 10336 5273 10364 12294
rect 10520 12220 10548 12786
rect 10428 12192 10548 12220
rect 10428 8945 10456 12192
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 10062 10548 11630
rect 10612 10470 10640 13280
rect 10692 12368 10744 12374
rect 10888 12345 10916 13670
rect 10692 12310 10744 12316
rect 10874 12336 10930 12345
rect 10704 10742 10732 12310
rect 10874 12271 10930 12280
rect 10980 11642 11008 21984
rect 11072 19825 11100 22052
rect 11058 19816 11114 19825
rect 11058 19751 11114 19760
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11072 18766 11100 19450
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 18426 11100 18702
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11164 17270 11192 28018
rect 11256 27606 11284 28562
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 11256 27130 11284 27542
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11256 25702 11284 26726
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 11256 25430 11284 25638
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 11256 24070 11284 25366
rect 11348 24682 11376 39520
rect 11808 37754 11836 39520
rect 12176 37890 12204 39520
rect 12176 37862 12388 37890
rect 11808 37726 12296 37754
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11428 34604 11480 34610
rect 11428 34546 11480 34552
rect 11440 34406 11468 34546
rect 11428 34400 11480 34406
rect 11428 34342 11480 34348
rect 11440 34202 11468 34342
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11428 34196 11480 34202
rect 11428 34138 11480 34144
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 12072 31816 12124 31822
rect 11978 31784 12034 31793
rect 12072 31758 12124 31764
rect 11978 31719 12034 31728
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11428 31204 11480 31210
rect 11428 31146 11480 31152
rect 11440 28082 11468 31146
rect 11532 31142 11560 31622
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11992 30326 12020 31719
rect 12084 30802 12112 31758
rect 12176 30870 12204 32302
rect 12164 30864 12216 30870
rect 12164 30806 12216 30812
rect 12072 30796 12124 30802
rect 12072 30738 12124 30744
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 11980 30320 12032 30326
rect 11980 30262 12032 30268
rect 11428 28076 11480 28082
rect 11428 28018 11480 28024
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11440 26790 11468 27406
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 11428 26308 11480 26314
rect 11428 26250 11480 26256
rect 11440 24818 11468 26250
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 11336 24676 11388 24682
rect 11336 24618 11388 24624
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11256 23186 11284 24006
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11256 21894 11284 23122
rect 11348 22438 11376 23190
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 19922 11284 21830
rect 11348 21554 11376 22374
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11334 21040 11390 21049
rect 11334 20975 11390 20984
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 15910 11100 16594
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15706 11100 15846
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13870 11100 14214
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 13530 11100 13806
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11164 12374 11192 16186
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11256 12714 11284 13262
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10888 11614 11008 11642
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9382 10548 9998
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8362 10456 8774
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10322 5264 10378 5273
rect 10322 5199 10378 5208
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4826 10180 4966
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 4457 10088 4626
rect 10046 4448 10102 4457
rect 10046 4383 10102 4392
rect 10152 4078 10180 4762
rect 10336 4706 10364 5199
rect 10244 4678 10364 4706
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10244 3602 10272 4678
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4282 10364 4558
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10428 3942 10456 8298
rect 10520 6361 10548 9318
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10612 8090 10640 8434
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10704 6769 10732 10678
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10796 10266 10824 10610
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10888 7313 10916 11614
rect 11060 11552 11112 11558
rect 10980 11500 11060 11506
rect 10980 11494 11112 11500
rect 10980 11478 11100 11494
rect 10980 10810 11008 11478
rect 11164 11286 11192 12174
rect 11256 11898 11284 12242
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11256 11354 11284 11834
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11256 10674 11284 11290
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 10968 8424 11020 8430
rect 11020 8384 11100 8412
rect 10968 8366 11020 8372
rect 10874 7304 10930 7313
rect 10874 7239 10930 7248
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6866 11008 7142
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11072 6798 11100 8384
rect 11150 7168 11206 7177
rect 11150 7103 11206 7112
rect 11060 6792 11112 6798
rect 10690 6760 10746 6769
rect 11060 6734 11112 6740
rect 10690 6695 10746 6704
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6361 11100 6598
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10874 6080 10930 6089
rect 10874 6015 10930 6024
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 5030 10640 5510
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10520 4729 10548 4966
rect 10506 4720 10562 4729
rect 10506 4655 10562 4664
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4146 10548 4422
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10520 3738 10548 4082
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10612 3641 10640 4966
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10704 4146 10732 4422
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 3738 10732 4082
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10598 3632 10654 3641
rect 10232 3596 10284 3602
rect 10598 3567 10654 3576
rect 10232 3538 10284 3544
rect 10782 3496 10838 3505
rect 10232 3460 10284 3466
rect 10782 3431 10838 3440
rect 10232 3402 10284 3408
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 2961 10180 3334
rect 10138 2952 10194 2961
rect 10138 2887 10194 2896
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10152 2446 10180 2518
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10244 2378 10272 3402
rect 10796 2582 10824 3431
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 9784 480 9812 2314
rect 9954 2272 10010 2281
rect 9954 2207 10010 2216
rect 9968 610 9996 2207
rect 10888 610 10916 6015
rect 11072 4826 11100 6122
rect 11164 5148 11192 7103
rect 11242 7032 11298 7041
rect 11242 6967 11298 6976
rect 11256 6458 11284 6967
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11348 6236 11376 20975
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11440 19990 11468 20402
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11440 19514 11468 19926
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11532 15722 11560 30262
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 12084 29782 12112 30738
rect 12072 29776 12124 29782
rect 11978 29744 12034 29753
rect 12072 29718 12124 29724
rect 11978 29679 12034 29688
rect 11992 29238 12020 29679
rect 11980 29232 12032 29238
rect 11978 29200 11980 29209
rect 12032 29200 12034 29209
rect 11978 29135 12034 29144
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 11992 28218 12020 28698
rect 12176 28558 12204 30806
rect 12268 30054 12296 37726
rect 12360 33017 12388 37862
rect 12544 35714 12572 39520
rect 13004 35714 13032 39520
rect 12544 35686 12664 35714
rect 12346 33008 12402 33017
rect 12346 32943 12402 32952
rect 12532 32768 12584 32774
rect 12532 32710 12584 32716
rect 12544 32434 12572 32710
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 12532 32292 12584 32298
rect 12532 32234 12584 32240
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 12452 31929 12480 32166
rect 12438 31920 12494 31929
rect 12348 31884 12400 31890
rect 12438 31855 12494 31864
rect 12348 31826 12400 31832
rect 12360 31278 12388 31826
rect 12544 31482 12572 32234
rect 12532 31476 12584 31482
rect 12532 31418 12584 31424
rect 12348 31272 12400 31278
rect 12348 31214 12400 31220
rect 12348 31136 12400 31142
rect 12400 31096 12480 31124
rect 12348 31078 12400 31084
rect 12452 30394 12480 31096
rect 12440 30388 12492 30394
rect 12440 30330 12492 30336
rect 12348 30184 12400 30190
rect 12348 30126 12400 30132
rect 12256 30048 12308 30054
rect 12360 30036 12388 30126
rect 12308 30008 12388 30036
rect 12256 29990 12308 29996
rect 12256 29776 12308 29782
rect 12256 29718 12308 29724
rect 12268 29170 12296 29718
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12164 28552 12216 28558
rect 12164 28494 12216 28500
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 12176 28150 12204 28494
rect 12164 28144 12216 28150
rect 12164 28086 12216 28092
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 12254 27568 12310 27577
rect 12254 27503 12310 27512
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11992 22234 12020 22374
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11900 21962 11928 22102
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11900 21622 11928 21898
rect 11992 21690 12020 22170
rect 12084 21690 12112 26998
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 12070 21584 12126 21593
rect 12070 21519 12126 21528
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 12084 21010 12112 21519
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11624 20602 11652 20810
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 12084 20534 12112 20946
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11624 15978 11652 16594
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11440 15694 11560 15722
rect 11440 13530 11468 15694
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15162 11560 15506
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11532 14074 11560 15098
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11440 12986 11468 13466
rect 11532 13326 11560 14010
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11532 12986 11560 13262
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11426 12744 11482 12753
rect 11426 12679 11428 12688
rect 11480 12679 11482 12688
rect 11428 12650 11480 12656
rect 11256 6208 11376 6236
rect 11256 5409 11284 6208
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5914 11376 6054
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11242 5400 11298 5409
rect 11242 5335 11298 5344
rect 11348 5234 11376 5510
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11164 5120 11284 5148
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4622 11100 4762
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4282 11100 4558
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11072 3602 11100 4218
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10966 2952 11022 2961
rect 11072 2922 11100 3538
rect 11164 3126 11192 3538
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 10966 2887 11022 2896
rect 11060 2916 11112 2922
rect 9956 604 10008 610
rect 9956 546 10008 552
rect 10140 604 10192 610
rect 10140 546 10192 552
rect 10600 604 10652 610
rect 10600 546 10652 552
rect 10876 604 10928 610
rect 10876 546 10928 552
rect 10152 480 10180 546
rect 10612 480 10640 546
rect 10980 480 11008 2887
rect 11060 2858 11112 2864
rect 11164 2446 11192 3062
rect 11256 2836 11284 5120
rect 11348 5030 11376 5170
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4690 11376 4966
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11348 3942 11376 4626
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3738 11376 3878
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11440 3194 11468 12650
rect 11532 12646 11560 12922
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11992 10713 12020 17206
rect 11978 10704 12034 10713
rect 11978 10639 12034 10648
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7546 11836 7890
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11992 6662 12020 6938
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11808 5370 11836 5646
rect 11992 5642 12020 6598
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11256 2808 11356 2836
rect 11440 2825 11468 2858
rect 12084 2825 12112 20470
rect 12176 15162 12204 22442
rect 12268 22030 12296 27503
rect 12360 26489 12388 30008
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 12544 28762 12572 29650
rect 12532 28756 12584 28762
rect 12532 28698 12584 28704
rect 12544 28665 12572 28698
rect 12530 28656 12586 28665
rect 12530 28591 12586 28600
rect 12532 28416 12584 28422
rect 12532 28358 12584 28364
rect 12544 26897 12572 28358
rect 12636 27577 12664 35686
rect 12820 35686 13032 35714
rect 12820 31385 12848 35686
rect 12900 32428 12952 32434
rect 12900 32370 12952 32376
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 12806 31376 12862 31385
rect 12806 31311 12862 31320
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12820 30598 12848 31214
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12820 29510 12848 30534
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12820 29170 12848 29446
rect 12912 29306 12940 32370
rect 13096 32026 13124 32370
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 13372 31362 13400 39520
rect 13740 35714 13768 39520
rect 13004 31334 13400 31362
rect 13464 35686 13768 35714
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12898 29200 12954 29209
rect 12808 29164 12860 29170
rect 12898 29135 12954 29144
rect 12808 29106 12860 29112
rect 12820 27674 12848 29106
rect 12912 29102 12940 29135
rect 12900 29096 12952 29102
rect 12900 29038 12952 29044
rect 12900 28960 12952 28966
rect 12900 28902 12952 28908
rect 12912 28422 12940 28902
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12808 27668 12860 27674
rect 12808 27610 12860 27616
rect 12622 27568 12678 27577
rect 12622 27503 12678 27512
rect 13004 27010 13032 31334
rect 13266 31240 13322 31249
rect 13084 31204 13136 31210
rect 13266 31175 13322 31184
rect 13084 31146 13136 31152
rect 13096 28762 13124 31146
rect 13280 31142 13308 31175
rect 13268 31136 13320 31142
rect 13268 31078 13320 31084
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 13082 28520 13138 28529
rect 13082 28455 13138 28464
rect 12728 26982 13032 27010
rect 12530 26888 12586 26897
rect 12530 26823 12586 26832
rect 12346 26480 12402 26489
rect 12346 26415 12402 26424
rect 12360 26058 12388 26415
rect 12360 26030 12664 26058
rect 12636 22098 12664 26030
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12360 21146 12388 21626
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12360 20602 12388 21082
rect 12452 21049 12480 21966
rect 12438 21040 12494 21049
rect 12438 20975 12494 20984
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 12268 15366 12296 15914
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12176 14958 12204 15098
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 14618 12204 14758
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12268 14414 12296 15302
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12176 14074 12204 14350
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12268 13462 12296 14350
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 12162 11792 12218 11801
rect 12162 11727 12164 11736
rect 12216 11727 12218 11736
rect 12164 11698 12216 11704
rect 12176 11558 12204 11698
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12176 5370 12204 5850
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 11328 2666 11356 2808
rect 11426 2816 11482 2825
rect 12070 2816 12126 2825
rect 11426 2751 11482 2760
rect 11622 2748 11918 2768
rect 12070 2751 12126 2760
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 12268 2666 12296 12854
rect 12360 7698 12388 20538
rect 12530 16688 12586 16697
rect 12530 16623 12586 16632
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16153 12480 16390
rect 12438 16144 12494 16153
rect 12438 16079 12494 16088
rect 12438 12336 12494 12345
rect 12438 12271 12494 12280
rect 12452 11898 12480 12271
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11694 12572 16623
rect 12728 15337 12756 26982
rect 12990 22536 13046 22545
rect 13096 22506 13124 28455
rect 13174 26888 13230 26897
rect 13174 26823 13230 26832
rect 12990 22471 13046 22480
rect 13084 22500 13136 22506
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12820 22166 12848 22374
rect 13004 22234 13032 22471
rect 13084 22442 13136 22448
rect 13188 22386 13216 26823
rect 13096 22358 13216 22386
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12820 21554 12848 22102
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12714 15328 12770 15337
rect 12714 15263 12770 15272
rect 12912 15094 12940 22034
rect 13004 21690 13032 22170
rect 13096 21962 13124 22358
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 13188 21690 13216 21966
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12728 14618 12756 14962
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 14618 12848 14826
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12728 13938 12756 14554
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12102 12664 12582
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11762 12664 12038
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12636 11354 12664 11698
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12360 7670 12572 7698
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12452 6730 12480 7482
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12544 6610 12572 7670
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12360 6582 12572 6610
rect 12360 2961 12388 6582
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12544 6118 12572 6190
rect 12636 6186 12664 6870
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4593 12664 4966
rect 12622 4584 12678 4593
rect 12622 4519 12678 4528
rect 12728 4486 12756 6734
rect 12820 6662 12848 13398
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5914 12848 6190
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12820 5710 12848 5850
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 4480 12768 4486
rect 12438 4448 12494 4457
rect 12716 4422 12768 4428
rect 12438 4383 12494 4392
rect 12452 3194 12480 4383
rect 12622 4040 12678 4049
rect 12622 3975 12678 3984
rect 12636 3942 12664 3975
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12622 3632 12678 3641
rect 12532 3596 12584 3602
rect 12622 3567 12678 3576
rect 12532 3538 12584 3544
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12346 2952 12402 2961
rect 12402 2910 12480 2938
rect 12346 2887 12402 2896
rect 12360 2827 12388 2887
rect 11328 2638 11376 2666
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11348 480 11376 2638
rect 12084 2638 12296 2666
rect 12452 2650 12480 2910
rect 12440 2644 12492 2650
rect 11886 2544 11942 2553
rect 11886 2479 11888 2488
rect 11940 2479 11942 2488
rect 11888 2450 11940 2456
rect 12084 1578 12112 2638
rect 12440 2586 12492 2592
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 11808 1550 12112 1578
rect 11808 480 11836 1550
rect 12176 480 12204 2518
rect 12544 480 12572 3538
rect 12636 2650 12664 3567
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12728 3369 12756 3470
rect 12714 3360 12770 3369
rect 12714 3295 12770 3304
rect 12716 3120 12768 3126
rect 12820 3097 12848 5510
rect 12912 5370 12940 14758
rect 13004 13802 13032 21626
rect 13174 17776 13230 17785
rect 13174 17711 13230 17720
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13096 13870 13124 15030
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12912 5166 12940 5306
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 13004 4146 13032 13466
rect 13096 13462 13124 13806
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13096 3641 13124 11630
rect 13082 3632 13138 3641
rect 13188 3602 13216 17711
rect 13280 5778 13308 31078
rect 13464 30682 13492 35686
rect 13820 32020 13872 32026
rect 13820 31962 13872 31968
rect 13464 30654 13584 30682
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 13464 30433 13492 30534
rect 13450 30424 13506 30433
rect 13450 30359 13506 30368
rect 13452 30252 13504 30258
rect 13452 30194 13504 30200
rect 13464 30054 13492 30194
rect 13452 30048 13504 30054
rect 13452 29990 13504 29996
rect 13464 29646 13492 29990
rect 13452 29640 13504 29646
rect 13452 29582 13504 29588
rect 13464 29306 13492 29582
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13372 22030 13400 22578
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13372 13530 13400 21830
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6458 13400 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13360 6112 13412 6118
rect 13464 6066 13492 28970
rect 13556 18873 13584 30654
rect 13832 30326 13860 31962
rect 13820 30320 13872 30326
rect 13820 30262 13872 30268
rect 14200 29034 14228 39520
rect 14568 37210 14596 39520
rect 14936 39494 15056 39520
rect 14568 37182 14688 37210
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14660 32337 14688 37182
rect 14646 32328 14702 32337
rect 14646 32263 14702 32272
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14188 29028 14240 29034
rect 14188 28970 14240 28976
rect 15028 28529 15056 39494
rect 15396 35290 15424 39520
rect 15384 35284 15436 35290
rect 15384 35226 15436 35232
rect 15764 31249 15792 39520
rect 15750 31240 15806 31249
rect 15750 31175 15806 31184
rect 15014 28520 15070 28529
rect 15014 28455 15070 28464
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13648 21690 13676 21966
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 13542 18864 13598 18873
rect 13542 18799 13598 18808
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13412 6060 13492 6066
rect 13360 6054 13492 6060
rect 13372 6038 13492 6054
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13280 5370 13308 5714
rect 13464 5681 13492 6038
rect 13450 5672 13506 5681
rect 13450 5607 13506 5616
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13556 4808 13584 9415
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13280 4780 13584 4808
rect 13082 3567 13138 3576
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13280 3482 13308 4780
rect 13358 4720 13414 4729
rect 13358 4655 13414 4664
rect 13004 3454 13308 3482
rect 12716 3062 12768 3068
rect 12806 3088 12862 3097
rect 12728 2990 12756 3062
rect 12806 3023 12862 3032
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 13004 480 13032 3454
rect 13372 480 13400 4655
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13464 2854 13492 2994
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13464 2446 13492 2790
rect 13452 2440 13504 2446
rect 13648 2417 13676 6598
rect 13740 2990 13768 11494
rect 13832 3058 13860 13738
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14186 10704 14242 10713
rect 14186 10639 14242 10648
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13452 2382 13504 2388
rect 13634 2408 13690 2417
rect 13634 2343 13690 2352
rect 13726 2000 13782 2009
rect 13726 1935 13782 1944
rect 13740 480 13768 1935
rect 14200 480 14228 10639
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 15750 5672 15806 5681
rect 15750 5607 15806 5616
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14646 5128 14702 5137
rect 14646 5063 14702 5072
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 5063
rect 15382 3632 15438 3641
rect 15382 3567 15438 3576
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 2994
rect 15396 480 15424 3567
rect 15764 480 15792 5607
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 1582 38664 1638 38720
rect 1490 34584 1546 34640
rect 1674 36352 1730 36408
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3330 35672 3386 35728
rect 2962 35536 3018 35592
rect 1582 34040 1638 34096
rect 2410 33516 2466 33552
rect 2410 33496 2412 33516
rect 2412 33496 2464 33516
rect 2464 33496 2466 33516
rect 2226 33224 2282 33280
rect 2042 32408 2098 32464
rect 2226 31864 2282 31920
rect 1582 31592 1638 31648
rect 2042 30132 2044 30152
rect 2044 30132 2096 30152
rect 2096 30132 2098 30152
rect 2042 30096 2098 30132
rect 1674 29280 1730 29336
rect 1582 26968 1638 27024
rect 2226 22636 2282 22672
rect 2226 22616 2228 22636
rect 2228 22616 2280 22636
rect 2280 22616 2282 22636
rect 1674 22208 1730 22264
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 4066 34740 4122 34776
rect 4066 34720 4068 34740
rect 4068 34720 4120 34740
rect 4120 34720 4122 34740
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 2778 24520 2834 24576
rect 2502 24112 2558 24168
rect 1582 19896 1638 19952
rect 2778 19624 2834 19680
rect 1674 17584 1730 17640
rect 3054 19624 3110 19680
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 1398 16652 1454 16688
rect 1398 16632 1400 16652
rect 1400 16632 1452 16652
rect 1452 16632 1454 16652
rect 1674 15136 1730 15192
rect 1674 13948 1676 13968
rect 1676 13948 1728 13968
rect 1728 13948 1730 13968
rect 1674 13912 1730 13948
rect 1582 12824 1638 12880
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3698 18164 3700 18184
rect 3700 18164 3752 18184
rect 3752 18164 3754 18184
rect 3698 18128 3754 18164
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3974 17196 4030 17232
rect 3974 17176 3976 17196
rect 3976 17176 4028 17196
rect 4028 17176 4030 17196
rect 3974 17060 4030 17096
rect 3974 17040 3976 17060
rect 3976 17040 4028 17060
rect 4028 17040 4030 17060
rect 3330 16496 3386 16552
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3790 15852 3792 15872
rect 3792 15852 3844 15872
rect 3844 15852 3846 15872
rect 3790 15816 3846 15852
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3790 14764 3792 14784
rect 3792 14764 3844 14784
rect 3844 14764 3846 14784
rect 3790 14728 3846 14764
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 4434 30232 4490 30288
rect 4802 24112 4858 24168
rect 5354 31320 5410 31376
rect 4986 30132 4988 30152
rect 4988 30132 5040 30152
rect 5040 30132 5042 30152
rect 4986 30096 5042 30132
rect 5170 29688 5226 29744
rect 5262 29144 5318 29200
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 5722 31320 5778 31376
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6090 33260 6092 33280
rect 6092 33260 6144 33280
rect 6144 33260 6146 33280
rect 6090 33224 6146 33260
rect 7470 35436 7472 35456
rect 7472 35436 7524 35456
rect 7524 35436 7526 35456
rect 7470 35400 7526 35436
rect 8022 35708 8024 35728
rect 8024 35708 8076 35728
rect 8076 35708 8078 35728
rect 8022 35672 8078 35708
rect 7562 34720 7618 34776
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 7286 33496 7342 33552
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 5998 30640 6054 30696
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6826 30912 6882 30968
rect 6826 30776 6882 30832
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6090 27512 6146 27568
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 5078 24248 5134 24304
rect 5446 21392 5502 21448
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 5170 19760 5226 19816
rect 2226 11620 2282 11656
rect 2226 11600 2228 11620
rect 2228 11600 2280 11620
rect 2280 11600 2282 11620
rect 1674 10512 1730 10568
rect 1490 8064 1546 8120
rect 2410 7948 2466 7984
rect 2410 7928 2412 7948
rect 2412 7928 2464 7948
rect 2464 7928 2466 7948
rect 2870 8336 2926 8392
rect 1582 5752 1638 5808
rect 2410 6296 2466 6352
rect 1490 4120 1546 4176
rect 1398 1400 1454 1456
rect 1674 3440 1730 3496
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 5078 18844 5080 18864
rect 5080 18844 5132 18864
rect 5132 18844 5134 18864
rect 5078 18808 5134 18844
rect 4894 12280 4950 12336
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3238 6160 3294 6216
rect 2778 4528 2834 4584
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 5078 15816 5134 15872
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6550 19760 6606 19816
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 5538 14728 5594 14784
rect 5078 12688 5134 12744
rect 4894 9696 4950 9752
rect 4434 9560 4490 9616
rect 4710 8336 4766 8392
rect 5078 7792 5134 7848
rect 5354 7248 5410 7304
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3330 3712 3386 3768
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 4250 4120 4306 4176
rect 3882 4004 3938 4040
rect 4526 4256 4582 4312
rect 3882 3984 3884 4004
rect 3884 3984 3936 4004
rect 3936 3984 3938 4004
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4342 3848 4398 3904
rect 4158 2896 4214 2952
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 3330 1672 3386 1728
rect 2962 1536 3018 1592
rect 3790 1400 3846 1456
rect 4986 4120 5042 4176
rect 4802 3984 4858 4040
rect 4710 3440 4766 3496
rect 5630 6432 5686 6488
rect 5538 5108 5540 5128
rect 5540 5108 5592 5128
rect 5592 5108 5594 5128
rect 5538 5072 5594 5108
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 7010 29824 7066 29880
rect 7470 29824 7526 29880
rect 7470 28600 7526 28656
rect 7286 26852 7342 26888
rect 7286 26832 7288 26852
rect 7288 26832 7340 26852
rect 7340 26832 7342 26852
rect 7378 26424 7434 26480
rect 7102 24656 7158 24712
rect 6918 19216 6974 19272
rect 6826 18672 6882 18728
rect 7010 17176 7066 17232
rect 6090 9968 6146 10024
rect 5998 6432 6054 6488
rect 5998 6296 6054 6352
rect 5722 4800 5778 4856
rect 5906 5244 5908 5264
rect 5908 5244 5960 5264
rect 5960 5244 5962 5264
rect 5906 5208 5962 5244
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 7654 29688 7710 29744
rect 7654 29416 7710 29472
rect 8206 34720 8262 34776
rect 8114 29008 8170 29064
rect 7838 28600 7894 28656
rect 7746 28500 7748 28520
rect 7748 28500 7800 28520
rect 7800 28500 7802 28520
rect 7746 28464 7802 28500
rect 7654 24556 7656 24576
rect 7656 24556 7708 24576
rect 7708 24556 7710 24576
rect 7654 24520 7710 24556
rect 7286 20032 7342 20088
rect 7286 19760 7342 19816
rect 7378 16632 7434 16688
rect 7838 22616 7894 22672
rect 7746 22480 7802 22536
rect 7562 20168 7618 20224
rect 7562 18672 7618 18728
rect 8482 34620 8484 34640
rect 8484 34620 8536 34640
rect 8536 34620 8538 34640
rect 8482 34584 8538 34620
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 9218 35536 9274 35592
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8482 32272 8538 32328
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8390 31864 8446 31920
rect 8666 31728 8722 31784
rect 8574 30932 8630 30968
rect 8574 30912 8576 30932
rect 8576 30912 8628 30932
rect 8628 30912 8630 30932
rect 8758 30776 8814 30832
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8850 30232 8906 30288
rect 8390 30096 8446 30152
rect 8574 29588 8576 29608
rect 8576 29588 8628 29608
rect 8628 29588 8630 29608
rect 8574 29552 8630 29588
rect 8482 29164 8538 29200
rect 8482 29144 8484 29164
rect 8484 29144 8536 29164
rect 8536 29144 8538 29164
rect 8390 26188 8392 26208
rect 8392 26188 8444 26208
rect 8444 26188 8446 26208
rect 8390 26152 8446 26188
rect 8666 29008 8722 29064
rect 8298 24792 8354 24848
rect 8482 24792 8538 24848
rect 8390 24656 8446 24712
rect 9770 33768 9826 33824
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 9494 31320 9550 31376
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 10230 34584 10286 34640
rect 9770 30368 9826 30424
rect 9678 30132 9680 30152
rect 9680 30132 9732 30152
rect 9732 30132 9734 30152
rect 9678 30096 9734 30132
rect 9586 29552 9642 29608
rect 9678 29416 9734 29472
rect 9862 29008 9918 29064
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8022 20032 8078 20088
rect 7102 12688 7158 12744
rect 7010 11736 7066 11792
rect 7010 9560 7066 9616
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6734 8336 6790 8392
rect 6734 6976 6790 7032
rect 6090 3884 6092 3904
rect 6092 3884 6144 3904
rect 6144 3884 6146 3904
rect 6090 3848 6146 3884
rect 6090 3712 6146 3768
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6826 6704 6882 6760
rect 7286 8880 7342 8936
rect 7010 7248 7066 7304
rect 7378 6840 7434 6896
rect 6826 5752 6882 5808
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6182 3576 6238 3632
rect 5814 1400 5870 1456
rect 6642 3168 6698 3224
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6274 2372 6330 2408
rect 6274 2352 6276 2372
rect 6276 2352 6328 2372
rect 6328 2352 6330 2372
rect 7102 4528 7158 4584
rect 7470 6024 7526 6080
rect 7746 11600 7802 11656
rect 8114 19352 8170 19408
rect 8114 17176 8170 17232
rect 8022 16652 8078 16688
rect 8022 16632 8024 16652
rect 8024 16632 8076 16652
rect 8076 16632 8078 16652
rect 7930 11328 7986 11384
rect 8390 12280 8446 12336
rect 8666 20984 8722 21040
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 9862 24812 9918 24848
rect 9862 24792 9864 24812
rect 9864 24792 9916 24812
rect 9916 24792 9918 24812
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8758 17992 8814 18048
rect 8666 16496 8722 16552
rect 8758 8880 8814 8936
rect 7838 7148 7840 7168
rect 7840 7148 7892 7168
rect 7892 7148 7894 7168
rect 7838 7112 7894 7148
rect 7838 6196 7840 6216
rect 7840 6196 7892 6216
rect 7892 6196 7894 6216
rect 7838 6160 7894 6196
rect 7838 5616 7894 5672
rect 7746 3440 7802 3496
rect 7746 3032 7802 3088
rect 7654 1536 7710 1592
rect 8390 7112 8446 7168
rect 8206 6296 8262 6352
rect 8022 4392 8078 4448
rect 8206 4392 8262 4448
rect 8022 2508 8078 2544
rect 8022 2488 8024 2508
rect 8024 2488 8076 2508
rect 8076 2488 8078 2508
rect 8482 4120 8538 4176
rect 8666 6840 8722 6896
rect 8666 6704 8722 6760
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 9218 19352 9274 19408
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 9678 24520 9734 24576
rect 9678 24268 9734 24304
rect 9678 24248 9680 24268
rect 9680 24248 9732 24268
rect 9732 24248 9734 24268
rect 9678 22072 9734 22128
rect 9678 21800 9734 21856
rect 10046 29416 10102 29472
rect 10506 32408 10562 32464
rect 10322 30640 10378 30696
rect 10322 30368 10378 30424
rect 10506 29960 10562 30016
rect 10506 29824 10562 29880
rect 10782 32988 10784 33008
rect 10784 32988 10836 33008
rect 10836 32988 10838 33008
rect 10782 32952 10838 32988
rect 10874 31884 10930 31920
rect 10874 31864 10876 31884
rect 10876 31864 10928 31884
rect 10928 31864 10930 31884
rect 11150 30368 11206 30424
rect 11150 30096 11206 30152
rect 11150 29572 11206 29608
rect 11150 29552 11152 29572
rect 11152 29552 11204 29572
rect 11204 29552 11206 29572
rect 10046 21412 10102 21448
rect 10046 21392 10048 21412
rect 10048 21392 10100 21412
rect 10100 21392 10102 21412
rect 9494 17040 9550 17096
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 9218 15000 9274 15056
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 9034 8336 9090 8392
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8942 7248 8998 7304
rect 8942 6724 8998 6760
rect 8942 6704 8944 6724
rect 8944 6704 8996 6724
rect 8996 6704 8998 6724
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 9678 16632 9734 16688
rect 10138 20204 10140 20224
rect 10140 20204 10192 20224
rect 10192 20204 10194 20224
rect 10138 20168 10194 20204
rect 10138 20032 10194 20088
rect 9862 18808 9918 18864
rect 10046 17992 10102 18048
rect 9862 16088 9918 16144
rect 10506 21528 10562 21584
rect 10690 19760 10746 19816
rect 10874 19388 10876 19408
rect 10876 19388 10928 19408
rect 10928 19388 10930 19408
rect 10874 19352 10930 19388
rect 10782 19216 10838 19272
rect 10598 17720 10654 17776
rect 10138 13912 10194 13968
rect 9586 11328 9642 11384
rect 9954 12280 10010 12336
rect 9678 7792 9734 7848
rect 9402 6704 9458 6760
rect 8758 4256 8814 4312
rect 8574 3188 8630 3224
rect 8574 3168 8576 3188
rect 8576 3168 8628 3188
rect 8628 3168 8630 3188
rect 8666 1944 8722 2000
rect 8758 1672 8814 1728
rect 9678 5752 9734 5808
rect 9954 7928 10010 7984
rect 10506 16632 10562 16688
rect 10690 16088 10746 16144
rect 10138 9424 10194 9480
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 9402 5364 9458 5400
rect 9402 5344 9404 5364
rect 9404 5344 9456 5364
rect 9456 5344 9458 5364
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 9034 4020 9036 4040
rect 9036 4020 9088 4040
rect 9088 4020 9090 4040
rect 9034 3984 9090 4020
rect 9402 3304 9458 3360
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9402 2760 9458 2816
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9770 2624 9826 2680
rect 10230 6196 10232 6216
rect 10232 6196 10284 6216
rect 10284 6196 10286 6216
rect 10230 6160 10286 6196
rect 10046 5636 10102 5672
rect 10046 5616 10048 5636
rect 10048 5616 10100 5636
rect 10100 5616 10102 5636
rect 10874 12280 10930 12336
rect 11058 19760 11114 19816
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11978 31728 12034 31784
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11334 20984 11390 21040
rect 10414 8880 10470 8936
rect 10322 5208 10378 5264
rect 10046 4392 10102 4448
rect 10874 7248 10930 7304
rect 11150 7112 11206 7168
rect 10690 6704 10746 6760
rect 10506 6296 10562 6352
rect 11058 6296 11114 6352
rect 10874 6024 10930 6080
rect 10506 4664 10562 4720
rect 10598 3576 10654 3632
rect 10782 3440 10838 3496
rect 10138 2896 10194 2952
rect 9954 2216 10010 2272
rect 11242 6976 11298 7032
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11978 29688 12034 29744
rect 11978 29180 11980 29200
rect 11980 29180 12032 29200
rect 12032 29180 12034 29200
rect 11978 29144 12034 29180
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 12346 32952 12402 33008
rect 12438 31864 12494 31920
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 12254 27512 12310 27568
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 12070 21528 12126 21584
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11426 12708 11482 12744
rect 11426 12688 11428 12708
rect 11428 12688 11480 12708
rect 11480 12688 11482 12708
rect 11242 5344 11298 5400
rect 10966 2896 11022 2952
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11978 10648 12034 10704
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 12530 28600 12586 28656
rect 12806 31320 12862 31376
rect 12898 29144 12954 29200
rect 12622 27512 12678 27568
rect 13266 31184 13322 31240
rect 13082 28464 13138 28520
rect 12530 26832 12586 26888
rect 12346 26424 12402 26480
rect 12438 20984 12494 21040
rect 12162 11756 12218 11792
rect 12162 11736 12164 11756
rect 12164 11736 12216 11756
rect 12216 11736 12218 11756
rect 11426 2760 11482 2816
rect 12070 2760 12126 2816
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12530 16632 12586 16688
rect 12438 16088 12494 16144
rect 12438 12280 12494 12336
rect 12990 22480 13046 22536
rect 13174 26832 13230 26888
rect 12714 15272 12770 15328
rect 12622 4528 12678 4584
rect 12438 4392 12494 4448
rect 12622 3984 12678 4040
rect 12622 3576 12678 3632
rect 12346 2896 12402 2952
rect 11886 2508 11942 2544
rect 11886 2488 11888 2508
rect 11888 2488 11940 2508
rect 11940 2488 11942 2508
rect 12714 3304 12770 3360
rect 13174 17720 13230 17776
rect 13082 3576 13138 3632
rect 13450 30368 13506 30424
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14646 32272 14702 32328
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 15750 31184 15806 31240
rect 15014 28464 15070 28520
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 13542 18808 13598 18864
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 13542 9424 13598 9480
rect 13450 5616 13506 5672
rect 13358 4664 13414 4720
rect 12806 3032 12862 3088
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14186 10648 14242 10704
rect 13634 2352 13690 2408
rect 13726 1944 13782 2000
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 15750 5616 15806 5672
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14646 5072 14702 5128
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 15382 3576 15438 3632
<< metal3 >>
rect 0 38722 480 38752
rect 1577 38722 1643 38725
rect 0 38720 1643 38722
rect 0 38664 1582 38720
rect 1638 38664 1643 38720
rect 0 38662 1643 38664
rect 0 38632 480 38662
rect 1577 38659 1643 38662
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 0 36410 480 36440
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 1669 36410 1735 36413
rect 0 36408 1735 36410
rect 0 36352 1674 36408
rect 1730 36352 1735 36408
rect 0 36350 1735 36352
rect 0 36320 480 36350
rect 1669 36347 1735 36350
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 3325 35730 3391 35733
rect 8017 35730 8083 35733
rect 3325 35728 8083 35730
rect 3325 35672 3330 35728
rect 3386 35672 8022 35728
rect 8078 35672 8083 35728
rect 3325 35670 8083 35672
rect 3325 35667 3391 35670
rect 8017 35667 8083 35670
rect 2957 35594 3023 35597
rect 9213 35594 9279 35597
rect 2957 35592 9279 35594
rect 2957 35536 2962 35592
rect 3018 35536 9218 35592
rect 9274 35536 9279 35592
rect 2957 35534 9279 35536
rect 2957 35531 3023 35534
rect 9213 35531 9279 35534
rect 7465 35458 7531 35461
rect 7598 35458 7604 35460
rect 7465 35456 7604 35458
rect 7465 35400 7470 35456
rect 7526 35400 7604 35456
rect 7465 35398 7604 35400
rect 7465 35395 7531 35398
rect 7598 35396 7604 35398
rect 7668 35396 7674 35460
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 4061 34778 4127 34781
rect 7557 34778 7623 34781
rect 4061 34776 7623 34778
rect 4061 34720 4066 34776
rect 4122 34720 7562 34776
rect 7618 34720 7623 34776
rect 4061 34718 7623 34720
rect 4061 34715 4127 34718
rect 7557 34715 7623 34718
rect 8201 34778 8267 34781
rect 8201 34776 8770 34778
rect 8201 34720 8206 34776
rect 8262 34720 8770 34776
rect 8201 34718 8770 34720
rect 8201 34715 8267 34718
rect 1485 34642 1551 34645
rect 8477 34642 8543 34645
rect 1485 34640 8543 34642
rect 1485 34584 1490 34640
rect 1546 34584 8482 34640
rect 8538 34584 8543 34640
rect 1485 34582 8543 34584
rect 8710 34642 8770 34718
rect 10225 34642 10291 34645
rect 8710 34640 10291 34642
rect 8710 34584 10230 34640
rect 10286 34584 10291 34640
rect 8710 34582 10291 34584
rect 1485 34579 1551 34582
rect 8477 34579 8543 34582
rect 10225 34579 10291 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 0 34098 480 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 480 34038
rect 1577 34035 1643 34038
rect 9622 33764 9628 33828
rect 9692 33826 9698 33828
rect 9765 33826 9831 33829
rect 9692 33824 9831 33826
rect 9692 33768 9770 33824
rect 9826 33768 9831 33824
rect 9692 33766 9831 33768
rect 9692 33764 9698 33766
rect 9765 33763 9831 33766
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 2405 33554 2471 33557
rect 7281 33554 7347 33557
rect 2405 33552 7347 33554
rect 2405 33496 2410 33552
rect 2466 33496 7286 33552
rect 7342 33496 7347 33552
rect 2405 33494 7347 33496
rect 2405 33491 2471 33494
rect 7281 33491 7347 33494
rect 2221 33282 2287 33285
rect 6085 33282 6151 33285
rect 2221 33280 6151 33282
rect 2221 33224 2226 33280
rect 2282 33224 6090 33280
rect 6146 33224 6151 33280
rect 2221 33222 6151 33224
rect 2221 33219 2287 33222
rect 6085 33219 6151 33222
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 10777 33010 10843 33013
rect 12341 33010 12407 33013
rect 10777 33008 12407 33010
rect 10777 32952 10782 33008
rect 10838 32952 12346 33008
rect 12402 32952 12407 33008
rect 10777 32950 12407 32952
rect 10777 32947 10843 32950
rect 12341 32947 12407 32950
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 2037 32466 2103 32469
rect 10501 32466 10567 32469
rect 2037 32464 10567 32466
rect 2037 32408 2042 32464
rect 2098 32408 10506 32464
rect 10562 32408 10567 32464
rect 2037 32406 10567 32408
rect 2037 32403 2103 32406
rect 10501 32403 10567 32406
rect 8477 32330 8543 32333
rect 14641 32330 14707 32333
rect 8477 32328 14707 32330
rect 8477 32272 8482 32328
rect 8538 32272 14646 32328
rect 14702 32272 14707 32328
rect 8477 32270 14707 32272
rect 8477 32267 8543 32270
rect 14641 32267 14707 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 2221 31922 2287 31925
rect 8385 31922 8451 31925
rect 2221 31920 8451 31922
rect 2221 31864 2226 31920
rect 2282 31864 8390 31920
rect 8446 31864 8451 31920
rect 2221 31862 8451 31864
rect 2221 31859 2287 31862
rect 8385 31859 8451 31862
rect 10869 31922 10935 31925
rect 12433 31922 12499 31925
rect 10869 31920 12499 31922
rect 10869 31864 10874 31920
rect 10930 31864 12438 31920
rect 12494 31864 12499 31920
rect 10869 31862 12499 31864
rect 10869 31859 10935 31862
rect 12433 31859 12499 31862
rect 8661 31786 8727 31789
rect 11973 31786 12039 31789
rect 8661 31784 12039 31786
rect 8661 31728 8666 31784
rect 8722 31728 11978 31784
rect 12034 31728 12039 31784
rect 8661 31726 12039 31728
rect 8661 31723 8727 31726
rect 11973 31723 12039 31726
rect 0 31650 480 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 480 31590
rect 1577 31587 1643 31590
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 5349 31378 5415 31381
rect 5717 31378 5783 31381
rect 9489 31378 9555 31381
rect 12801 31378 12867 31381
rect 5349 31376 12867 31378
rect 5349 31320 5354 31376
rect 5410 31320 5722 31376
rect 5778 31320 9494 31376
rect 9550 31320 12806 31376
rect 12862 31320 12867 31376
rect 5349 31318 12867 31320
rect 5349 31315 5415 31318
rect 5717 31315 5783 31318
rect 9489 31315 9555 31318
rect 12801 31315 12867 31318
rect 13261 31242 13327 31245
rect 15745 31242 15811 31245
rect 13261 31240 15811 31242
rect 13261 31184 13266 31240
rect 13322 31184 15750 31240
rect 15806 31184 15811 31240
rect 13261 31182 15811 31184
rect 13261 31179 13327 31182
rect 15745 31179 15811 31182
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 6821 30970 6887 30973
rect 8569 30970 8635 30973
rect 6821 30968 8635 30970
rect 6821 30912 6826 30968
rect 6882 30912 8574 30968
rect 8630 30912 8635 30968
rect 6821 30910 8635 30912
rect 6821 30907 6887 30910
rect 8569 30907 8635 30910
rect 6821 30834 6887 30837
rect 8753 30834 8819 30837
rect 6821 30832 8819 30834
rect 6821 30776 6826 30832
rect 6882 30776 8758 30832
rect 8814 30776 8819 30832
rect 6821 30774 8819 30776
rect 6821 30771 6887 30774
rect 8753 30771 8819 30774
rect 5993 30698 6059 30701
rect 10317 30698 10383 30701
rect 5993 30696 10383 30698
rect 5993 30640 5998 30696
rect 6054 30640 10322 30696
rect 10378 30640 10383 30696
rect 5993 30638 10383 30640
rect 5993 30635 6059 30638
rect 10317 30635 10383 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 9765 30426 9831 30429
rect 10317 30426 10383 30429
rect 9765 30424 10383 30426
rect 9765 30368 9770 30424
rect 9826 30368 10322 30424
rect 10378 30368 10383 30424
rect 9765 30366 10383 30368
rect 9765 30363 9831 30366
rect 10317 30363 10383 30366
rect 11145 30426 11211 30429
rect 13445 30426 13511 30429
rect 11145 30424 13738 30426
rect 11145 30368 11150 30424
rect 11206 30368 13450 30424
rect 13506 30368 13738 30424
rect 11145 30366 13738 30368
rect 11145 30363 11211 30366
rect 13445 30363 13511 30366
rect 4429 30290 4495 30293
rect 8845 30290 8911 30293
rect 4429 30288 8911 30290
rect 4429 30232 4434 30288
rect 4490 30232 8850 30288
rect 8906 30232 8911 30288
rect 4429 30230 8911 30232
rect 4429 30227 4495 30230
rect 8845 30227 8911 30230
rect 2037 30154 2103 30157
rect 4981 30154 5047 30157
rect 8385 30154 8451 30157
rect 2037 30152 8451 30154
rect 2037 30096 2042 30152
rect 2098 30096 4986 30152
rect 5042 30096 8390 30152
rect 8446 30096 8451 30152
rect 2037 30094 8451 30096
rect 2037 30091 2103 30094
rect 4981 30091 5047 30094
rect 8385 30091 8451 30094
rect 9673 30154 9739 30157
rect 11145 30154 11211 30157
rect 9673 30152 11211 30154
rect 9673 30096 9678 30152
rect 9734 30096 11150 30152
rect 11206 30096 11211 30152
rect 9673 30094 11211 30096
rect 9673 30091 9739 30094
rect 11145 30091 11211 30094
rect 10501 30018 10567 30021
rect 6686 30016 10567 30018
rect 6686 29960 10506 30016
rect 10562 29960 10567 30016
rect 6686 29958 10567 29960
rect 13678 30018 13738 30366
rect 15520 30018 16000 30048
rect 13678 29958 16000 30018
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 5165 29746 5231 29749
rect 6686 29746 6746 29958
rect 10501 29955 10567 29958
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 7005 29882 7071 29885
rect 7465 29882 7531 29885
rect 10501 29882 10567 29885
rect 7005 29880 10567 29882
rect 7005 29824 7010 29880
rect 7066 29824 7470 29880
rect 7526 29824 10506 29880
rect 10562 29824 10567 29880
rect 7005 29822 10567 29824
rect 7005 29819 7071 29822
rect 7465 29819 7531 29822
rect 10501 29819 10567 29822
rect 5165 29744 6746 29746
rect 5165 29688 5170 29744
rect 5226 29688 6746 29744
rect 5165 29686 6746 29688
rect 7649 29746 7715 29749
rect 11973 29746 12039 29749
rect 7649 29744 12039 29746
rect 7649 29688 7654 29744
rect 7710 29688 11978 29744
rect 12034 29688 12039 29744
rect 7649 29686 12039 29688
rect 5165 29683 5231 29686
rect 7649 29683 7715 29686
rect 11973 29683 12039 29686
rect 8569 29610 8635 29613
rect 9581 29610 9647 29613
rect 11145 29610 11211 29613
rect 8569 29608 11211 29610
rect 8569 29552 8574 29608
rect 8630 29552 9586 29608
rect 9642 29552 11150 29608
rect 11206 29552 11211 29608
rect 8569 29550 11211 29552
rect 8569 29547 8635 29550
rect 9581 29547 9647 29550
rect 11145 29547 11211 29550
rect 7649 29476 7715 29477
rect 9673 29476 9739 29477
rect 7598 29474 7604 29476
rect 7558 29414 7604 29474
rect 7668 29472 7715 29476
rect 7710 29416 7715 29472
rect 7598 29412 7604 29414
rect 7668 29412 7715 29416
rect 9622 29412 9628 29476
rect 9692 29474 9739 29476
rect 10041 29474 10107 29477
rect 9692 29472 9784 29474
rect 9734 29416 9784 29472
rect 9692 29414 9784 29416
rect 9998 29472 10107 29474
rect 9998 29416 10046 29472
rect 10102 29416 10107 29472
rect 9692 29412 9739 29414
rect 7649 29411 7715 29412
rect 9673 29411 9739 29412
rect 9998 29411 10107 29416
rect 3610 29408 3930 29409
rect 0 29338 480 29368
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 1669 29338 1735 29341
rect 0 29336 1735 29338
rect 0 29280 1674 29336
rect 1730 29280 1735 29336
rect 0 29278 1735 29280
rect 0 29248 480 29278
rect 1669 29275 1735 29278
rect 5257 29202 5323 29205
rect 8477 29202 8543 29205
rect 5257 29200 8543 29202
rect 5257 29144 5262 29200
rect 5318 29144 8482 29200
rect 8538 29144 8543 29200
rect 5257 29142 8543 29144
rect 5257 29139 5323 29142
rect 8477 29139 8543 29142
rect 8109 29066 8175 29069
rect 8661 29066 8727 29069
rect 8109 29064 8727 29066
rect 8109 29008 8114 29064
rect 8170 29008 8666 29064
rect 8722 29008 8727 29064
rect 8109 29006 8727 29008
rect 8109 29003 8175 29006
rect 8661 29003 8727 29006
rect 9857 29066 9923 29069
rect 9998 29066 10058 29411
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 11973 29202 12039 29205
rect 12893 29202 12959 29205
rect 11973 29200 12959 29202
rect 11973 29144 11978 29200
rect 12034 29144 12898 29200
rect 12954 29144 12959 29200
rect 11973 29142 12959 29144
rect 11973 29139 12039 29142
rect 12893 29139 12959 29142
rect 9857 29064 10058 29066
rect 9857 29008 9862 29064
rect 9918 29008 10058 29064
rect 9857 29006 10058 29008
rect 9857 29003 9923 29006
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 7465 28658 7531 28661
rect 7833 28658 7899 28661
rect 12525 28658 12591 28661
rect 7465 28656 12591 28658
rect 7465 28600 7470 28656
rect 7526 28600 7838 28656
rect 7894 28600 12530 28656
rect 12586 28600 12591 28656
rect 7465 28598 12591 28600
rect 7465 28595 7531 28598
rect 7833 28595 7899 28598
rect 12525 28595 12591 28598
rect 7741 28522 7807 28525
rect 13077 28522 13143 28525
rect 15009 28522 15075 28525
rect 7741 28520 15075 28522
rect 7741 28464 7746 28520
rect 7802 28464 13082 28520
rect 13138 28464 15014 28520
rect 15070 28464 15075 28520
rect 7741 28462 15075 28464
rect 7741 28459 7807 28462
rect 13077 28459 13143 28462
rect 15009 28459 15075 28462
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 6085 27570 6151 27573
rect 12249 27570 12315 27573
rect 12617 27570 12683 27573
rect 6085 27568 12683 27570
rect 6085 27512 6090 27568
rect 6146 27512 12254 27568
rect 12310 27512 12622 27568
rect 12678 27512 12683 27568
rect 6085 27510 12683 27512
rect 6085 27507 6151 27510
rect 12249 27507 12315 27510
rect 12617 27507 12683 27510
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 0 27026 480 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 480 26966
rect 1577 26963 1643 26966
rect 7281 26890 7347 26893
rect 12525 26890 12591 26893
rect 13169 26890 13235 26893
rect 7281 26888 13235 26890
rect 7281 26832 7286 26888
rect 7342 26832 12530 26888
rect 12586 26832 13174 26888
rect 13230 26832 13235 26888
rect 7281 26830 13235 26832
rect 7281 26827 7347 26830
rect 12525 26827 12591 26830
rect 13169 26827 13235 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 7373 26482 7439 26485
rect 12341 26482 12407 26485
rect 7373 26480 12407 26482
rect 7373 26424 7378 26480
rect 7434 26424 12346 26480
rect 12402 26424 12407 26480
rect 7373 26422 12407 26424
rect 7373 26419 7439 26422
rect 12341 26419 12407 26422
rect 8385 26210 8451 26213
rect 8518 26210 8524 26212
rect 8385 26208 8524 26210
rect 8385 26152 8390 26208
rect 8446 26152 8524 26208
rect 8385 26150 8524 26152
rect 8385 26147 8451 26150
rect 8518 26148 8524 26150
rect 8588 26148 8594 26212
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 8293 24850 8359 24853
rect 8477 24850 8543 24853
rect 9857 24850 9923 24853
rect 8293 24848 9923 24850
rect 8293 24792 8298 24848
rect 8354 24792 8482 24848
rect 8538 24792 9862 24848
rect 9918 24792 9923 24848
rect 8293 24790 9923 24792
rect 8293 24787 8359 24790
rect 8477 24787 8543 24790
rect 9857 24787 9923 24790
rect 7097 24714 7163 24717
rect 8385 24714 8451 24717
rect 7097 24712 8451 24714
rect 7097 24656 7102 24712
rect 7158 24656 8390 24712
rect 8446 24656 8451 24712
rect 7097 24654 8451 24656
rect 7097 24651 7163 24654
rect 8385 24651 8451 24654
rect 0 24578 480 24608
rect 2773 24578 2839 24581
rect 0 24576 2839 24578
rect 0 24520 2778 24576
rect 2834 24520 2839 24576
rect 0 24518 2839 24520
rect 0 24488 480 24518
rect 2773 24515 2839 24518
rect 7649 24578 7715 24581
rect 9673 24578 9739 24581
rect 7649 24576 9739 24578
rect 7649 24520 7654 24576
rect 7710 24520 9678 24576
rect 9734 24520 9739 24576
rect 7649 24518 9739 24520
rect 7649 24515 7715 24518
rect 9673 24515 9739 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 5073 24306 5139 24309
rect 9673 24306 9739 24309
rect 5073 24304 9739 24306
rect 5073 24248 5078 24304
rect 5134 24248 9678 24304
rect 9734 24248 9739 24304
rect 5073 24246 9739 24248
rect 5073 24243 5139 24246
rect 9673 24243 9739 24246
rect 2497 24170 2563 24173
rect 4797 24170 4863 24173
rect 2497 24168 4863 24170
rect 2497 24112 2502 24168
rect 2558 24112 4802 24168
rect 4858 24112 4863 24168
rect 2497 24110 4863 24112
rect 2497 24107 2563 24110
rect 4797 24107 4863 24110
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 2221 22674 2287 22677
rect 7833 22674 7899 22677
rect 2221 22672 7899 22674
rect 2221 22616 2226 22672
rect 2282 22616 7838 22672
rect 7894 22616 7899 22672
rect 2221 22614 7899 22616
rect 2221 22611 2287 22614
rect 7833 22611 7899 22614
rect 7741 22538 7807 22541
rect 12985 22538 13051 22541
rect 7741 22536 13051 22538
rect 7741 22480 7746 22536
rect 7802 22480 12990 22536
rect 13046 22480 13051 22536
rect 7741 22478 13051 22480
rect 7741 22475 7807 22478
rect 12985 22475 13051 22478
rect 6277 22336 6597 22337
rect 0 22266 480 22296
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 1669 22266 1735 22269
rect 0 22264 1735 22266
rect 0 22208 1674 22264
rect 1730 22208 1735 22264
rect 0 22206 1735 22208
rect 0 22176 480 22206
rect 1669 22203 1735 22206
rect 9673 22128 9739 22133
rect 9673 22072 9678 22128
rect 9734 22072 9739 22128
rect 9673 22067 9739 22072
rect 9676 21861 9736 22067
rect 9673 21856 9739 21861
rect 9673 21800 9678 21856
rect 9734 21800 9739 21856
rect 9673 21795 9739 21800
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 10501 21586 10567 21589
rect 12065 21586 12131 21589
rect 10501 21584 12131 21586
rect 10501 21528 10506 21584
rect 10562 21528 12070 21584
rect 12126 21528 12131 21584
rect 10501 21526 12131 21528
rect 10501 21523 10567 21526
rect 12065 21523 12131 21526
rect 5441 21450 5507 21453
rect 10041 21450 10107 21453
rect 5441 21448 10107 21450
rect 5441 21392 5446 21448
rect 5502 21392 10046 21448
rect 10102 21392 10107 21448
rect 5441 21390 10107 21392
rect 5441 21387 5507 21390
rect 10041 21387 10107 21390
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 8518 20980 8524 21044
rect 8588 21042 8594 21044
rect 8661 21042 8727 21045
rect 8588 21040 8727 21042
rect 8588 20984 8666 21040
rect 8722 20984 8727 21040
rect 8588 20982 8727 20984
rect 8588 20980 8594 20982
rect 8661 20979 8727 20982
rect 11329 21042 11395 21045
rect 12433 21042 12499 21045
rect 11329 21040 12499 21042
rect 11329 20984 11334 21040
rect 11390 20984 12438 21040
rect 12494 20984 12499 21040
rect 11329 20982 12499 20984
rect 11329 20979 11395 20982
rect 12433 20979 12499 20982
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 7557 20226 7623 20229
rect 10133 20226 10199 20229
rect 7557 20224 10199 20226
rect 7557 20168 7562 20224
rect 7618 20168 10138 20224
rect 10194 20168 10199 20224
rect 7557 20166 10199 20168
rect 7557 20163 7623 20166
rect 10133 20163 10199 20166
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 7281 20090 7347 20093
rect 8017 20090 8083 20093
rect 10133 20090 10199 20093
rect 7281 20088 10199 20090
rect 7281 20032 7286 20088
rect 7342 20032 8022 20088
rect 8078 20032 10138 20088
rect 10194 20032 10199 20088
rect 7281 20030 10199 20032
rect 7281 20027 7347 20030
rect 8017 20027 8083 20030
rect 10133 20027 10199 20030
rect 0 19954 480 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 480 19894
rect 1577 19891 1643 19894
rect 5165 19818 5231 19821
rect 6545 19818 6611 19821
rect 7281 19818 7347 19821
rect 10685 19818 10751 19821
rect 11053 19818 11119 19821
rect 5165 19816 11119 19818
rect 5165 19760 5170 19816
rect 5226 19760 6550 19816
rect 6606 19760 7286 19816
rect 7342 19760 10690 19816
rect 10746 19760 11058 19816
rect 11114 19760 11119 19816
rect 5165 19758 11119 19760
rect 5165 19755 5231 19758
rect 6545 19755 6611 19758
rect 7281 19755 7347 19758
rect 10685 19755 10751 19758
rect 11053 19755 11119 19758
rect 2773 19682 2839 19685
rect 3049 19682 3115 19685
rect 2773 19680 3115 19682
rect 2773 19624 2778 19680
rect 2834 19624 3054 19680
rect 3110 19624 3115 19680
rect 2773 19622 3115 19624
rect 2773 19619 2839 19622
rect 3049 19619 3115 19622
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 8109 19410 8175 19413
rect 9213 19410 9279 19413
rect 10869 19410 10935 19413
rect 8109 19408 10935 19410
rect 8109 19352 8114 19408
rect 8170 19352 9218 19408
rect 9274 19352 10874 19408
rect 10930 19352 10935 19408
rect 8109 19350 10935 19352
rect 8109 19347 8175 19350
rect 9213 19347 9279 19350
rect 10869 19347 10935 19350
rect 6913 19274 6979 19277
rect 10777 19274 10843 19277
rect 6913 19272 10843 19274
rect 6913 19216 6918 19272
rect 6974 19216 10782 19272
rect 10838 19216 10843 19272
rect 6913 19214 10843 19216
rect 6913 19211 6979 19214
rect 10777 19211 10843 19214
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 5073 18866 5139 18869
rect 9857 18866 9923 18869
rect 13537 18866 13603 18869
rect 5073 18864 13603 18866
rect 5073 18808 5078 18864
rect 5134 18808 9862 18864
rect 9918 18808 13542 18864
rect 13598 18808 13603 18864
rect 5073 18806 13603 18808
rect 5073 18803 5139 18806
rect 9857 18803 9923 18806
rect 13537 18803 13603 18806
rect 6821 18730 6887 18733
rect 7557 18730 7623 18733
rect 6821 18728 7623 18730
rect 6821 18672 6826 18728
rect 6882 18672 7562 18728
rect 7618 18672 7623 18728
rect 6821 18670 7623 18672
rect 6821 18667 6887 18670
rect 7557 18667 7623 18670
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 3693 18186 3759 18189
rect 3693 18184 7666 18186
rect 3693 18128 3698 18184
rect 3754 18128 7666 18184
rect 3693 18126 7666 18128
rect 3693 18123 3759 18126
rect 7606 18050 7666 18126
rect 8753 18050 8819 18053
rect 10041 18050 10107 18053
rect 7606 18048 10107 18050
rect 7606 17992 8758 18048
rect 8814 17992 10046 18048
rect 10102 17992 10107 18048
rect 7606 17990 10107 17992
rect 8753 17987 8819 17990
rect 10041 17987 10107 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 10593 17778 10659 17781
rect 13169 17778 13235 17781
rect 10593 17776 13235 17778
rect 10593 17720 10598 17776
rect 10654 17720 13174 17776
rect 13230 17720 13235 17776
rect 10593 17718 13235 17720
rect 10593 17715 10659 17718
rect 13169 17715 13235 17718
rect 0 17642 480 17672
rect 1669 17642 1735 17645
rect 0 17640 1735 17642
rect 0 17584 1674 17640
rect 1730 17584 1735 17640
rect 0 17582 1735 17584
rect 0 17552 480 17582
rect 1669 17579 1735 17582
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 3969 17234 4035 17237
rect 7005 17234 7071 17237
rect 8109 17234 8175 17237
rect 3969 17232 8175 17234
rect 3969 17176 3974 17232
rect 4030 17176 7010 17232
rect 7066 17176 8114 17232
rect 8170 17176 8175 17232
rect 3969 17174 8175 17176
rect 3969 17171 4035 17174
rect 7005 17171 7071 17174
rect 8109 17171 8175 17174
rect 3969 17098 4035 17101
rect 9489 17098 9555 17101
rect 3969 17096 9555 17098
rect 3969 17040 3974 17096
rect 4030 17040 9494 17096
rect 9550 17040 9555 17096
rect 3969 17038 9555 17040
rect 3969 17035 4035 17038
rect 9489 17035 9555 17038
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 1393 16690 1459 16693
rect 7373 16690 7439 16693
rect 1393 16688 7439 16690
rect 1393 16632 1398 16688
rect 1454 16632 7378 16688
rect 7434 16632 7439 16688
rect 1393 16630 7439 16632
rect 1393 16627 1459 16630
rect 7373 16627 7439 16630
rect 8017 16690 8083 16693
rect 9673 16690 9739 16693
rect 8017 16688 9739 16690
rect 8017 16632 8022 16688
rect 8078 16632 9678 16688
rect 9734 16632 9739 16688
rect 8017 16630 9739 16632
rect 8017 16627 8083 16630
rect 9673 16627 9739 16630
rect 10501 16690 10567 16693
rect 12525 16690 12591 16693
rect 10501 16688 12591 16690
rect 10501 16632 10506 16688
rect 10562 16632 12530 16688
rect 12586 16632 12591 16688
rect 10501 16630 12591 16632
rect 10501 16627 10567 16630
rect 12525 16627 12591 16630
rect 3325 16554 3391 16557
rect 8661 16554 8727 16557
rect 3325 16552 8727 16554
rect 3325 16496 3330 16552
rect 3386 16496 8666 16552
rect 8722 16496 8727 16552
rect 3325 16494 8727 16496
rect 3325 16491 3391 16494
rect 8661 16491 8727 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 9857 16146 9923 16149
rect 10685 16146 10751 16149
rect 12433 16146 12499 16149
rect 9857 16144 12499 16146
rect 9857 16088 9862 16144
rect 9918 16088 10690 16144
rect 10746 16088 12438 16144
rect 12494 16088 12499 16144
rect 9857 16086 12499 16088
rect 9857 16083 9923 16086
rect 10685 16083 10751 16086
rect 12433 16083 12499 16086
rect 3785 15874 3851 15877
rect 5073 15874 5139 15877
rect 3785 15872 5139 15874
rect 3785 15816 3790 15872
rect 3846 15816 5078 15872
rect 5134 15816 5139 15872
rect 3785 15814 5139 15816
rect 3785 15811 3851 15814
rect 5073 15811 5139 15814
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 9622 15268 9628 15332
rect 9692 15330 9698 15332
rect 12709 15330 12775 15333
rect 9692 15328 12775 15330
rect 9692 15272 12714 15328
rect 12770 15272 12775 15328
rect 9692 15270 12775 15272
rect 9692 15268 9698 15270
rect 12709 15267 12775 15270
rect 3610 15264 3930 15265
rect 0 15194 480 15224
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 480 15134
rect 1669 15131 1735 15134
rect 9213 15058 9279 15061
rect 9622 15058 9628 15060
rect 9213 15056 9628 15058
rect 9213 15000 9218 15056
rect 9274 15000 9628 15056
rect 9213 14998 9628 15000
rect 9213 14995 9279 14998
rect 9622 14996 9628 14998
rect 9692 14996 9698 15060
rect 3785 14786 3851 14789
rect 5533 14786 5599 14789
rect 3785 14784 5599 14786
rect 3785 14728 3790 14784
rect 3846 14728 5538 14784
rect 5594 14728 5599 14784
rect 3785 14726 5599 14728
rect 3785 14723 3851 14726
rect 5533 14723 5599 14726
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 1669 13970 1735 13973
rect 10133 13970 10199 13973
rect 1669 13968 10199 13970
rect 1669 13912 1674 13968
rect 1730 13912 10138 13968
rect 10194 13912 10199 13968
rect 1669 13910 10199 13912
rect 1669 13907 1735 13910
rect 10133 13907 10199 13910
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 0 12882 480 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 480 12822
rect 1577 12819 1643 12822
rect 5073 12746 5139 12749
rect 7097 12746 7163 12749
rect 11421 12746 11487 12749
rect 5073 12744 11487 12746
rect 5073 12688 5078 12744
rect 5134 12688 7102 12744
rect 7158 12688 11426 12744
rect 11482 12688 11487 12744
rect 5073 12686 11487 12688
rect 5073 12683 5139 12686
rect 7097 12683 7163 12686
rect 11421 12683 11487 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 4889 12338 4955 12341
rect 8385 12338 8451 12341
rect 9949 12338 10015 12341
rect 4889 12336 10015 12338
rect 4889 12280 4894 12336
rect 4950 12280 8390 12336
rect 8446 12280 9954 12336
rect 10010 12280 10015 12336
rect 4889 12278 10015 12280
rect 4889 12275 4955 12278
rect 8385 12275 8451 12278
rect 9949 12275 10015 12278
rect 10869 12338 10935 12341
rect 12433 12338 12499 12341
rect 10869 12336 12499 12338
rect 10869 12280 10874 12336
rect 10930 12280 12438 12336
rect 12494 12280 12499 12336
rect 10869 12278 12499 12280
rect 10869 12275 10935 12278
rect 12433 12275 12499 12278
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 7005 11794 7071 11797
rect 12157 11794 12223 11797
rect 7005 11792 12223 11794
rect 7005 11736 7010 11792
rect 7066 11736 12162 11792
rect 12218 11736 12223 11792
rect 7005 11734 12223 11736
rect 7005 11731 7071 11734
rect 12157 11731 12223 11734
rect 2221 11658 2287 11661
rect 7741 11658 7807 11661
rect 2221 11656 7807 11658
rect 2221 11600 2226 11656
rect 2282 11600 7746 11656
rect 7802 11600 7807 11656
rect 2221 11598 7807 11600
rect 2221 11595 2287 11598
rect 7741 11595 7807 11598
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 7925 11386 7991 11389
rect 9581 11386 9647 11389
rect 7925 11384 9647 11386
rect 7925 11328 7930 11384
rect 7986 11328 9586 11384
rect 9642 11328 9647 11384
rect 7925 11326 9647 11328
rect 7925 11323 7991 11326
rect 9581 11323 9647 11326
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 11973 10706 12039 10709
rect 14181 10706 14247 10709
rect 11973 10704 14247 10706
rect 11973 10648 11978 10704
rect 12034 10648 14186 10704
rect 14242 10648 14247 10704
rect 11973 10646 14247 10648
rect 11973 10643 12039 10646
rect 14181 10643 14247 10646
rect 0 10570 480 10600
rect 1669 10570 1735 10573
rect 0 10568 1735 10570
rect 0 10512 1674 10568
rect 1730 10512 1735 10568
rect 0 10510 1735 10512
rect 0 10480 480 10510
rect 1669 10507 1735 10510
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 6085 10026 6151 10029
rect 15520 10026 16000 10056
rect 6085 10024 16000 10026
rect 6085 9968 6090 10024
rect 6146 9968 16000 10024
rect 6085 9966 16000 9968
rect 6085 9963 6151 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 4889 9754 4955 9757
rect 4889 9752 8402 9754
rect 4889 9696 4894 9752
rect 4950 9696 8402 9752
rect 4889 9694 8402 9696
rect 4889 9691 4955 9694
rect 4429 9618 4495 9621
rect 7005 9618 7071 9621
rect 4429 9616 7071 9618
rect 4429 9560 4434 9616
rect 4490 9560 7010 9616
rect 7066 9560 7071 9616
rect 4429 9558 7071 9560
rect 8342 9618 8402 9694
rect 9806 9618 9812 9620
rect 8342 9558 9812 9618
rect 4429 9555 4495 9558
rect 7005 9555 7071 9558
rect 9806 9556 9812 9558
rect 9876 9556 9882 9620
rect 10133 9482 10199 9485
rect 13537 9482 13603 9485
rect 10133 9480 13603 9482
rect 10133 9424 10138 9480
rect 10194 9424 13542 9480
rect 13598 9424 13603 9480
rect 10133 9422 13603 9424
rect 10133 9419 10199 9422
rect 13537 9419 13603 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 7281 8938 7347 8941
rect 8753 8938 8819 8941
rect 10409 8938 10475 8941
rect 7281 8936 10475 8938
rect 7281 8880 7286 8936
rect 7342 8880 8758 8936
rect 8814 8880 10414 8936
rect 10470 8880 10475 8936
rect 7281 8878 10475 8880
rect 7281 8875 7347 8878
rect 8753 8875 8819 8878
rect 10409 8875 10475 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 2865 8394 2931 8397
rect 4705 8394 4771 8397
rect 2865 8392 4771 8394
rect 2865 8336 2870 8392
rect 2926 8336 4710 8392
rect 4766 8336 4771 8392
rect 2865 8334 4771 8336
rect 2865 8331 2931 8334
rect 4705 8331 4771 8334
rect 6729 8394 6795 8397
rect 9029 8394 9095 8397
rect 6729 8392 9095 8394
rect 6729 8336 6734 8392
rect 6790 8336 9034 8392
rect 9090 8336 9095 8392
rect 6729 8334 9095 8336
rect 6729 8331 6795 8334
rect 9029 8331 9095 8334
rect 6277 8192 6597 8193
rect 0 8122 480 8152
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 480 8062
rect 1485 8059 1551 8062
rect 2405 7986 2471 7989
rect 9949 7986 10015 7989
rect 2405 7984 10015 7986
rect 2405 7928 2410 7984
rect 2466 7928 9954 7984
rect 10010 7928 10015 7984
rect 2405 7926 10015 7928
rect 2405 7923 2471 7926
rect 9949 7923 10015 7926
rect 5073 7850 5139 7853
rect 9673 7852 9739 7853
rect 9622 7850 9628 7852
rect 5073 7848 9628 7850
rect 9692 7850 9739 7852
rect 9692 7848 9820 7850
rect 5073 7792 5078 7848
rect 5134 7792 9628 7848
rect 9734 7792 9820 7848
rect 5073 7790 9628 7792
rect 5073 7787 5139 7790
rect 9622 7788 9628 7790
rect 9692 7790 9820 7792
rect 9692 7788 9739 7790
rect 9673 7787 9739 7788
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 5349 7306 5415 7309
rect 7005 7306 7071 7309
rect 5349 7304 7071 7306
rect 5349 7248 5354 7304
rect 5410 7248 7010 7304
rect 7066 7248 7071 7304
rect 5349 7246 7071 7248
rect 5349 7243 5415 7246
rect 7005 7243 7071 7246
rect 8937 7306 9003 7309
rect 10869 7306 10935 7309
rect 8937 7304 10935 7306
rect 8937 7248 8942 7304
rect 8998 7248 10874 7304
rect 10930 7248 10935 7304
rect 8937 7246 10935 7248
rect 8937 7243 9003 7246
rect 10869 7243 10935 7246
rect 7833 7170 7899 7173
rect 8385 7170 8451 7173
rect 11145 7170 11211 7173
rect 7833 7168 11211 7170
rect 7833 7112 7838 7168
rect 7894 7112 8390 7168
rect 8446 7112 11150 7168
rect 11206 7112 11211 7168
rect 7833 7110 11211 7112
rect 7833 7107 7899 7110
rect 8385 7107 8451 7110
rect 11145 7107 11211 7110
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 6729 7034 6795 7037
rect 11237 7034 11303 7037
rect 6729 7032 11303 7034
rect 6729 6976 6734 7032
rect 6790 6976 11242 7032
rect 11298 6976 11303 7032
rect 6729 6974 11303 6976
rect 6729 6971 6795 6974
rect 11237 6971 11303 6974
rect 7373 6898 7439 6901
rect 8661 6898 8727 6901
rect 7373 6896 8727 6898
rect 7373 6840 7378 6896
rect 7434 6840 8666 6896
rect 8722 6840 8727 6896
rect 7373 6838 8727 6840
rect 7373 6835 7439 6838
rect 8661 6835 8727 6838
rect 6821 6762 6887 6765
rect 8661 6762 8727 6765
rect 6821 6760 8727 6762
rect 6821 6704 6826 6760
rect 6882 6704 8666 6760
rect 8722 6704 8727 6760
rect 6821 6702 8727 6704
rect 6821 6699 6887 6702
rect 8661 6699 8727 6702
rect 8937 6762 9003 6765
rect 9397 6762 9463 6765
rect 10685 6762 10751 6765
rect 8937 6760 10751 6762
rect 8937 6704 8942 6760
rect 8998 6704 9402 6760
rect 9458 6704 10690 6760
rect 10746 6704 10751 6760
rect 8937 6702 10751 6704
rect 8937 6699 9003 6702
rect 9397 6699 9463 6702
rect 10685 6699 10751 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 5625 6490 5691 6493
rect 5993 6490 6059 6493
rect 5625 6488 8080 6490
rect 5625 6432 5630 6488
rect 5686 6432 5998 6488
rect 6054 6432 8080 6488
rect 5625 6430 8080 6432
rect 5625 6427 5691 6430
rect 5993 6427 6059 6430
rect 2405 6354 2471 6357
rect 5993 6354 6059 6357
rect 2405 6352 6059 6354
rect 2405 6296 2410 6352
rect 2466 6296 5998 6352
rect 6054 6296 6059 6352
rect 2405 6294 6059 6296
rect 2405 6291 2471 6294
rect 5993 6291 6059 6294
rect 3233 6218 3299 6221
rect 7833 6218 7899 6221
rect 3233 6216 7899 6218
rect 3233 6160 3238 6216
rect 3294 6160 7838 6216
rect 7894 6160 7899 6216
rect 3233 6158 7899 6160
rect 8020 6218 8080 6430
rect 8201 6354 8267 6357
rect 10501 6354 10567 6357
rect 11053 6354 11119 6357
rect 8201 6352 11119 6354
rect 8201 6296 8206 6352
rect 8262 6296 10506 6352
rect 10562 6296 11058 6352
rect 11114 6296 11119 6352
rect 8201 6294 11119 6296
rect 8201 6291 8267 6294
rect 10501 6291 10567 6294
rect 11053 6291 11119 6294
rect 10225 6218 10291 6221
rect 8020 6216 10291 6218
rect 8020 6160 10230 6216
rect 10286 6160 10291 6216
rect 8020 6158 10291 6160
rect 3233 6155 3299 6158
rect 7833 6155 7899 6158
rect 10225 6155 10291 6158
rect 7465 6082 7531 6085
rect 10869 6082 10935 6085
rect 7465 6080 10935 6082
rect 7465 6024 7470 6080
rect 7526 6024 10874 6080
rect 10930 6024 10935 6080
rect 7465 6022 10935 6024
rect 7465 6019 7531 6022
rect 10869 6019 10935 6022
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 0 5810 480 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 480 5750
rect 1577 5747 1643 5750
rect 6821 5810 6887 5813
rect 9673 5810 9739 5813
rect 6821 5808 9739 5810
rect 6821 5752 6826 5808
rect 6882 5752 9678 5808
rect 9734 5752 9739 5808
rect 6821 5750 9739 5752
rect 6821 5747 6887 5750
rect 9673 5747 9739 5750
rect 7833 5674 7899 5677
rect 10041 5674 10107 5677
rect 7833 5672 10107 5674
rect 7833 5616 7838 5672
rect 7894 5616 10046 5672
rect 10102 5616 10107 5672
rect 7833 5614 10107 5616
rect 7833 5611 7899 5614
rect 10041 5611 10107 5614
rect 13445 5674 13511 5677
rect 15745 5674 15811 5677
rect 13445 5672 15811 5674
rect 13445 5616 13450 5672
rect 13506 5616 15750 5672
rect 15806 5616 15811 5672
rect 13445 5614 15811 5616
rect 13445 5611 13511 5614
rect 15745 5611 15811 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 9397 5402 9463 5405
rect 11237 5402 11303 5405
rect 9397 5400 11303 5402
rect 9397 5344 9402 5400
rect 9458 5344 11242 5400
rect 11298 5344 11303 5400
rect 9397 5342 11303 5344
rect 9397 5339 9463 5342
rect 11237 5339 11303 5342
rect 5901 5266 5967 5269
rect 10317 5266 10383 5269
rect 5901 5264 10383 5266
rect 5901 5208 5906 5264
rect 5962 5208 10322 5264
rect 10378 5208 10383 5264
rect 5901 5206 10383 5208
rect 5901 5203 5967 5206
rect 10317 5203 10383 5206
rect 5533 5130 5599 5133
rect 14641 5130 14707 5133
rect 5533 5128 14707 5130
rect 5533 5072 5538 5128
rect 5594 5072 14646 5128
rect 14702 5072 14707 5128
rect 5533 5070 14707 5072
rect 5533 5067 5599 5070
rect 14641 5067 14707 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 5717 4858 5783 4861
rect 5717 4856 5826 4858
rect 5717 4800 5722 4856
rect 5778 4800 5826 4856
rect 5717 4795 5826 4800
rect 5766 4722 5826 4795
rect 10501 4722 10567 4725
rect 13353 4722 13419 4725
rect 5766 4720 13419 4722
rect 5766 4664 10506 4720
rect 10562 4664 13358 4720
rect 13414 4664 13419 4720
rect 5766 4662 13419 4664
rect 10501 4659 10567 4662
rect 13353 4659 13419 4662
rect 2773 4586 2839 4589
rect 7097 4586 7163 4589
rect 12617 4586 12683 4589
rect 2773 4584 6930 4586
rect 2773 4528 2778 4584
rect 2834 4528 6930 4584
rect 2773 4526 6930 4528
rect 2773 4523 2839 4526
rect 6870 4450 6930 4526
rect 7097 4584 12683 4586
rect 7097 4528 7102 4584
rect 7158 4528 12622 4584
rect 12678 4528 12683 4584
rect 7097 4526 12683 4528
rect 7097 4523 7163 4526
rect 12617 4523 12683 4526
rect 8017 4450 8083 4453
rect 8201 4450 8267 4453
rect 6870 4448 8267 4450
rect 6870 4392 8022 4448
rect 8078 4392 8206 4448
rect 8262 4392 8267 4448
rect 6870 4390 8267 4392
rect 8017 4387 8083 4390
rect 8201 4387 8267 4390
rect 10041 4450 10107 4453
rect 12433 4450 12499 4453
rect 10041 4448 12499 4450
rect 10041 4392 10046 4448
rect 10102 4392 12438 4448
rect 12494 4392 12499 4448
rect 10041 4390 12499 4392
rect 10041 4387 10107 4390
rect 12433 4387 12499 4390
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 4521 4314 4587 4317
rect 8753 4314 8819 4317
rect 4521 4312 8819 4314
rect 4521 4256 4526 4312
rect 4582 4256 8758 4312
rect 8814 4256 8819 4312
rect 4521 4254 8819 4256
rect 4521 4251 4587 4254
rect 8753 4251 8819 4254
rect 1485 4178 1551 4181
rect 4245 4178 4311 4181
rect 1485 4176 4311 4178
rect 1485 4120 1490 4176
rect 1546 4120 4250 4176
rect 4306 4120 4311 4176
rect 1485 4118 4311 4120
rect 1485 4115 1551 4118
rect 4245 4115 4311 4118
rect 4981 4178 5047 4181
rect 8477 4178 8543 4181
rect 4981 4176 8543 4178
rect 4981 4120 4986 4176
rect 5042 4120 8482 4176
rect 8538 4120 8543 4176
rect 4981 4118 8543 4120
rect 4981 4115 5047 4118
rect 8477 4115 8543 4118
rect 3877 4042 3943 4045
rect 4797 4042 4863 4045
rect 9029 4042 9095 4045
rect 12617 4042 12683 4045
rect 3877 4040 9095 4042
rect 3877 3984 3882 4040
rect 3938 3984 4802 4040
rect 4858 3984 9034 4040
rect 9090 3984 9095 4040
rect 3877 3982 9095 3984
rect 3877 3979 3943 3982
rect 4797 3979 4863 3982
rect 9029 3979 9095 3982
rect 9262 4040 12683 4042
rect 9262 3984 12622 4040
rect 12678 3984 12683 4040
rect 9262 3982 12683 3984
rect 4337 3906 4403 3909
rect 6085 3906 6151 3909
rect 4337 3904 6151 3906
rect 4337 3848 4342 3904
rect 4398 3848 6090 3904
rect 6146 3848 6151 3904
rect 4337 3846 6151 3848
rect 4337 3843 4403 3846
rect 6085 3843 6151 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 3325 3770 3391 3773
rect 6085 3770 6151 3773
rect 3325 3768 6151 3770
rect 3325 3712 3330 3768
rect 3386 3712 6090 3768
rect 6146 3712 6151 3768
rect 3325 3710 6151 3712
rect 3325 3707 3391 3710
rect 6085 3707 6151 3710
rect 6177 3634 6243 3637
rect 9262 3634 9322 3982
rect 12617 3979 12683 3982
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 6177 3632 9322 3634
rect 6177 3576 6182 3632
rect 6238 3576 9322 3632
rect 6177 3574 9322 3576
rect 10593 3634 10659 3637
rect 12617 3634 12683 3637
rect 10593 3632 12683 3634
rect 10593 3576 10598 3632
rect 10654 3576 12622 3632
rect 12678 3576 12683 3632
rect 10593 3574 12683 3576
rect 6177 3571 6243 3574
rect 10593 3571 10659 3574
rect 12617 3571 12683 3574
rect 13077 3634 13143 3637
rect 15377 3634 15443 3637
rect 13077 3632 15443 3634
rect 13077 3576 13082 3632
rect 13138 3576 15382 3632
rect 15438 3576 15443 3632
rect 13077 3574 15443 3576
rect 13077 3571 13143 3574
rect 15377 3571 15443 3574
rect 0 3498 480 3528
rect 1669 3498 1735 3501
rect 0 3496 1735 3498
rect 0 3440 1674 3496
rect 1730 3440 1735 3496
rect 0 3438 1735 3440
rect 0 3408 480 3438
rect 1669 3435 1735 3438
rect 4705 3498 4771 3501
rect 7741 3498 7807 3501
rect 10777 3498 10843 3501
rect 4705 3496 10843 3498
rect 4705 3440 4710 3496
rect 4766 3440 7746 3496
rect 7802 3440 10782 3496
rect 10838 3440 10843 3496
rect 4705 3438 10843 3440
rect 4705 3435 4771 3438
rect 7741 3435 7807 3438
rect 10777 3435 10843 3438
rect 9397 3362 9463 3365
rect 12709 3362 12775 3365
rect 9397 3360 12775 3362
rect 9397 3304 9402 3360
rect 9458 3304 12714 3360
rect 12770 3304 12775 3360
rect 9397 3302 12775 3304
rect 9397 3299 9463 3302
rect 12709 3299 12775 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 6637 3226 6703 3229
rect 8569 3226 8635 3229
rect 6637 3224 8635 3226
rect 6637 3168 6642 3224
rect 6698 3168 8574 3224
rect 8630 3168 8635 3224
rect 6637 3166 8635 3168
rect 6637 3163 6703 3166
rect 8569 3163 8635 3166
rect 7741 3090 7807 3093
rect 12801 3090 12867 3093
rect 7741 3088 12867 3090
rect 7741 3032 7746 3088
rect 7802 3032 12806 3088
rect 12862 3032 12867 3088
rect 7741 3030 12867 3032
rect 7741 3027 7807 3030
rect 12801 3027 12867 3030
rect 4153 2954 4219 2957
rect 10133 2954 10199 2957
rect 4153 2952 10199 2954
rect 4153 2896 4158 2952
rect 4214 2896 10138 2952
rect 10194 2896 10199 2952
rect 4153 2894 10199 2896
rect 4153 2891 4219 2894
rect 10133 2891 10199 2894
rect 10961 2954 11027 2957
rect 12341 2954 12407 2957
rect 10961 2952 12407 2954
rect 10961 2896 10966 2952
rect 11022 2896 12346 2952
rect 12402 2896 12407 2952
rect 10961 2894 12407 2896
rect 10961 2891 11027 2894
rect 12341 2891 12407 2894
rect 9397 2818 9463 2821
rect 11421 2818 11487 2821
rect 12065 2818 12131 2821
rect 9397 2816 11487 2818
rect 9397 2760 9402 2816
rect 9458 2760 11426 2816
rect 11482 2760 11487 2816
rect 9397 2758 11487 2760
rect 9397 2755 9463 2758
rect 11421 2755 11487 2758
rect 12022 2816 12131 2818
rect 12022 2760 12070 2816
rect 12126 2760 12131 2816
rect 12022 2755 12131 2760
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 9622 2620 9628 2684
rect 9692 2682 9698 2684
rect 9765 2682 9831 2685
rect 9692 2680 9831 2682
rect 9692 2624 9770 2680
rect 9826 2624 9831 2680
rect 9692 2622 9831 2624
rect 9692 2620 9698 2622
rect 9765 2619 9831 2622
rect 8017 2546 8083 2549
rect 11881 2546 11947 2549
rect 12022 2546 12082 2755
rect 8017 2544 12082 2546
rect 8017 2488 8022 2544
rect 8078 2488 11886 2544
rect 11942 2488 12082 2544
rect 8017 2486 12082 2488
rect 8017 2483 8083 2486
rect 11881 2483 11947 2486
rect 6269 2410 6335 2413
rect 13629 2410 13695 2413
rect 6269 2408 13695 2410
rect 6269 2352 6274 2408
rect 6330 2352 13634 2408
rect 13690 2352 13695 2408
rect 6269 2350 13695 2352
rect 6269 2347 6335 2350
rect 13629 2347 13695 2350
rect 9806 2212 9812 2276
rect 9876 2274 9882 2276
rect 9949 2274 10015 2277
rect 9876 2272 10015 2274
rect 9876 2216 9954 2272
rect 10010 2216 10015 2272
rect 9876 2214 10015 2216
rect 9876 2212 9882 2214
rect 9949 2211 10015 2214
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 8661 2002 8727 2005
rect 13721 2002 13787 2005
rect 8661 2000 13787 2002
rect 8661 1944 8666 2000
rect 8722 1944 13726 2000
rect 13782 1944 13787 2000
rect 8661 1942 13787 1944
rect 8661 1939 8727 1942
rect 13721 1939 13787 1942
rect 3325 1730 3391 1733
rect 8753 1730 8819 1733
rect 3325 1728 8819 1730
rect 3325 1672 3330 1728
rect 3386 1672 8758 1728
rect 8814 1672 8819 1728
rect 3325 1670 8819 1672
rect 3325 1667 3391 1670
rect 8753 1667 8819 1670
rect 2957 1594 3023 1597
rect 7649 1594 7715 1597
rect 2957 1592 7715 1594
rect 2957 1536 2962 1592
rect 3018 1536 7654 1592
rect 7710 1536 7715 1592
rect 2957 1534 7715 1536
rect 2957 1531 3023 1534
rect 7649 1531 7715 1534
rect 1393 1458 1459 1461
rect 1350 1456 1459 1458
rect 1350 1400 1398 1456
rect 1454 1400 1459 1456
rect 1350 1395 1459 1400
rect 3785 1458 3851 1461
rect 5809 1458 5875 1461
rect 3785 1456 5875 1458
rect 3785 1400 3790 1456
rect 3846 1400 5814 1456
rect 5870 1400 5875 1456
rect 3785 1398 5875 1400
rect 3785 1395 3851 1398
rect 5809 1395 5875 1398
rect 0 1186 480 1216
rect 1350 1186 1410 1395
rect 0 1126 1410 1186
rect 0 1096 480 1126
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 7604 35396 7668 35460
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 9628 33764 9692 33828
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 7604 29472 7668 29476
rect 7604 29416 7654 29472
rect 7654 29416 7668 29472
rect 7604 29412 7668 29416
rect 9628 29472 9692 29476
rect 9628 29416 9678 29472
rect 9678 29416 9692 29472
rect 9628 29412 9692 29416
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 8524 26148 8588 26212
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 8524 20980 8588 21044
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 9628 15268 9692 15332
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 9628 14996 9692 15060
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 9812 9556 9876 9620
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 9628 7848 9692 7852
rect 9628 7792 9678 7848
rect 9678 7792 9692 7848
rect 9628 7788 9692 7792
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 9628 2620 9692 2684
rect 9812 2212 9876 2276
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 7603 35460 7669 35461
rect 7603 35396 7604 35460
rect 7668 35396 7669 35460
rect 7603 35395 7669 35396
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 7606 29477 7666 35395
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 9627 33828 9693 33829
rect 9627 33764 9628 33828
rect 9692 33764 9693 33828
rect 9627 33763 9693 33764
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 7603 29476 7669 29477
rect 7603 29412 7604 29476
rect 7668 29412 7669 29476
rect 7603 29411 7669 29412
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 8944 29408 9264 30432
rect 9630 29477 9690 33763
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 9627 29476 9693 29477
rect 9627 29412 9628 29476
rect 9692 29412 9693 29476
rect 9627 29411 9693 29412
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8523 26212 8589 26213
rect 8523 26148 8524 26212
rect 8588 26148 8589 26212
rect 8523 26147 8589 26148
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 8526 21045 8586 26147
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8523 21044 8589 21045
rect 8523 20980 8524 21044
rect 8588 20980 8589 21044
rect 8523 20979 8589 20980
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 9627 15332 9693 15333
rect 9627 15268 9628 15332
rect 9692 15268 9693 15332
rect 9627 15267 9693 15268
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 9630 15061 9690 15267
rect 9627 15060 9693 15061
rect 9627 14996 9628 15060
rect 9692 14996 9693 15060
rect 9627 14995 9693 14996
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 9811 9620 9877 9621
rect 9811 9556 9812 9620
rect 9876 9556 9877 9620
rect 9811 9555 9877 9556
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 9630 2685 9690 7787
rect 9627 2684 9693 2685
rect 9627 2620 9628 2684
rect 9692 2620 9693 2684
rect 9627 2619 9693 2620
rect 9814 2277 9874 9555
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 9811 2276 9877 2277
rect 9811 2212 9812 2276
rect 9876 2212 9877 2276
rect 9811 2211 9877 2212
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_11
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1472 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_24
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1604681595
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1604681595
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1604681595
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73
timestamp 1604681595
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1604681595
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1604681595
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_112
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_108
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_75
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1604681595
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_83
timestamp 1604681595
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_87
timestamp 1604681595
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1604681595
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13524 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_127
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_138
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_48
timestamp 1604681595
transform 1 0 5520 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_52
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_55
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1604681595
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1604681595
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_116
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_131 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1604681595
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1604681595
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_49
timestamp 1604681595
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1604681595
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_87
timestamp 1604681595
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_18
timestamp 1604681595
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 3496 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_22
timestamp 1604681595
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_45
timestamp 1604681595
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_49
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6992 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_80
timestamp 1604681595
transform 1 0 8464 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_89
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1604681595
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1604681595
transform 1 0 10948 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1604681595
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_117
timestamp 1604681595
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1604681595
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1604681595
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_13
timestamp 1604681595
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_16
timestamp 1604681595
transform 1 0 2576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 2668 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1604681595
transform 1 0 3404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_25
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1604681595
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_40
timestamp 1604681595
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp 1604681595
transform 1 0 5520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_44
timestamp 1604681595
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1604681595
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_77
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 8280 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1604681595
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_6_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_95
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1604681595
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 10212 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1604681595
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 13248 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_140
timestamp 1604681595
transform 1 0 13984 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_136
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_24
timestamp 1604681595
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1604681595
transform 1 0 4508 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4600 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_47
timestamp 1604681595
transform 1 0 5428 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1604681595
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_112
timestamp 1604681595
transform 1 0 11408 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_50
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_54
timestamp 1604681595
transform 1 0 6072 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1604681595
transform 1 0 1932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp 1604681595
transform 1 0 2300 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_16
timestamp 1604681595
transform 1 0 2576 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_22
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1604681595
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1604681595
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_102
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1604681595
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_122
timestamp 1604681595
transform 1 0 12328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_134
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_33
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 1604681595
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1604681595
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1604681595
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_95
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4324 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 5888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1604681595
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1604681595
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1604681595
transform 1 0 10120 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_110
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_122
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_134
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1604681595
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_36
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1604681595
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_40
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_52
timestamp 1604681595
transform 1 0 5888 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604681595
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 6624 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1604681595
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_103
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1604681595
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_118
timestamp 1604681595
transform 1 0 11960 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_130
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4508 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_29
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_33
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_54
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_58
timestamp 1604681595
transform 1 0 6440 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_81
timestamp 1604681595
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1604681595
transform 1 0 8924 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1604681595
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_112
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_143
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 4784 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1604681595
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_116
timestamp 1604681595
transform 1 0 11776 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_122
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_13
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_21
timestamp 1604681595
transform 1 0 3036 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_67
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_94
timestamp 1604681595
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_111
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_115
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_43
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_55
timestamp 1604681595
transform 1 0 6164 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_67
timestamp 1604681595
transform 1 0 7268 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_96
timestamp 1604681595
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_100
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_128
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_140
timestamp 1604681595
transform 1 0 13984 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_70
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_72
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_76
timestamp 1604681595
transform 1 0 8096 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_82
timestamp 1604681595
transform 1 0 8648 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1604681595
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1604681595
transform 1 0 9660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_100
timestamp 1604681595
transform 1 0 10304 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_100
timestamp 1604681595
transform 1 0 10304 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_108
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_116
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_137
timestamp 1604681595
transform 1 0 13708 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1604681595
transform 1 0 2852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1604681595
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_49
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_43
timestamp 1604681595
transform 1 0 5060 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1604681595
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_100
timestamp 1604681595
transform 1 0 10304 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_112
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_144
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_9
timestamp 1604681595
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_21
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5888 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11684 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1604681595
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1604681595
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1604681595
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_143
timestamp 1604681595
transform 1 0 14260 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_79
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1604681595
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1604681595
transform 1 0 5796 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_62
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_67
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11592 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_133
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_19
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_23
timestamp 1604681595
transform 1 0 3220 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp 1604681595
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7084 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9568 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_84
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_88
timestamp 1604681595
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_111
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1604681595
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_9
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1604681595
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1604681595
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1604681595
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_36
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_41
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_50
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_46
timestamp 1604681595
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_58
timestamp 1604681595
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_48
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1604681595
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1604681595
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1604681595
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_101
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11040 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_127
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_139
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1604681595
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_55
timestamp 1604681595
transform 1 0 6164 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_61
timestamp 1604681595
transform 1 0 6716 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_114
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_126
timestamp 1604681595
transform 1 0 12696 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_77
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 9108 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp 1604681595
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_90
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1604681595
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_19
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_22
timestamp 1604681595
transform 1 0 3128 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1604681595
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1604681595
transform 1 0 6072 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1604681595
transform 1 0 6716 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1604681595
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_110
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_122
timestamp 1604681595
transform 1 0 12328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_134
timestamp 1604681595
transform 1 0 13432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2944 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_29
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_81
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9292 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_108
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_112
timestamp 1604681595
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_116
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_143
timestamp 1604681595
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1604681595
transform 1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_13
timestamp 1604681595
transform 1 0 2300 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1604681595
transform 1 0 2576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4324 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_26
timestamp 1604681595
transform 1 0 3496 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_46
timestamp 1604681595
transform 1 0 5336 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_54
timestamp 1604681595
transform 1 0 6072 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_72
timestamp 1604681595
transform 1 0 7728 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_77
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_100
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1604681595
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_108
timestamp 1604681595
transform 1 0 11040 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_128
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_140
timestamp 1604681595
transform 1 0 13984 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_11
timestamp 1604681595
transform 1 0 2116 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2668 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_40
timestamp 1604681595
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_47
timestamp 1604681595
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_57
timestamp 1604681595
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1604681595
transform 1 0 5980 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6992 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_66
timestamp 1604681595
transform 1 0 7176 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_72
timestamp 1604681595
transform 1 0 7728 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_77
timestamp 1604681595
transform 1 0 8188 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_82
timestamp 1604681595
transform 1 0 8648 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10304 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1604681595
transform 1 0 11132 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_111
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1604681595
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1604681595
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_139
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_145
timestamp 1604681595
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_126
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_138
timestamp 1604681595
transform 1 0 13800 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_34
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_42
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_45
timestamp 1604681595
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_49
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_53
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_68
timestamp 1604681595
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_72
timestamp 1604681595
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_76
timestamp 1604681595
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_89
timestamp 1604681595
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp 1604681595
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_112
timestamp 1604681595
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_116
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_126
timestamp 1604681595
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_130
timestamp 1604681595
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_134
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_138
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_40
timestamp 1604681595
transform 1 0 4784 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5060 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7544 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_64
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_79
timestamp 1604681595
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_83
timestamp 1604681595
transform 1 0 8740 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1604681595
transform 1 0 9292 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1604681595
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_106
timestamp 1604681595
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1604681595
transform 1 0 12052 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_125
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_136
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_144
timestamp 1604681595
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_9
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_13
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_46
timestamp 1604681595
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_50
timestamp 1604681595
transform 1 0 5704 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_54
timestamp 1604681595
transform 1 0 6072 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 8648 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604681595
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_79
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_85
timestamp 1604681595
transform 1 0 8924 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_91
timestamp 1604681595
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_104
timestamp 1604681595
transform 1 0 10672 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_108
timestamp 1604681595
transform 1 0 11040 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_111
timestamp 1604681595
transform 1 0 11316 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_115
timestamp 1604681595
transform 1 0 11684 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_132
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_144
timestamp 1604681595
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_38
timestamp 1604681595
transform 1 0 4600 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_41
timestamp 1604681595
transform 1 0 4876 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1604681595
transform 1 0 5244 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_65
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_69
timestamp 1604681595
transform 1 0 7452 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_82
timestamp 1604681595
transform 1 0 8648 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9292 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1604681595
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_101
timestamp 1604681595
transform 1 0 10396 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11132 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_38_128
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_140
timestamp 1604681595
transform 1 0 13984 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_31
timestamp 1604681595
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_35
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4876 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_52
timestamp 1604681595
transform 1 0 5888 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_60
timestamp 1604681595
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_48
timestamp 1604681595
transform 1 0 5520 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_64
timestamp 1604681595
transform 1 0 6992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_85
timestamp 1604681595
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_102
timestamp 1604681595
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_102
timestamp 1604681595
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_106
timestamp 1604681595
transform 1 0 10856 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_106
timestamp 1604681595
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_110
timestamp 1604681595
transform 1 0 11224 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_122
timestamp 1604681595
transform 1 0 12328 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_143
timestamp 1604681595
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_134
timestamp 1604681595
transform 1 0 13432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_9
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_13
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4508 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4140 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 6072 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_48
timestamp 1604681595
transform 1 0 5520 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_52
timestamp 1604681595
transform 1 0 5888 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_56
timestamp 1604681595
transform 1 0 6256 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8740 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_75
timestamp 1604681595
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_79
timestamp 1604681595
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_92
timestamp 1604681595
transform 1 0 9568 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_96
timestamp 1604681595
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11316 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_109
timestamp 1604681595
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1604681595
transform 1 0 11500 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1604681595
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_143
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2576 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2944 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_18
timestamp 1604681595
transform 1 0 2760 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_22
timestamp 1604681595
transform 1 0 3128 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1604681595
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_41
timestamp 1604681595
transform 1 0 4876 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 5612 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_45
timestamp 1604681595
transform 1 0 5244 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_52
timestamp 1604681595
transform 1 0 5888 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_64
timestamp 1604681595
transform 1 0 6992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_71
timestamp 1604681595
transform 1 0 7636 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10028 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_84
timestamp 1604681595
transform 1 0 8832 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1604681595
transform 1 0 9200 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_99
timestamp 1604681595
transform 1 0 10212 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_119
timestamp 1604681595
transform 1 0 12052 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_131
timestamp 1604681595
transform 1 0 13156 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_143
timestamp 1604681595
transform 1 0 14260 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2576 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 1656 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_8
timestamp 1604681595
transform 1 0 1840 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_12
timestamp 1604681595
transform 1 0 2208 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4876 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_35
timestamp 1604681595
transform 1 0 4324 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_39
timestamp 1604681595
transform 1 0 4692 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5060 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6072 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_52
timestamp 1604681595
transform 1 0 5888 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_56
timestamp 1604681595
transform 1 0 6256 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_60
timestamp 1604681595
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8648 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_74
timestamp 1604681595
transform 1 0 7912 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_77
timestamp 1604681595
transform 1 0 8188 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_81
timestamp 1604681595
transform 1 0 8556 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9108 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 8832 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_106
timestamp 1604681595
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_110
timestamp 1604681595
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_135
timestamp 1604681595
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_143
timestamp 1604681595
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_11
timestamp 1604681595
transform 1 0 2116 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4876 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_23
timestamp 1604681595
transform 1 0 3220 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604681595
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_32
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_40
timestamp 1604681595
transform 1 0 4784 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6808 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_60
timestamp 1604681595
transform 1 0 6624 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8648 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7268 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7636 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_64
timestamp 1604681595
transform 1 0 6992 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_69
timestamp 1604681595
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_73
timestamp 1604681595
transform 1 0 7820 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_81
timestamp 1604681595
transform 1 0 8556 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10028 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_84
timestamp 1604681595
transform 1 0 8832 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_89
timestamp 1604681595
transform 1 0 9292 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_93
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_116
timestamp 1604681595
transform 1 0 11776 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_128
timestamp 1604681595
transform 1 0 12880 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_140
timestamp 1604681595
transform 1 0 13984 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1604681595
transform 1 0 1748 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_19
timestamp 1604681595
transform 1 0 2852 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3220 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_44
timestamp 1604681595
transform 1 0 5152 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_48
timestamp 1604681595
transform 1 0 5520 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_51
timestamp 1604681595
transform 1 0 5796 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_55
timestamp 1604681595
transform 1 0 6164 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8464 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_71
timestamp 1604681595
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_75
timestamp 1604681595
transform 1 0 8004 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_79
timestamp 1604681595
transform 1 0 8372 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9660 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_91
timestamp 1604681595
transform 1 0 9476 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_95
timestamp 1604681595
transform 1 0 9844 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1604681595
transform 1 0 10948 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1604681595
transform 1 0 11316 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_114
timestamp 1604681595
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1604681595
transform 1 0 11960 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1604681595
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1604681595
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_9
timestamp 1604681595
transform 1 0 1932 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1604681595
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_21
timestamp 1604681595
transform 1 0 3036 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1604681595
transform 1 0 3772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1604681595
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_39
timestamp 1604681595
transform 1 0 4692 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_48
timestamp 1604681595
transform 1 0 5520 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_45
timestamp 1604681595
transform 1 0 5244 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 5336 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5152 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 5336 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 5704 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1604681595
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_53
timestamp 1604681595
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_58
timestamp 1604681595
transform 1 0 6440 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6808 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7268 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8740 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8648 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_64
timestamp 1604681595
transform 1 0 6992 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_76
timestamp 1604681595
transform 1 0 8096 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_81
timestamp 1604681595
transform 1 0 8556 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 9292 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 9108 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_84
timestamp 1604681595
transform 1 0 8832 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_90
timestamp 1604681595
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_85
timestamp 1604681595
transform 1 0 8924 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_92
timestamp 1604681595
transform 1 0 9568 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_104
timestamp 1604681595
transform 1 0 10672 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_111
timestamp 1604681595
transform 1 0 11316 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_108
timestamp 1604681595
transform 1 0 11040 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_111
timestamp 1604681595
transform 1 0 11316 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_105
timestamp 1604681595
transform 1 0 10764 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_119
timestamp 1604681595
transform 1 0 12052 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_115
timestamp 1604681595
transform 1 0 11684 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11408 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_46_131
timestamp 1604681595
transform 1 0 13156 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_143
timestamp 1604681595
transform 1 0 14260 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1604681595
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_143
timestamp 1604681595
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1604681595
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4508 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4876 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1604681595
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_32
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_36
timestamp 1604681595
transform 1 0 4416 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_39
timestamp 1604681595
transform 1 0 4692 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6808 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_43
timestamp 1604681595
transform 1 0 5060 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_51
timestamp 1604681595
transform 1 0 5796 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_56
timestamp 1604681595
transform 1 0 6256 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_60
timestamp 1604681595
transform 1 0 6624 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7268 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 6992 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_76
timestamp 1604681595
transform 1 0 8096 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_80
timestamp 1604681595
transform 1 0 8464 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_88
timestamp 1604681595
transform 1 0 9200 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_84
timestamp 1604681595
transform 1 0 8832 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_97
timestamp 1604681595
transform 1 0 10028 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_101
timestamp 1604681595
transform 1 0 10396 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 10212 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11500 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12512 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10948 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_105
timestamp 1604681595
transform 1 0 10764 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_109
timestamp 1604681595
transform 1 0 11132 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_122
timestamp 1604681595
transform 1 0 12328 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 13064 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12880 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_126
timestamp 1604681595
transform 1 0 12696 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_133
timestamp 1604681595
transform 1 0 13340 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1604681595
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1604681595
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4508 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4324 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3956 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1604681595
transform 1 0 3588 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_33
timestamp 1604681595
transform 1 0 4140 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5520 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_46
timestamp 1604681595
transform 1 0 5336 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_50
timestamp 1604681595
transform 1 0 5704 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_54
timestamp 1604681595
transform 1 0 6072 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1604681595
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8648 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_71
timestamp 1604681595
transform 1 0 7636 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_77
timestamp 1604681595
transform 1 0 8188 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 10212 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_91
timestamp 1604681595
transform 1 0 9476 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_95
timestamp 1604681595
transform 1 0 9844 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_102
timestamp 1604681595
transform 1 0 10488 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12512 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_112
timestamp 1604681595
transform 1 0 11408 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_118
timestamp 1604681595
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_123
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13524 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_133
timestamp 1604681595
transform 1 0 13340 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_137
timestamp 1604681595
transform 1 0 13708 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_145
timestamp 1604681595
transform 1 0 14444 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1604681595
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1604681595
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_32
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_36
timestamp 1604681595
transform 1 0 4416 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6808 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_58
timestamp 1604681595
transform 1 0 6440 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_64
timestamp 1604681595
transform 1 0 6992 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_69
timestamp 1604681595
transform 1 0 7452 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_84
timestamp 1604681595
transform 1 0 8832 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_112
timestamp 1604681595
transform 1 0 11408 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13156 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_129
timestamp 1604681595
transform 1 0 12972 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_133
timestamp 1604681595
transform 1 0 13340 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1604681595
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 1932 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_11
timestamp 1604681595
transform 1 0 2116 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3772 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3220 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_25
timestamp 1604681595
transform 1 0 3404 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_38
timestamp 1604681595
transform 1 0 4600 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_42
timestamp 1604681595
transform 1 0 4968 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 5336 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_49
timestamp 1604681595
transform 1 0 5612 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 5796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_53
timestamp 1604681595
transform 1 0 5980 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1604681595
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_62
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7268 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_86
timestamp 1604681595
transform 1 0 9016 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_90
timestamp 1604681595
transform 1 0 9384 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1604681595
transform 1 0 11500 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1604681595
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 13800 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_132
timestamp 1604681595
transform 1 0 13248 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_136
timestamp 1604681595
transform 1 0 13616 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_140
timestamp 1604681595
transform 1 0 13984 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_13
timestamp 1604681595
transform 1 0 2300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1604681595
transform 1 0 1932 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_13
timestamp 1604681595
transform 1 0 2300 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_7
timestamp 1604681595
transform 1 0 1748 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1932 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_20
timestamp 1604681595
transform 1 0 2944 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_16
timestamp 1604681595
transform 1 0 2576 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_17
timestamp 1604681595
transform 1 0 2668 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2852 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_26
timestamp 1604681595
transform 1 0 3496 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_21
timestamp 1604681595
transform 1 0 3036 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3128 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3312 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_37
timestamp 1604681595
transform 1 0 4508 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_33
timestamp 1604681595
transform 1 0 4140 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4692 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_41
timestamp 1604681595
transform 1 0 4876 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4876 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_50
timestamp 1604681595
transform 1 0 5704 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_52
timestamp 1604681595
transform 1 0 5888 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_47
timestamp 1604681595
transform 1 0 5428 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5244 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5888 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 5612 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_58
timestamp 1604681595
transform 1 0 6440 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_54
timestamp 1604681595
transform 1 0 6072 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_56
timestamp 1604681595
transform 1 0 6256 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6624 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8188 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8556 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_79
timestamp 1604681595
transform 1 0 8372 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_83
timestamp 1604681595
transform 1 0 8740 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_71
timestamp 1604681595
transform 1 0 7636 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_75
timestamp 1604681595
transform 1 0 8004 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_92
timestamp 1604681595
transform 1 0 9568 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_88
timestamp 1604681595
transform 1 0 9200 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_93
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1604681595
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_100
timestamp 1604681595
transform 1 0 10304 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_96
timestamp 1604681595
transform 1 0 9936 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_98
timestamp 1604681595
transform 1 0 10120 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9752 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10304 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10120 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10488 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_53_104
timestamp 1604681595
transform 1 0 10672 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_114
timestamp 1604681595
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_111
timestamp 1604681595
transform 1 0 11316 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11500 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_53_123
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_118
timestamp 1604681595
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_115
timestamp 1604681595
transform 1 0 11684 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11868 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12512 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12052 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13524 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_138
timestamp 1604681595
transform 1 0 13800 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_133
timestamp 1604681595
transform 1 0 13340 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_137
timestamp 1604681595
transform 1 0 13708 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_145
timestamp 1604681595
transform 1 0 14444 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_3
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_11
timestamp 1604681595
transform 1 0 2116 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4876 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_23
timestamp 1604681595
transform 1 0 3220 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_32
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_36
timestamp 1604681595
transform 1 0 4416 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_39
timestamp 1604681595
transform 1 0 4692 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5244 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_43
timestamp 1604681595
transform 1 0 5060 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_54
timestamp 1604681595
transform 1 0 6072 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_58
timestamp 1604681595
transform 1 0 6440 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_71
timestamp 1604681595
transform 1 0 7636 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_75
timestamp 1604681595
transform 1 0 8004 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1604681595
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_86
timestamp 1604681595
transform 1 0 9016 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_93
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_99
timestamp 1604681595
transform 1 0 10212 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12052 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11500 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_111
timestamp 1604681595
transform 1 0 11316 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_115
timestamp 1604681595
transform 1 0 11684 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_138
timestamp 1604681595
transform 1 0 13800 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_9
timestamp 1604681595
transform 1 0 1932 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_13
timestamp 1604681595
transform 1 0 2300 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_17
timestamp 1604681595
transform 1 0 2668 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_20
timestamp 1604681595
transform 1 0 2944 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3312 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4876 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3128 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_33
timestamp 1604681595
transform 1 0 4140 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_37
timestamp 1604681595
transform 1 0 4508 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_40
timestamp 1604681595
transform 1 0 4784 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_50
timestamp 1604681595
transform 1 0 5704 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_54
timestamp 1604681595
transform 1 0 6072 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1604681595
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_62
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7268 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8648 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8280 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_66
timestamp 1604681595
transform 1 0 7176 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_76
timestamp 1604681595
transform 1 0 8096 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_80
timestamp 1604681595
transform 1 0 8464 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8832 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10488 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_93
timestamp 1604681595
transform 1 0 9660 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_97
timestamp 1604681595
transform 1 0 10028 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_100
timestamp 1604681595
transform 1 0 10304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_104
timestamp 1604681595
transform 1 0 10672 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10856 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_108
timestamp 1604681595
transform 1 0 11040 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_118
timestamp 1604681595
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_132
timestamp 1604681595
transform 1 0 13248 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_144
timestamp 1604681595
transform 1 0 14352 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2944 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_15
timestamp 1604681595
transform 1 0 2484 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_19
timestamp 1604681595
transform 1 0 2852 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 4600 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4416 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_22
timestamp 1604681595
transform 1 0 3128 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1604681595
transform 1 0 3496 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_30
timestamp 1604681595
transform 1 0 3864 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_32
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6624 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5520 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_42
timestamp 1604681595
transform 1 0 4968 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_46
timestamp 1604681595
transform 1 0 5336 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_50
timestamp 1604681595
transform 1 0 5704 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_58
timestamp 1604681595
transform 1 0 6440 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_62
timestamp 1604681595
transform 1 0 6808 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_56_72
timestamp 1604681595
transform 1 0 7728 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10120 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9844 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_86
timestamp 1604681595
transform 1 0 9016 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_90
timestamp 1604681595
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_97
timestamp 1604681595
transform 1 0 10028 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_107
timestamp 1604681595
transform 1 0 10948 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_119
timestamp 1604681595
transform 1 0 12052 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_125
timestamp 1604681595
transform 1 0 12604 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_137
timestamp 1604681595
transform 1 0 13708 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_145
timestamp 1604681595
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 1748 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_19
timestamp 1604681595
transform 1 0 2852 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_15
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_11
timestamp 1604681595
transform 1 0 2116 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 2668 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 2300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2944 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4876 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_39
timestamp 1604681595
transform 1 0 4692 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 5428 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5244 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_43
timestamp 1604681595
transform 1 0 5060 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_51
timestamp 1604681595
transform 1 0 5796 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_55
timestamp 1604681595
transform 1 0 6164 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 8648 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1604681595
transform 1 0 7636 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_75
timestamp 1604681595
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_79
timestamp 1604681595
transform 1 0 8372 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8832 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_57_103
timestamp 1604681595
transform 1 0 10580 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 11316 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10764 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_107
timestamp 1604681595
transform 1 0 10948 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_114
timestamp 1604681595
transform 1 0 11592 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1604681595
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_143
timestamp 1604681595
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 2668 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_9
timestamp 1604681595
transform 1 0 1932 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4140 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3404 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_21
timestamp 1604681595
transform 1 0 3036 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1604681595
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_32
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6624 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_52
timestamp 1604681595
transform 1 0 5888 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8556 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_79
timestamp 1604681595
transform 1 0 8372 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_83
timestamp 1604681595
transform 1 0 8740 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9844 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_87
timestamp 1604681595
transform 1 0 9108 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_91
timestamp 1604681595
transform 1 0 9476 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_114
timestamp 1604681595
transform 1 0 11592 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_126
timestamp 1604681595
transform 1 0 12696 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_138
timestamp 1604681595
transform 1 0 13800 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_11
timestamp 1604681595
transform 1 0 2116 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_7
timestamp 1604681595
transform 1 0 1748 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_13
timestamp 1604681595
transform 1 0 2300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_9
timestamp 1604681595
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 2116 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_19
timestamp 1604681595
transform 1 0 2852 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_17
timestamp 1604681595
transform 1 0 2668 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 2484 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3404 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 3220 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1604681595
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_36
timestamp 1604681595
transform 1 0 4416 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 5796 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 5796 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_44
timestamp 1604681595
transform 1 0 5152 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_50
timestamp 1604681595
transform 1 0 5704 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_53
timestamp 1604681595
transform 1 0 5980 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_62
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_48
timestamp 1604681595
transform 1 0 5520 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_55
timestamp 1604681595
transform 1 0 6164 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_71
timestamp 1604681595
transform 1 0 7636 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_67
timestamp 1604681595
transform 1 0 7268 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_72
timestamp 1604681595
transform 1 0 7728 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_66
timestamp 1604681595
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 6992 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 7360 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 6900 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_76
timestamp 1604681595
transform 1 0 8096 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8280 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 7912 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_60_93
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_88
timestamp 1604681595
transform 1 0 9200 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_84
timestamp 1604681595
transform 1 0 8832 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_93
timestamp 1604681595
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_89
timestamp 1604681595
transform 1 0 9292 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9476 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9936 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10028 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10120 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_59_114
timestamp 1604681595
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1604681595
transform 1 0 11224 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_106
timestamp 1604681595
transform 1 0 10856 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11040 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_118
timestamp 1604681595
transform 1 0 11960 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_119
timestamp 1604681595
transform 1 0 12052 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_107
timestamp 1604681595
transform 1 0 10948 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_135
timestamp 1604681595
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_143
timestamp 1604681595
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_131
timestamp 1604681595
transform 1 0 13156 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_143
timestamp 1604681595
transform 1 0 14260 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 1932 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_7
timestamp 1604681595
transform 1 0 1748 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_11
timestamp 1604681595
transform 1 0 2116 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_19
timestamp 1604681595
transform 1 0 2852 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 4232 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 4784 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 3036 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 4048 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_23
timestamp 1604681595
transform 1 0 3220 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_31
timestamp 1604681595
transform 1 0 3956 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_38
timestamp 1604681595
transform 1 0 4600 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 5612 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 5336 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 6164 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_42
timestamp 1604681595
transform 1 0 4968 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_48
timestamp 1604681595
transform 1 0 5520 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_53
timestamp 1604681595
transform 1 0 5980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 1604681595
transform 1 0 6348 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 7912 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 7360 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 8464 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_66
timestamp 1604681595
transform 1 0 7176 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_70
timestamp 1604681595
transform 1 0 7544 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_78
timestamp 1604681595
transform 1 0 8280 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_82
timestamp 1604681595
transform 1 0 8648 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 9016 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 9568 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_90
timestamp 1604681595
transform 1 0 9384 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1604681595
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_106
timestamp 1604681595
transform 1 0 10856 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_118
timestamp 1604681595
transform 1 0 11960 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604681595
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604681595
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 4232 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_38
timestamp 1604681595
transform 1 0 4600 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 5336 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_50
timestamp 1604681595
transform 1 0 5704 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_62
timestamp 1604681595
transform 1 0 6808 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_74
timestamp 1604681595
transform 1 0 7912 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_86
timestamp 1604681595
transform 1 0 9016 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604681595
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604681595
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1604681595
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1604681595
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604681595
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604681595
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604681595
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604681595
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604681595
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604681595
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604681595
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604681595
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604681595
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 1096 480 1216 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 29928 16000 30048 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_16_
port 82 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 left_grid_pin_17_
port 83 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_18_
port 84 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 left_grid_pin_19_
port 85 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_20_
port 86 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_21_
port 87 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_22_
port 88 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 left_grid_pin_23_
port 89 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 left_grid_pin_24_
port 90 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 left_grid_pin_25_
port 91 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_26_
port 92 nsew default tristate
rlabel metal3 s 0 29248 480 29368 6 left_grid_pin_27_
port 93 nsew default tristate
rlabel metal3 s 0 31560 480 31680 6 left_grid_pin_28_
port 94 nsew default tristate
rlabel metal3 s 0 34008 480 34128 6 left_grid_pin_29_
port 95 nsew default tristate
rlabel metal3 s 0 36320 480 36440 6 left_grid_pin_30_
port 96 nsew default tristate
rlabel metal3 s 0 38632 480 38752 6 left_grid_pin_31_
port 97 nsew default tristate
rlabel metal3 s 15520 9936 16000 10056 6 prog_clk
port 98 nsew default input
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 99 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
