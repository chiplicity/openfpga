magic
tech EFS8A
magscale 1 2
timestamp 1603803781
<< locali >>
rect 2789 12631 2823 12733
rect 8677 10455 8711 10557
rect 28457 8823 28491 9129
rect 34437 8347 34471 8585
rect 21465 7191 21499 7497
rect 26617 5083 26651 5253
<< viali >>
rect 1593 12937 1627 12971
rect 35633 12937 35667 12971
rect 1409 12733 1443 12767
rect 2580 12733 2614 12767
rect 2789 12733 2823 12767
rect 4972 12733 5006 12767
rect 13001 12733 13035 12767
rect 35449 12733 35483 12767
rect 36001 12733 36035 12767
rect 2053 12665 2087 12699
rect 2651 12597 2685 12631
rect 2789 12597 2823 12631
rect 3065 12597 3099 12631
rect 5043 12597 5077 12631
rect 5457 12597 5491 12631
rect 13185 12597 13219 12631
rect 13553 12597 13587 12631
rect 1593 12393 1627 12427
rect 1409 12257 1443 12291
rect 2513 12257 2547 12291
rect 4144 12257 4178 12291
rect 5952 12257 5986 12291
rect 10241 12257 10275 12291
rect 11320 12257 11354 12291
rect 13093 12257 13127 12291
rect 2053 12053 2087 12087
rect 2421 12053 2455 12087
rect 2697 12053 2731 12087
rect 4215 12053 4249 12087
rect 6055 12053 6089 12087
rect 10425 12053 10459 12087
rect 11391 12053 11425 12087
rect 13277 12053 13311 12087
rect 14289 12053 14323 12087
rect 2881 11849 2915 11883
rect 2053 11645 2087 11679
rect 2421 11645 2455 11679
rect 3433 11645 3467 11679
rect 4940 11645 4974 11679
rect 5365 11645 5399 11679
rect 6904 11645 6938 11679
rect 7297 11645 7331 11679
rect 10241 11645 10275 11679
rect 11069 11645 11103 11679
rect 11288 11645 11322 11679
rect 11713 11645 11747 11679
rect 14289 11645 14323 11679
rect 14749 11645 14783 11679
rect 18464 11645 18498 11679
rect 18889 11645 18923 11679
rect 19752 11645 19786 11679
rect 20177 11645 20211 11679
rect 2605 11577 2639 11611
rect 4169 11577 4203 11611
rect 10701 11577 10735 11611
rect 15025 11577 15059 11611
rect 1685 11509 1719 11543
rect 3341 11509 3375 11543
rect 3617 11509 3651 11543
rect 5043 11509 5077 11543
rect 5917 11509 5951 11543
rect 6975 11509 7009 11543
rect 10425 11509 10459 11543
rect 11391 11509 11425 11543
rect 12173 11509 12207 11543
rect 12449 11509 12483 11543
rect 13185 11509 13219 11543
rect 14105 11509 14139 11543
rect 18567 11509 18601 11543
rect 19855 11509 19889 11543
rect 17003 11305 17037 11339
rect 35633 11305 35667 11339
rect 1869 11169 1903 11203
rect 2421 11169 2455 11203
rect 4144 11169 4178 11203
rect 4629 11169 4663 11203
rect 5156 11169 5190 11203
rect 6168 11169 6202 11203
rect 7148 11169 7182 11203
rect 8192 11169 8226 11203
rect 9689 11169 9723 11203
rect 10768 11169 10802 11203
rect 11805 11169 11839 11203
rect 13645 11169 13679 11203
rect 14105 11169 14139 11203
rect 16900 11169 16934 11203
rect 18496 11169 18530 11203
rect 19508 11169 19542 11203
rect 22084 11169 22118 11203
rect 26652 11169 26686 11203
rect 34380 11169 34414 11203
rect 35449 11169 35483 11203
rect 2329 11101 2363 11135
rect 12449 11101 12483 11135
rect 14381 11101 14415 11135
rect 15669 11101 15703 11135
rect 4215 11033 4249 11067
rect 5227 11033 5261 11067
rect 6239 11033 6273 11067
rect 7251 11033 7285 11067
rect 9873 11033 9907 11067
rect 10839 11033 10873 11067
rect 18567 11033 18601 11067
rect 19579 11033 19613 11067
rect 22155 11033 22189 11067
rect 26755 11033 26789 11067
rect 1777 10965 1811 10999
rect 8263 10965 8297 10999
rect 13461 10965 13495 10999
rect 34483 10965 34517 10999
rect 1593 10761 1627 10795
rect 4537 10761 4571 10795
rect 5871 10761 5905 10795
rect 7481 10761 7515 10795
rect 8585 10761 8619 10795
rect 15301 10761 15335 10795
rect 18521 10761 18555 10795
rect 26249 10761 26283 10795
rect 35633 10761 35667 10795
rect 2605 10693 2639 10727
rect 4169 10625 4203 10659
rect 13645 10625 13679 10659
rect 15761 10625 15795 10659
rect 19533 10625 19567 10659
rect 1409 10557 1443 10591
rect 2789 10557 2823 10591
rect 3341 10557 3375 10591
rect 4353 10557 4387 10591
rect 5800 10557 5834 10591
rect 6561 10557 6595 10591
rect 8033 10557 8067 10591
rect 8677 10557 8711 10591
rect 10368 10557 10402 10591
rect 10793 10557 10827 10591
rect 11380 10557 11414 10591
rect 11805 10557 11839 10591
rect 12265 10557 12299 10591
rect 12541 10557 12575 10591
rect 14105 10557 14139 10591
rect 14565 10557 14599 10591
rect 15853 10557 15887 10591
rect 16313 10557 16347 10591
rect 18096 10557 18130 10591
rect 18889 10557 18923 10591
rect 19108 10557 19142 10591
rect 19901 10557 19935 10591
rect 20856 10557 20890 10591
rect 21281 10557 21315 10591
rect 21868 10557 21902 10591
rect 25732 10557 25766 10591
rect 25835 10557 25869 10591
rect 26744 10557 26778 10591
rect 27169 10557 27203 10591
rect 27788 10557 27822 10591
rect 28181 10557 28215 10591
rect 33308 10557 33342 10591
rect 35265 10557 35299 10591
rect 35449 10557 35483 10591
rect 36001 10557 36035 10591
rect 3525 10489 3559 10523
rect 9321 10489 9355 10523
rect 11483 10489 11517 10523
rect 14841 10489 14875 10523
rect 22661 10489 22695 10523
rect 26847 10489 26881 10523
rect 2053 10421 2087 10455
rect 5181 10421 5215 10455
rect 6193 10421 6227 10455
rect 7021 10421 7055 10455
rect 8217 10421 8251 10455
rect 8677 10421 8711 10455
rect 8953 10421 8987 10455
rect 9781 10421 9815 10455
rect 10471 10421 10505 10455
rect 11253 10421 11287 10455
rect 12909 10421 12943 10455
rect 16129 10421 16163 10455
rect 16865 10421 16899 10455
rect 18199 10421 18233 10455
rect 19211 10421 19245 10455
rect 20959 10421 20993 10455
rect 21971 10421 22005 10455
rect 22385 10421 22419 10455
rect 26617 10421 26651 10455
rect 27859 10421 27893 10455
rect 33379 10421 33413 10455
rect 33793 10421 33827 10455
rect 34437 10421 34471 10455
rect 2421 10217 2455 10251
rect 3525 10217 3559 10251
rect 6929 10217 6963 10251
rect 10793 10217 10827 10251
rect 13461 10217 13495 10251
rect 14105 10217 14139 10251
rect 27169 10217 27203 10251
rect 35633 10217 35667 10251
rect 27445 10149 27479 10183
rect 1685 10081 1719 10115
rect 1869 10081 1903 10115
rect 3040 10081 3074 10115
rect 4261 10081 4295 10115
rect 4537 10081 4571 10115
rect 5708 10081 5742 10115
rect 6653 10081 6687 10115
rect 7113 10081 7147 10115
rect 8652 10081 8686 10115
rect 10517 10081 10551 10115
rect 11069 10081 11103 10115
rect 12817 10081 12851 10115
rect 15853 10081 15887 10115
rect 16313 10081 16347 10115
rect 17969 10081 18003 10115
rect 18245 10081 18279 10115
rect 19384 10081 19418 10115
rect 20948 10081 20982 10115
rect 21960 10081 21994 10115
rect 22937 10081 22971 10115
rect 24409 10081 24443 10115
rect 25488 10081 25522 10115
rect 28892 10081 28926 10115
rect 33460 10081 33494 10115
rect 34504 10081 34538 10115
rect 35449 10081 35483 10115
rect 36620 10081 36654 10115
rect 1961 10013 1995 10047
rect 4629 10013 4663 10047
rect 13185 10013 13219 10047
rect 16405 10013 16439 10047
rect 18337 10013 18371 10047
rect 21465 10013 21499 10047
rect 27353 10013 27387 10047
rect 27997 10013 28031 10047
rect 12955 9945 12989 9979
rect 22063 9945 22097 9979
rect 2789 9877 2823 9911
rect 3111 9877 3145 9911
rect 5779 9877 5813 9911
rect 8723 9877 8757 9911
rect 11713 9877 11747 9911
rect 12541 9877 12575 9911
rect 13093 9877 13127 9911
rect 14473 9877 14507 9911
rect 19487 9877 19521 9911
rect 19901 9877 19935 9911
rect 21051 9877 21085 9911
rect 21741 9877 21775 9911
rect 23121 9877 23155 9911
rect 24133 9877 24167 9911
rect 24593 9877 24627 9911
rect 25559 9877 25593 9911
rect 28963 9877 28997 9911
rect 33563 9877 33597 9911
rect 34575 9877 34609 9911
rect 36691 9877 36725 9911
rect 2881 9673 2915 9707
rect 6285 9673 6319 9707
rect 8217 9673 8251 9707
rect 10241 9673 10275 9707
rect 11529 9673 11563 9707
rect 13461 9673 13495 9707
rect 15393 9673 15427 9707
rect 19349 9673 19383 9707
rect 20913 9673 20947 9707
rect 25513 9673 25547 9707
rect 33425 9673 33459 9707
rect 3985 9605 4019 9639
rect 6561 9605 6595 9639
rect 11805 9605 11839 9639
rect 13829 9605 13863 9639
rect 15853 9605 15887 9639
rect 32321 9605 32355 9639
rect 35541 9605 35575 9639
rect 36645 9605 36679 9639
rect 3065 9537 3099 9571
rect 7205 9537 7239 9571
rect 12265 9537 12299 9571
rect 12541 9537 12575 9571
rect 14381 9537 14415 9571
rect 16037 9537 16071 9571
rect 16957 9537 16991 9571
rect 21741 9537 21775 9571
rect 24777 9537 24811 9571
rect 27445 9537 27479 9571
rect 32597 9537 32631 9571
rect 35173 9537 35207 9571
rect 1685 9469 1719 9503
rect 1961 9469 1995 9503
rect 4445 9469 4479 9503
rect 4629 9469 4663 9503
rect 8401 9469 8435 9503
rect 8861 9469 8895 9503
rect 10517 9469 10551 9503
rect 10977 9469 11011 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 19625 9469 19659 9503
rect 20085 9469 20119 9503
rect 22477 9469 22511 9503
rect 24409 9469 24443 9503
rect 24593 9469 24627 9503
rect 26408 9469 26442 9503
rect 29352 9469 29386 9503
rect 30297 9469 30331 9503
rect 30757 9469 30791 9503
rect 31836 9469 31870 9503
rect 32816 9469 32850 9503
rect 33860 9469 33894 9503
rect 35357 9469 35391 9503
rect 36461 9469 36495 9503
rect 37013 9469 37047 9503
rect 2145 9401 2179 9435
rect 3157 9401 3191 9435
rect 3709 9401 3743 9435
rect 5273 9401 5307 9435
rect 6929 9401 6963 9435
rect 7021 9401 7055 9435
rect 9965 9401 9999 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 16129 9401 16163 9435
rect 16681 9401 16715 9435
rect 21465 9401 21499 9435
rect 21557 9401 21591 9435
rect 22937 9401 22971 9435
rect 24041 9401 24075 9435
rect 27261 9401 27295 9435
rect 27537 9401 27571 9435
rect 28089 9401 28123 9435
rect 34345 9401 34379 9435
rect 2513 9333 2547 9367
rect 5733 9333 5767 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 9413 9333 9447 9367
rect 10517 9333 10551 9367
rect 17417 9333 17451 9367
rect 17785 9333 17819 9367
rect 18153 9333 18187 9367
rect 19901 9333 19935 9367
rect 26479 9333 26513 9367
rect 26893 9333 26927 9367
rect 28365 9333 28399 9367
rect 28825 9333 28859 9367
rect 29423 9333 29457 9367
rect 29837 9333 29871 9367
rect 30481 9333 30515 9367
rect 31907 9333 31941 9367
rect 32919 9333 32953 9367
rect 33931 9333 33965 9367
rect 34713 9333 34747 9367
rect 35909 9333 35943 9367
rect 37381 9333 37415 9367
rect 1961 9129 1995 9163
rect 3893 9129 3927 9163
rect 11069 9129 11103 9163
rect 11437 9129 11471 9163
rect 12817 9129 12851 9163
rect 16221 9129 16255 9163
rect 16497 9129 16531 9163
rect 18061 9129 18095 9163
rect 18705 9129 18739 9163
rect 20085 9129 20119 9163
rect 23903 9129 23937 9163
rect 28273 9129 28307 9163
rect 28457 9129 28491 9163
rect 33609 9129 33643 9163
rect 2605 9061 2639 9095
rect 3157 9061 3191 9095
rect 4261 9061 4295 9095
rect 7389 9061 7423 9095
rect 11805 9061 11839 9095
rect 13369 9061 13403 9095
rect 15622 9061 15656 9095
rect 17233 9061 17267 9095
rect 18521 9061 18555 9095
rect 21281 9061 21315 9095
rect 21373 9061 21407 9095
rect 27445 9061 27479 9095
rect 1476 8993 1510 9027
rect 5641 8993 5675 9027
rect 5917 8993 5951 9027
rect 10057 8993 10091 9027
rect 10517 8993 10551 9027
rect 15301 8993 15335 9027
rect 18613 8993 18647 9027
rect 19165 8993 19199 9027
rect 22820 8993 22854 9027
rect 23832 8993 23866 9027
rect 24869 8993 24903 9027
rect 25329 8993 25363 9027
rect 2513 8925 2547 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 5181 8925 5215 8959
rect 6101 8925 6135 8959
rect 7297 8925 7331 8959
rect 7573 8925 7607 8959
rect 10609 8925 10643 8959
rect 11713 8925 11747 8959
rect 13277 8925 13311 8959
rect 13553 8925 13587 8959
rect 16865 8925 16899 8959
rect 17141 8925 17175 8959
rect 17417 8925 17451 8959
rect 25605 8925 25639 8959
rect 27353 8925 27387 8959
rect 27997 8925 28031 8959
rect 5733 8857 5767 8891
rect 8493 8857 8527 8891
rect 12265 8857 12299 8891
rect 21833 8857 21867 8891
rect 28641 9061 28675 9095
rect 29009 9061 29043 9095
rect 34069 9061 34103 9095
rect 35633 9061 35667 9095
rect 30424 8993 30458 9027
rect 32321 8993 32355 9027
rect 32689 8993 32723 9027
rect 28917 8925 28951 8959
rect 29193 8925 29227 8959
rect 32873 8925 32907 8959
rect 33977 8925 34011 8959
rect 34253 8925 34287 8959
rect 35541 8925 35575 8959
rect 36093 8857 36127 8891
rect 1547 8789 1581 8823
rect 2329 8789 2363 8823
rect 3525 8789 3559 8823
rect 6929 8789 6963 8823
rect 8861 8789 8895 8823
rect 19717 8789 19751 8823
rect 22293 8789 22327 8823
rect 22891 8789 22925 8823
rect 24409 8789 24443 8823
rect 27169 8789 27203 8823
rect 28457 8789 28491 8823
rect 30527 8789 30561 8823
rect 31309 8789 31343 8823
rect 33333 8789 33367 8823
rect 34989 8789 35023 8823
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 6193 8585 6227 8619
rect 8033 8585 8067 8619
rect 8677 8585 8711 8619
rect 10149 8585 10183 8619
rect 13461 8585 13495 8619
rect 17095 8585 17129 8619
rect 17877 8585 17911 8619
rect 19257 8585 19291 8619
rect 22385 8585 22419 8619
rect 22845 8585 22879 8619
rect 23949 8585 23983 8619
rect 26801 8585 26835 8619
rect 28733 8585 28767 8619
rect 34253 8585 34287 8619
rect 34437 8585 34471 8619
rect 35909 8585 35943 8619
rect 36277 8585 36311 8619
rect 36645 8585 36679 8619
rect 2421 8517 2455 8551
rect 4997 8517 5031 8551
rect 5825 8517 5859 8551
rect 8309 8517 8343 8551
rect 10425 8517 10459 8551
rect 11437 8517 11471 8551
rect 13829 8517 13863 8551
rect 15117 8517 15151 8551
rect 16497 8517 16531 8551
rect 18889 8517 18923 8551
rect 33885 8517 33919 8551
rect 1501 8449 1535 8483
rect 2145 8449 2179 8483
rect 3065 8449 3099 8483
rect 3709 8449 3743 8483
rect 5273 8449 5307 8483
rect 10885 8449 10919 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 15209 8449 15243 8483
rect 16773 8449 16807 8483
rect 18337 8449 18371 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 21465 8449 21499 8483
rect 21833 8449 21867 8483
rect 27721 8449 27755 8483
rect 29377 8449 29411 8483
rect 29653 8449 29687 8483
rect 33333 8449 33367 8483
rect 7113 8381 7147 8415
rect 8861 8381 8895 8415
rect 9321 8381 9355 8415
rect 14064 8381 14098 8415
rect 14565 8381 14599 8415
rect 16992 8381 17026 8415
rect 21189 8381 21223 8415
rect 24409 8381 24443 8415
rect 24869 8381 24903 8415
rect 25053 8381 25087 8415
rect 25881 8381 25915 8415
rect 31217 8381 31251 8415
rect 32137 8381 32171 8415
rect 35541 8517 35575 8551
rect 34989 8449 35023 8483
rect 37703 8449 37737 8483
rect 36461 8381 36495 8415
rect 37013 8381 37047 8415
rect 37600 8381 37634 8415
rect 38025 8381 38059 8415
rect 1593 8313 1627 8347
rect 2881 8313 2915 8347
rect 3157 8313 3191 8347
rect 5365 8313 5399 8347
rect 7434 8313 7468 8347
rect 10977 8313 11011 8347
rect 11897 8313 11931 8347
rect 12633 8313 12667 8347
rect 14151 8313 14185 8347
rect 15530 8313 15564 8347
rect 17417 8313 17451 8347
rect 18429 8313 18463 8347
rect 19625 8313 19659 8347
rect 19993 8313 20027 8347
rect 20821 8313 20855 8347
rect 21557 8313 21591 8347
rect 23489 8313 23523 8347
rect 25421 8313 25455 8347
rect 26243 8313 26277 8347
rect 27813 8313 27847 8347
rect 28365 8313 28399 8347
rect 29009 8313 29043 8347
rect 29469 8313 29503 8347
rect 30389 8313 30423 8347
rect 31538 8313 31572 8347
rect 32413 8313 32447 8347
rect 32781 8313 32815 8347
rect 33425 8313 33459 8347
rect 34437 8313 34471 8347
rect 34713 8313 34747 8347
rect 35081 8313 35115 8347
rect 6653 8245 6687 8279
rect 8953 8245 8987 8279
rect 12265 8245 12299 8279
rect 16129 8245 16163 8279
rect 25789 8245 25823 8279
rect 27261 8245 27295 8279
rect 31125 8245 31159 8279
rect 2053 8041 2087 8075
rect 3065 8041 3099 8075
rect 3341 8041 3375 8075
rect 3801 8041 3835 8075
rect 6653 8041 6687 8075
rect 7665 8041 7699 8075
rect 8033 8041 8067 8075
rect 8401 8041 8435 8075
rect 10517 8041 10551 8075
rect 10885 8041 10919 8075
rect 11897 8041 11931 8075
rect 12541 8041 12575 8075
rect 15117 8041 15151 8075
rect 16221 8041 16255 8075
rect 19809 8041 19843 8075
rect 22109 8041 22143 8075
rect 23673 8041 23707 8075
rect 25881 8041 25915 8075
rect 27445 8041 27479 8075
rect 27813 8041 27847 8075
rect 28089 8041 28123 8075
rect 33425 8041 33459 8075
rect 34345 8041 34379 8075
rect 35909 8041 35943 8075
rect 36645 8041 36679 8075
rect 2507 7973 2541 8007
rect 4169 7973 4203 8007
rect 4261 7973 4295 8007
rect 4813 7973 4847 8007
rect 7107 7973 7141 8007
rect 11339 7973 11373 8007
rect 12909 7973 12943 8007
rect 15642 7973 15676 8007
rect 17233 7973 17267 8007
rect 17785 7973 17819 8007
rect 18975 7973 19009 8007
rect 21281 7973 21315 8007
rect 21833 7973 21867 8007
rect 22845 7973 22879 8007
rect 26846 7973 26880 8007
rect 28641 7973 28675 8007
rect 32458 7973 32492 8007
rect 35081 7973 35115 8007
rect 2145 7905 2179 7939
rect 5641 7905 5675 7939
rect 6745 7905 6779 7939
rect 8493 7905 8527 7939
rect 10000 7905 10034 7939
rect 10977 7905 11011 7939
rect 15301 7905 15335 7939
rect 18613 7905 18647 7939
rect 19533 7905 19567 7939
rect 24869 7905 24903 7939
rect 25329 7905 25363 7939
rect 30757 7905 30791 7939
rect 31033 7905 31067 7939
rect 33057 7905 33091 7939
rect 33920 7905 33954 7939
rect 36461 7905 36495 7939
rect 6285 7837 6319 7871
rect 10103 7837 10137 7871
rect 12173 7837 12207 7871
rect 12817 7837 12851 7871
rect 13461 7837 13495 7871
rect 16497 7837 16531 7871
rect 17141 7837 17175 7871
rect 21189 7837 21223 7871
rect 22753 7837 22787 7871
rect 23397 7837 23431 7871
rect 24777 7837 24811 7871
rect 25605 7837 25639 7871
rect 26525 7837 26559 7871
rect 28549 7837 28583 7871
rect 29193 7837 29227 7871
rect 31217 7837 31251 7871
rect 32137 7837 32171 7871
rect 34989 7837 35023 7871
rect 35633 7837 35667 7871
rect 5825 7769 5859 7803
rect 20729 7769 20763 7803
rect 34805 7769 34839 7803
rect 1685 7701 1719 7735
rect 5273 7701 5307 7735
rect 8677 7701 8711 7735
rect 16865 7701 16899 7735
rect 18337 7701 18371 7735
rect 24409 7701 24443 7735
rect 29469 7701 29503 7735
rect 34023 7701 34057 7735
rect 3157 7497 3191 7531
rect 4905 7497 4939 7531
rect 6285 7497 6319 7531
rect 7757 7497 7791 7531
rect 13829 7497 13863 7531
rect 15393 7497 15427 7531
rect 17509 7497 17543 7531
rect 18981 7497 19015 7531
rect 20913 7497 20947 7531
rect 21281 7497 21315 7531
rect 21465 7497 21499 7531
rect 21557 7497 21591 7531
rect 26985 7497 27019 7531
rect 27629 7497 27663 7531
rect 28641 7497 28675 7531
rect 32505 7497 32539 7531
rect 33057 7497 33091 7531
rect 34253 7497 34287 7531
rect 36277 7497 36311 7531
rect 3801 7429 3835 7463
rect 4169 7429 4203 7463
rect 8033 7429 8067 7463
rect 11529 7429 11563 7463
rect 13461 7429 13495 7463
rect 2237 7361 2271 7395
rect 3525 7361 3559 7395
rect 5273 7361 5307 7395
rect 5641 7361 5675 7395
rect 6837 7361 6871 7395
rect 10609 7361 10643 7395
rect 14289 7361 14323 7395
rect 16037 7361 16071 7395
rect 16681 7361 16715 7395
rect 18061 7361 18095 7395
rect 19993 7361 20027 7395
rect 3985 7293 4019 7327
rect 4537 7293 4571 7327
rect 8585 7293 8619 7327
rect 9045 7293 9079 7327
rect 12173 7293 12207 7327
rect 12541 7293 12575 7327
rect 14565 7293 14599 7327
rect 14933 7293 14967 7327
rect 2558 7225 2592 7259
rect 5365 7225 5399 7259
rect 6653 7225 6687 7259
rect 7199 7225 7233 7259
rect 10517 7225 10551 7259
rect 10971 7225 11005 7259
rect 15117 7225 15151 7259
rect 16129 7225 16163 7259
rect 17877 7225 17911 7259
rect 18423 7225 18457 7259
rect 20314 7225 20348 7259
rect 27951 7429 27985 7463
rect 21833 7361 21867 7395
rect 23765 7361 23799 7395
rect 24041 7361 24075 7395
rect 26065 7361 26099 7395
rect 29377 7361 29411 7395
rect 29653 7361 29687 7395
rect 31401 7361 31435 7395
rect 33333 7361 33367 7395
rect 33977 7361 34011 7395
rect 34989 7361 35023 7395
rect 35633 7361 35667 7395
rect 36553 7361 36587 7395
rect 36829 7361 36863 7395
rect 27880 7293 27914 7327
rect 28273 7293 28307 7327
rect 30849 7293 30883 7327
rect 31309 7293 31343 7327
rect 21925 7225 21959 7259
rect 22477 7225 22511 7259
rect 23857 7225 23891 7259
rect 24869 7225 24903 7259
rect 25973 7225 26007 7259
rect 26427 7225 26461 7259
rect 29469 7225 29503 7259
rect 30665 7225 30699 7259
rect 33425 7225 33459 7259
rect 35081 7225 35115 7259
rect 36645 7225 36679 7259
rect 1777 7157 1811 7191
rect 2145 7157 2179 7191
rect 8401 7157 8435 7191
rect 8677 7157 8711 7191
rect 9965 7157 9999 7191
rect 11897 7157 11931 7191
rect 12909 7157 12943 7191
rect 15853 7157 15887 7191
rect 17141 7157 17175 7191
rect 19257 7157 19291 7191
rect 19809 7157 19843 7191
rect 21465 7157 21499 7191
rect 22845 7157 22879 7191
rect 23489 7157 23523 7191
rect 25329 7157 25363 7191
rect 27353 7157 27387 7191
rect 29101 7157 29135 7191
rect 30389 7157 30423 7191
rect 32229 7157 32263 7191
rect 34713 7157 34747 7191
rect 35909 7157 35943 7191
rect 4261 6953 4295 6987
rect 10609 6953 10643 6987
rect 14473 6953 14507 6987
rect 15761 6953 15795 6987
rect 18153 6953 18187 6987
rect 18613 6953 18647 6987
rect 19993 6953 20027 6987
rect 21833 6953 21867 6987
rect 23581 6953 23615 6987
rect 26065 6953 26099 6987
rect 27721 6953 27755 6987
rect 28733 6953 28767 6987
rect 29285 6953 29319 6987
rect 30481 6953 30515 6987
rect 36737 6953 36771 6987
rect 2558 6885 2592 6919
rect 4813 6885 4847 6919
rect 6377 6885 6411 6919
rect 7941 6885 7975 6919
rect 11431 6885 11465 6919
rect 13001 6885 13035 6919
rect 16838 6885 16872 6919
rect 18889 6885 18923 6919
rect 22655 6885 22689 6919
rect 24403 6885 24437 6919
rect 28175 6885 28209 6919
rect 29923 6885 29957 6919
rect 32873 6885 32907 6919
rect 34155 6885 34189 6919
rect 35903 6885 35937 6919
rect 2053 6817 2087 6851
rect 3157 6817 3191 6851
rect 5641 6817 5675 6851
rect 9724 6817 9758 6851
rect 11069 6817 11103 6851
rect 11989 6817 12023 6851
rect 15301 6817 15335 6851
rect 16313 6817 16347 6851
rect 20913 6817 20947 6851
rect 21097 6817 21131 6851
rect 21465 6817 21499 6851
rect 23213 6817 23247 6851
rect 24961 6817 24995 6851
rect 26836 6817 26870 6851
rect 26939 6817 26973 6851
rect 31125 6817 31159 6851
rect 32137 6817 32171 6851
rect 32597 6817 32631 6851
rect 33793 6817 33827 6851
rect 35357 6817 35391 6851
rect 36461 6817 36495 6851
rect 1685 6749 1719 6783
rect 2237 6749 2271 6783
rect 3433 6749 3467 6783
rect 4721 6749 4755 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 6561 6749 6595 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 12909 6749 12943 6783
rect 13185 6749 13219 6783
rect 16497 6749 16531 6783
rect 18797 6749 18831 6783
rect 19441 6749 19475 6783
rect 22293 6749 22327 6783
rect 24041 6749 24075 6783
rect 27813 6749 27847 6783
rect 29561 6749 29595 6783
rect 35541 6749 35575 6783
rect 5273 6681 5307 6715
rect 9137 6681 9171 6715
rect 20361 6681 20395 6715
rect 34713 6681 34747 6715
rect 7297 6613 7331 6647
rect 7665 6613 7699 6647
rect 8861 6613 8895 6647
rect 9827 6613 9861 6647
rect 10149 6613 10183 6647
rect 12541 6613 12575 6647
rect 15485 6613 15519 6647
rect 17417 6613 17451 6647
rect 23857 6613 23891 6647
rect 27261 6613 27295 6647
rect 30849 6613 30883 6647
rect 31493 6613 31527 6647
rect 33333 6613 33367 6647
rect 34989 6613 35023 6647
rect 3617 6409 3651 6443
rect 4353 6409 4387 6443
rect 6561 6409 6595 6443
rect 9137 6409 9171 6443
rect 9597 6409 9631 6443
rect 10793 6409 10827 6443
rect 11161 6409 11195 6443
rect 13461 6409 13495 6443
rect 15761 6409 15795 6443
rect 17141 6409 17175 6443
rect 18521 6409 18555 6443
rect 19717 6409 19751 6443
rect 21281 6409 21315 6443
rect 28089 6409 28123 6443
rect 30941 6409 30975 6443
rect 32137 6409 32171 6443
rect 34253 6409 34287 6443
rect 35909 6409 35943 6443
rect 6193 6341 6227 6375
rect 11529 6341 11563 6375
rect 13093 6341 13127 6375
rect 17509 6341 17543 6375
rect 20085 6341 20119 6375
rect 26801 6341 26835 6375
rect 2053 6273 2087 6307
rect 5273 6273 5307 6307
rect 5917 6273 5951 6307
rect 8217 6273 8251 6307
rect 12541 6273 12575 6307
rect 16221 6273 16255 6307
rect 20361 6273 20395 6307
rect 22385 6273 22419 6307
rect 22937 6273 22971 6307
rect 25237 6273 25271 6307
rect 27353 6273 27387 6307
rect 29009 6273 29043 6307
rect 34989 6273 35023 6307
rect 36829 6273 36863 6307
rect 3868 6205 3902 6239
rect 6904 6205 6938 6239
rect 7297 6205 7331 6239
rect 9689 6205 9723 6239
rect 10149 6205 10183 6239
rect 11345 6205 11379 6239
rect 13921 6205 13955 6239
rect 14105 6205 14139 6239
rect 21833 6205 21867 6239
rect 22293 6205 22327 6239
rect 23673 6205 23707 6239
rect 24225 6205 24259 6239
rect 29285 6205 29319 6239
rect 29745 6205 29779 6239
rect 31125 6205 31159 6239
rect 31585 6205 31619 6239
rect 33977 6205 34011 6239
rect 36277 6205 36311 6239
rect 1961 6137 1995 6171
rect 2415 6137 2449 6171
rect 3341 6137 3375 6171
rect 5365 6137 5399 6171
rect 7757 6137 7791 6171
rect 8309 6137 8343 6171
rect 8861 6137 8895 6171
rect 11897 6137 11931 6171
rect 12633 6137 12667 6171
rect 14013 6137 14047 6171
rect 16129 6137 16163 6171
rect 16583 6137 16617 6171
rect 17877 6137 17911 6171
rect 18797 6137 18831 6171
rect 18889 6137 18923 6171
rect 19441 6137 19475 6171
rect 20453 6137 20487 6171
rect 21005 6137 21039 6171
rect 24409 6137 24443 6171
rect 24777 6137 24811 6171
rect 25145 6137 25179 6171
rect 25599 6137 25633 6171
rect 26525 6137 26559 6171
rect 27077 6137 27111 6171
rect 27169 6137 27203 6171
rect 28457 6137 28491 6171
rect 31861 6137 31895 6171
rect 33333 6137 33367 6171
rect 33425 6137 33459 6171
rect 34621 6137 34655 6171
rect 35081 6137 35115 6171
rect 35633 6137 35667 6171
rect 36553 6137 36587 6171
rect 36645 6137 36679 6171
rect 2973 6069 3007 6103
rect 3939 6069 3973 6103
rect 4629 6069 4663 6103
rect 5089 6069 5123 6103
rect 6975 6069 7009 6103
rect 9781 6069 9815 6103
rect 12173 6069 12207 6103
rect 15393 6069 15427 6103
rect 21649 6069 21683 6103
rect 23397 6069 23431 6103
rect 26157 6069 26191 6103
rect 29377 6069 29411 6103
rect 30389 6069 30423 6103
rect 32505 6069 32539 6103
rect 33149 6069 33183 6103
rect 2881 5865 2915 5899
rect 4997 5865 5031 5899
rect 7481 5865 7515 5899
rect 8861 5865 8895 5899
rect 12449 5865 12483 5899
rect 12817 5865 12851 5899
rect 14657 5865 14691 5899
rect 15577 5865 15611 5899
rect 22385 5865 22419 5899
rect 23765 5865 23799 5899
rect 25237 5865 25271 5899
rect 29653 5865 29687 5899
rect 31217 5865 31251 5899
rect 33057 5865 33091 5899
rect 33701 5865 33735 5899
rect 34805 5865 34839 5899
rect 35081 5865 35115 5899
rect 36645 5865 36679 5899
rect 1777 5797 1811 5831
rect 2282 5797 2316 5831
rect 4439 5797 4473 5831
rect 5641 5797 5675 5831
rect 6285 5797 6319 5831
rect 8027 5797 8061 5831
rect 9873 5797 9907 5831
rect 11891 5797 11925 5831
rect 13461 5797 13495 5831
rect 16313 5797 16347 5831
rect 16767 5797 16801 5831
rect 18797 5797 18831 5831
rect 20269 5797 20303 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 23213 5797 23247 5831
rect 24403 5797 24437 5831
rect 26709 5797 26743 5831
rect 28273 5797 28307 5831
rect 30618 5797 30652 5831
rect 32458 5797 32492 5831
rect 34206 5797 34240 5831
rect 35449 5797 35483 5831
rect 35817 5797 35851 5831
rect 1961 5729 1995 5763
rect 3249 5729 3283 5763
rect 4077 5729 4111 5763
rect 7665 5729 7699 5763
rect 8585 5729 8619 5763
rect 15393 5729 15427 5763
rect 17325 5729 17359 5763
rect 18429 5729 18463 5763
rect 22753 5729 22787 5763
rect 22937 5729 22971 5763
rect 33885 5729 33919 5763
rect 5273 5661 5307 5695
rect 6193 5661 6227 5695
rect 6469 5661 6503 5695
rect 9413 5661 9447 5695
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 11529 5661 11563 5695
rect 13369 5661 13403 5695
rect 15025 5661 15059 5695
rect 16405 5661 16439 5695
rect 17969 5661 18003 5695
rect 18705 5661 18739 5695
rect 18981 5661 19015 5695
rect 21005 5661 21039 5695
rect 24041 5661 24075 5695
rect 26617 5661 26651 5695
rect 27261 5661 27295 5695
rect 28181 5661 28215 5695
rect 28457 5661 28491 5695
rect 29285 5661 29319 5695
rect 30297 5661 30331 5695
rect 32137 5661 32171 5695
rect 35725 5661 35759 5695
rect 36001 5661 36035 5695
rect 13921 5593 13955 5627
rect 22017 5593 22051 5627
rect 24961 5593 24995 5627
rect 10977 5525 11011 5559
rect 11437 5525 11471 5559
rect 14289 5525 14323 5559
rect 15853 5525 15887 5559
rect 17601 5525 17635 5559
rect 19717 5525 19751 5559
rect 20729 5525 20763 5559
rect 1593 5321 1627 5355
rect 2053 5321 2087 5355
rect 4169 5321 4203 5355
rect 5549 5321 5583 5355
rect 6193 5321 6227 5355
rect 7205 5321 7239 5355
rect 8585 5321 8619 5355
rect 8953 5321 8987 5355
rect 10425 5321 10459 5355
rect 13001 5321 13035 5355
rect 15209 5321 15243 5355
rect 16405 5321 16439 5355
rect 17049 5321 17083 5355
rect 22385 5321 22419 5355
rect 24869 5321 24903 5355
rect 26341 5321 26375 5355
rect 28089 5321 28123 5355
rect 28457 5321 28491 5355
rect 33517 5321 33551 5355
rect 34253 5321 34287 5355
rect 35909 5321 35943 5355
rect 2605 5253 2639 5287
rect 12633 5253 12667 5287
rect 13461 5253 13495 5287
rect 18245 5253 18279 5287
rect 22109 5253 22143 5287
rect 26617 5253 26651 5287
rect 26709 5253 26743 5287
rect 32137 5253 32171 5287
rect 33241 5253 33275 5287
rect 36277 5253 36311 5287
rect 2697 5185 2731 5219
rect 4537 5185 4571 5219
rect 4813 5185 4847 5219
rect 6469 5185 6503 5219
rect 7665 5185 7699 5219
rect 12265 5185 12299 5219
rect 13553 5185 13587 5219
rect 14841 5185 14875 5219
rect 15669 5185 15703 5219
rect 21097 5185 21131 5219
rect 21741 5185 21775 5219
rect 25973 5185 26007 5219
rect 1409 5117 1443 5151
rect 9597 5117 9631 5151
rect 9965 5117 9999 5151
rect 10885 5117 10919 5151
rect 11161 5117 11195 5151
rect 12449 5117 12483 5151
rect 16865 5117 16899 5151
rect 18061 5117 18095 5151
rect 18521 5117 18555 5151
rect 19165 5117 19199 5151
rect 19257 5117 19291 5151
rect 23673 5117 23707 5151
rect 26985 5185 27019 5219
rect 27261 5185 27295 5219
rect 29653 5185 29687 5219
rect 31769 5185 31803 5219
rect 32321 5185 32355 5219
rect 34989 5185 35023 5219
rect 35265 5185 35299 5219
rect 36829 5185 36863 5219
rect 30389 5117 30423 5151
rect 30849 5117 30883 5151
rect 31309 5117 31343 5151
rect 3059 5049 3093 5083
rect 4629 5049 4663 5083
rect 7573 5049 7607 5083
rect 8027 5049 8061 5083
rect 9321 5049 9355 5083
rect 10977 5049 11011 5083
rect 11529 5049 11563 5083
rect 13915 5049 13949 5083
rect 15393 5049 15427 5083
rect 15485 5049 15519 5083
rect 19578 5049 19612 5083
rect 21189 5049 21223 5083
rect 23489 5049 23523 5083
rect 24035 5049 24069 5083
rect 25421 5049 25455 5083
rect 26617 5049 26651 5083
rect 27077 5049 27111 5083
rect 29009 5049 29043 5083
rect 29377 5049 29411 5083
rect 29469 5049 29503 5083
rect 32642 5049 32676 5083
rect 33885 5049 33919 5083
rect 35081 5049 35115 5083
rect 36553 5049 36587 5083
rect 36645 5049 36679 5083
rect 3617 4981 3651 5015
rect 9689 4981 9723 5015
rect 11897 4981 11931 5015
rect 14473 4981 14507 5015
rect 17325 4981 17359 5015
rect 17785 4981 17819 5015
rect 20177 4981 20211 5015
rect 20453 4981 20487 5015
rect 20821 4981 20855 5015
rect 22569 4981 22603 5015
rect 23121 4981 23155 5015
rect 24593 4981 24627 5015
rect 30665 4981 30699 5015
rect 31033 4981 31067 5015
rect 34713 4981 34747 5015
rect 1685 4777 1719 4811
rect 3893 4777 3927 4811
rect 5825 4777 5859 4811
rect 12173 4777 12207 4811
rect 12541 4777 12575 4811
rect 14013 4777 14047 4811
rect 19625 4777 19659 4811
rect 21925 4777 21959 4811
rect 24317 4777 24351 4811
rect 24961 4777 24995 4811
rect 26341 4777 26375 4811
rect 29377 4777 29411 4811
rect 32965 4777 32999 4811
rect 34989 4777 35023 4811
rect 36093 4777 36127 4811
rect 36461 4777 36495 4811
rect 2139 4709 2173 4743
rect 4261 4709 4295 4743
rect 5089 4709 5123 4743
rect 8170 4709 8204 4743
rect 9873 4709 9907 4743
rect 10425 4709 10459 4743
rect 11615 4709 11649 4743
rect 12817 4709 12851 4743
rect 13093 4709 13127 4743
rect 13185 4709 13219 4743
rect 14381 4709 14415 4743
rect 19067 4709 19101 4743
rect 19901 4709 19935 4743
rect 20729 4709 20763 4743
rect 21097 4709 21131 4743
rect 21649 4709 21683 4743
rect 24041 4709 24075 4743
rect 24685 4709 24719 4743
rect 26709 4709 26743 4743
rect 28273 4709 28307 4743
rect 31217 4709 31251 4743
rect 33746 4709 33780 4743
rect 35494 4709 35528 4743
rect 6561 4641 6595 4675
rect 6837 4641 6871 4675
rect 7849 4641 7883 4675
rect 8769 4641 8803 4675
rect 15301 4641 15335 4675
rect 15853 4641 15887 4675
rect 16865 4641 16899 4675
rect 18705 4641 18739 4675
rect 20269 4641 20303 4675
rect 23581 4641 23615 4675
rect 23765 4641 23799 4675
rect 24961 4641 24995 4675
rect 25329 4641 25363 4675
rect 30481 4641 30515 4675
rect 30941 4641 30975 4675
rect 1777 4573 1811 4607
rect 3525 4573 3559 4607
rect 4169 4573 4203 4607
rect 4813 4573 4847 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 9781 4573 9815 4607
rect 11253 4573 11287 4607
rect 13461 4573 13495 4607
rect 15669 4573 15703 4607
rect 16405 4573 16439 4607
rect 17233 4573 17267 4607
rect 21005 4573 21039 4607
rect 26617 4573 26651 4607
rect 28181 4573 28215 4607
rect 28825 4573 28859 4607
rect 32137 4573 32171 4607
rect 33425 4573 33459 4607
rect 35173 4573 35207 4607
rect 9413 4505 9447 4539
rect 18061 4505 18095 4539
rect 27169 4505 27203 4539
rect 32597 4505 32631 4539
rect 2697 4437 2731 4471
rect 3065 4437 3099 4471
rect 7757 4437 7791 4471
rect 9045 4437 9079 4471
rect 10793 4437 10827 4471
rect 15117 4437 15151 4471
rect 16681 4437 16715 4471
rect 17003 4437 17037 4471
rect 17141 4437 17175 4471
rect 17325 4437 17359 4471
rect 18429 4437 18463 4471
rect 31493 4437 31527 4471
rect 34345 4437 34379 4471
rect 2421 4233 2455 4267
rect 3985 4233 4019 4267
rect 6377 4233 6411 4267
rect 9229 4233 9263 4267
rect 11897 4233 11931 4267
rect 12817 4233 12851 4267
rect 18199 4233 18233 4267
rect 20913 4233 20947 4267
rect 21281 4233 21315 4267
rect 21649 4233 21683 4267
rect 23397 4233 23431 4267
rect 27629 4233 27663 4267
rect 28181 4233 28215 4267
rect 30481 4233 30515 4267
rect 33701 4233 33735 4267
rect 35909 4233 35943 4267
rect 36277 4233 36311 4267
rect 5641 4165 5675 4199
rect 16589 4165 16623 4199
rect 17325 4165 17359 4199
rect 2697 4097 2731 4131
rect 3341 4097 3375 4131
rect 4537 4097 4571 4131
rect 7849 4097 7883 4131
rect 11345 4097 11379 4131
rect 11529 4097 11563 4131
rect 14749 4097 14783 4131
rect 15761 4097 15795 4131
rect 16460 4097 16494 4131
rect 16681 4097 16715 4131
rect 17785 4097 17819 4131
rect 18429 4097 18463 4131
rect 19441 4097 19475 4131
rect 19993 4097 20027 4131
rect 23029 4097 23063 4131
rect 24501 4097 24535 4131
rect 30941 4097 30975 4131
rect 32413 4097 32447 4131
rect 34621 4097 34655 4131
rect 34989 4097 35023 4131
rect 35265 4097 35299 4131
rect 1660 4029 1694 4063
rect 5733 4029 5767 4063
rect 6837 4029 6871 4063
rect 10701 4029 10735 4063
rect 11253 4029 11287 4063
rect 13185 4029 13219 4063
rect 13553 4029 13587 4063
rect 13829 4029 13863 4063
rect 14289 4029 14323 4063
rect 14933 4029 14967 4063
rect 15117 4029 15151 4063
rect 18291 4029 18325 4063
rect 18797 4029 18831 4063
rect 21833 4029 21867 4063
rect 22201 4029 22235 4063
rect 24961 4029 24995 4063
rect 25881 4029 25915 4063
rect 26709 4029 26743 4063
rect 29561 4029 29595 4063
rect 29929 4029 29963 4063
rect 32597 4029 32631 4063
rect 33057 4029 33091 4063
rect 36461 4029 36495 4063
rect 37013 4029 37047 4063
rect 37600 4029 37634 4063
rect 38025 4029 38059 4063
rect 2145 3961 2179 3995
rect 2789 3961 2823 3995
rect 4261 3961 4295 3995
rect 4353 3961 4387 3995
rect 7757 3961 7791 3995
rect 8211 3961 8245 3995
rect 9597 3961 9631 3995
rect 9965 3961 9999 3995
rect 12265 3961 12299 3995
rect 15485 3961 15519 3995
rect 16313 3961 16347 3995
rect 17049 3961 17083 3995
rect 18061 3961 18095 3995
rect 19165 3961 19199 3995
rect 20314 3961 20348 3995
rect 24869 3961 24903 3995
rect 25323 3961 25357 3995
rect 26617 3961 26651 3995
rect 27071 3961 27105 3995
rect 29101 3961 29135 3995
rect 30113 3961 30147 3995
rect 31125 3961 31159 3995
rect 31217 3961 31251 3995
rect 31769 3961 31803 3995
rect 33333 3961 33367 3995
rect 35081 3961 35115 3995
rect 1731 3893 1765 3927
rect 3709 3893 3743 3927
rect 5273 3893 5307 3927
rect 5917 3893 5951 3927
rect 7021 3893 7055 3927
rect 7389 3893 7423 3927
rect 8769 3893 8803 3927
rect 10241 3893 10275 3927
rect 13553 3893 13587 3927
rect 16129 3893 16163 3927
rect 19809 3893 19843 3927
rect 22017 3893 22051 3927
rect 23673 3893 23707 3927
rect 26249 3893 26283 3927
rect 28457 3893 28491 3927
rect 33977 3893 34011 3927
rect 36645 3893 36679 3927
rect 37703 3893 37737 3927
rect 3249 3689 3283 3723
rect 4169 3689 4203 3723
rect 5181 3689 5215 3723
rect 5733 3689 5767 3723
rect 6837 3689 6871 3723
rect 7573 3689 7607 3723
rect 9045 3689 9079 3723
rect 9873 3689 9907 3723
rect 11069 3689 11103 3723
rect 13461 3689 13495 3723
rect 13921 3689 13955 3723
rect 15025 3689 15059 3723
rect 15577 3689 15611 3723
rect 17877 3689 17911 3723
rect 20177 3689 20211 3723
rect 20545 3689 20579 3723
rect 22201 3689 22235 3723
rect 23305 3689 23339 3723
rect 25145 3689 25179 3723
rect 26249 3689 26283 3723
rect 28089 3689 28123 3723
rect 30113 3689 30147 3723
rect 31125 3689 31159 3723
rect 34621 3689 34655 3723
rect 1955 3621 1989 3655
rect 2881 3621 2915 3655
rect 3893 3621 3927 3655
rect 8217 3621 8251 3655
rect 10517 3621 10551 3655
rect 12817 3621 12851 3655
rect 16405 3621 16439 3655
rect 17233 3621 17267 3655
rect 18245 3621 18279 3655
rect 19901 3621 19935 3655
rect 20913 3621 20947 3655
rect 22747 3621 22781 3655
rect 24225 3621 24259 3655
rect 24317 3621 24351 3655
rect 25973 3621 26007 3655
rect 26801 3621 26835 3655
rect 27353 3621 27387 3655
rect 28543 3621 28577 3655
rect 30526 3621 30560 3655
rect 34022 3621 34056 3655
rect 35633 3621 35667 3655
rect 4077 3553 4111 3587
rect 4629 3553 4663 3587
rect 5825 3553 5859 3587
rect 6193 3553 6227 3587
rect 9689 3553 9723 3587
rect 11069 3553 11103 3587
rect 11345 3553 11379 3587
rect 11621 3553 11655 3587
rect 12964 3553 12998 3587
rect 15669 3553 15703 3587
rect 17380 3553 17414 3587
rect 19073 3553 19107 3587
rect 19441 3553 19475 3587
rect 19625 3553 19659 3587
rect 21097 3553 21131 3587
rect 22385 3553 22419 3587
rect 30205 3553 30239 3587
rect 31401 3553 31435 3587
rect 32229 3553 32263 3587
rect 32597 3553 32631 3587
rect 33701 3553 33735 3587
rect 1593 3485 1627 3519
rect 8125 3485 8159 3519
rect 8769 3485 8803 3519
rect 13185 3485 13219 3519
rect 14197 3485 14231 3519
rect 16037 3485 16071 3519
rect 16865 3485 16899 3519
rect 17601 3485 17635 3519
rect 21465 3485 21499 3519
rect 24501 3485 24535 3519
rect 26709 3485 26743 3519
rect 28181 3485 28215 3519
rect 32873 3485 32907 3519
rect 35173 3485 35207 3519
rect 35541 3485 35575 3519
rect 36001 3485 36035 3519
rect 13093 3417 13127 3451
rect 15945 3417 15979 3451
rect 17509 3417 17543 3451
rect 2513 3349 2547 3383
rect 7941 3349 7975 3383
rect 9505 3349 9539 3383
rect 12541 3349 12575 3383
rect 14565 3349 14599 3383
rect 15807 3349 15841 3383
rect 18613 3349 18647 3383
rect 21833 3349 21867 3383
rect 25513 3349 25547 3383
rect 29101 3349 29135 3383
rect 29469 3349 29503 3383
rect 1685 3145 1719 3179
rect 3709 3145 3743 3179
rect 4077 3145 4111 3179
rect 5089 3145 5123 3179
rect 6285 3145 6319 3179
rect 8125 3145 8159 3179
rect 9873 3145 9907 3179
rect 10517 3145 10551 3179
rect 12173 3145 12207 3179
rect 13461 3145 13495 3179
rect 16589 3145 16623 3179
rect 17233 3145 17267 3179
rect 17785 3145 17819 3179
rect 20913 3145 20947 3179
rect 21281 3145 21315 3179
rect 21833 3145 21867 3179
rect 23489 3145 23523 3179
rect 24225 3145 24259 3179
rect 26065 3145 26099 3179
rect 28089 3145 28123 3179
rect 28733 3145 28767 3179
rect 30297 3145 30331 3179
rect 31953 3145 31987 3179
rect 34069 3145 34103 3179
rect 34713 3145 34747 3179
rect 35909 3145 35943 3179
rect 36277 3145 36311 3179
rect 37611 3145 37645 3179
rect 2789 3077 2823 3111
rect 5273 3077 5307 3111
rect 12541 3077 12575 3111
rect 13921 3077 13955 3111
rect 14105 3077 14139 3111
rect 18153 3077 18187 3111
rect 27169 3077 27203 3111
rect 33701 3077 33735 3111
rect 2237 3009 2271 3043
rect 3157 3009 3191 3043
rect 13093 3009 13127 3043
rect 16037 3009 16071 3043
rect 18521 3009 18555 3043
rect 22753 3009 22787 3043
rect 23765 3009 23799 3043
rect 26341 3009 26375 3043
rect 26617 3009 26651 3043
rect 28319 3009 28353 3043
rect 29653 3009 29687 3043
rect 31585 3009 31619 3043
rect 33149 3009 33183 3043
rect 34989 3009 35023 3043
rect 35265 3009 35299 3043
rect 36461 3009 36495 3043
rect 4169 2941 4203 2975
rect 4629 2941 4663 2975
rect 5181 2941 5215 2975
rect 5457 2941 5491 2975
rect 6837 2941 6871 2975
rect 7297 2941 7331 2975
rect 8493 2941 8527 2975
rect 8953 2941 8987 2975
rect 10241 2941 10275 2975
rect 10701 2941 10735 2975
rect 10793 2941 10827 2975
rect 12449 2941 12483 2975
rect 12725 2941 12759 2975
rect 14013 2941 14047 2975
rect 14289 2941 14323 2975
rect 15577 2941 15611 2975
rect 15669 2941 15703 2975
rect 15853 2941 15887 2975
rect 18061 2941 18095 2975
rect 18337 2941 18371 2975
rect 19901 2941 19935 2975
rect 20085 2941 20119 2975
rect 22017 2941 22051 2975
rect 22569 2941 22603 2975
rect 24777 2941 24811 2975
rect 28216 2941 28250 2975
rect 30757 2941 30791 2975
rect 30849 2941 30883 2975
rect 31401 2941 31435 2975
rect 32321 2941 32355 2975
rect 32413 2941 32447 2975
rect 32873 2941 32907 2975
rect 37508 2941 37542 2975
rect 37933 2941 37967 2975
rect 2329 2873 2363 2907
rect 5917 2873 5951 2907
rect 8769 2873 8803 2907
rect 9274 2873 9308 2907
rect 11805 2873 11839 2907
rect 15393 2873 15427 2907
rect 19165 2873 19199 2907
rect 19533 2873 19567 2907
rect 23121 2873 23155 2907
rect 24685 2873 24719 2907
rect 25098 2873 25132 2907
rect 26709 2873 26743 2907
rect 29101 2873 29135 2907
rect 29377 2873 29411 2907
rect 29469 2873 29503 2907
rect 35081 2873 35115 2907
rect 2053 2805 2087 2839
rect 4353 2805 4387 2839
rect 6561 2805 6595 2839
rect 6929 2805 6963 2839
rect 14473 2805 14507 2839
rect 15025 2805 15059 2839
rect 19717 2805 19751 2839
rect 25697 2805 25731 2839
rect 27537 2805 27571 2839
rect 1685 2601 1719 2635
rect 2053 2601 2087 2635
rect 5365 2601 5399 2635
rect 6285 2601 6319 2635
rect 7113 2601 7147 2635
rect 9137 2601 9171 2635
rect 9505 2601 9539 2635
rect 10885 2601 10919 2635
rect 13277 2601 13311 2635
rect 14013 2601 14047 2635
rect 15209 2601 15243 2635
rect 16589 2601 16623 2635
rect 16957 2601 16991 2635
rect 17509 2601 17543 2635
rect 18061 2601 18095 2635
rect 19717 2601 19751 2635
rect 20913 2601 20947 2635
rect 21373 2601 21407 2635
rect 23397 2601 23431 2635
rect 23765 2601 23799 2635
rect 25421 2601 25455 2635
rect 26341 2601 26375 2635
rect 27261 2601 27295 2635
rect 28825 2601 28859 2635
rect 29469 2601 29503 2635
rect 30941 2601 30975 2635
rect 32597 2601 32631 2635
rect 33057 2601 33091 2635
rect 34069 2601 34103 2635
rect 34989 2601 35023 2635
rect 36001 2601 36035 2635
rect 2329 2533 2363 2567
rect 2881 2533 2915 2567
rect 4445 2533 4479 2567
rect 7941 2533 7975 2567
rect 8861 2533 8895 2567
rect 9965 2533 9999 2567
rect 10517 2533 10551 2567
rect 11161 2533 11195 2567
rect 12633 2533 12667 2567
rect 18337 2533 18371 2567
rect 20637 2533 20671 2567
rect 23121 2533 23155 2567
rect 25053 2533 25087 2567
rect 28181 2533 28215 2567
rect 32229 2533 32263 2567
rect 4905 2465 4939 2499
rect 5181 2465 5215 2499
rect 6009 2465 6043 2499
rect 6745 2465 6779 2499
rect 6929 2465 6963 2499
rect 7665 2465 7699 2499
rect 8401 2465 8435 2499
rect 8585 2465 8619 2499
rect 11380 2465 11414 2499
rect 13645 2465 13679 2499
rect 14197 2465 14231 2499
rect 15577 2465 15611 2499
rect 17049 2465 17083 2499
rect 18429 2465 18463 2499
rect 19901 2465 19935 2499
rect 21189 2465 21223 2499
rect 22661 2465 22695 2499
rect 22937 2465 22971 2499
rect 24041 2465 24075 2499
rect 24501 2465 24535 2499
rect 25640 2465 25674 2499
rect 26709 2465 26743 2499
rect 27721 2465 27755 2499
rect 27905 2465 27939 2499
rect 29745 2465 29779 2499
rect 30205 2465 30239 2499
rect 31344 2465 31378 2499
rect 31769 2465 31803 2499
rect 33676 2465 33710 2499
rect 35516 2465 35550 2499
rect 36496 2465 36530 2499
rect 36921 2465 36955 2499
rect 2237 2397 2271 2431
rect 3157 2397 3191 2431
rect 4997 2397 5031 2431
rect 9873 2397 9907 2431
rect 11483 2397 11517 2431
rect 12780 2397 12814 2431
rect 13001 2397 13035 2431
rect 15485 2397 15519 2431
rect 21741 2397 21775 2431
rect 22109 2397 22143 2431
rect 24685 2397 24719 2431
rect 29193 2397 29227 2431
rect 30297 2397 30331 2431
rect 36599 2397 36633 2431
rect 12081 2329 12115 2363
rect 14381 2329 14415 2363
rect 17233 2329 17267 2363
rect 35587 2329 35621 2363
rect 4721 2261 4755 2295
rect 12449 2261 12483 2295
rect 12909 2261 12943 2295
rect 14841 2261 14875 2295
rect 20085 2261 20119 2295
rect 25743 2261 25777 2295
rect 31447 2261 31481 2295
rect 33747 2261 33781 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 35618 12968 35624 12980
rect 35579 12940 35624 12968
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 2568 12767 2626 12773
rect 2568 12733 2580 12767
rect 2614 12764 2626 12767
rect 2777 12767 2835 12773
rect 2777 12764 2789 12767
rect 2614 12736 2789 12764
rect 2614 12733 2626 12736
rect 2568 12727 2626 12733
rect 2777 12733 2789 12736
rect 2823 12733 2835 12767
rect 2777 12727 2835 12733
rect 4960 12767 5018 12773
rect 4960 12733 4972 12767
rect 5006 12764 5018 12767
rect 5442 12764 5448 12776
rect 5006 12736 5448 12764
rect 5006 12733 5018 12736
rect 4960 12727 5018 12733
rect 1412 12696 1440 12727
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 35434 12764 35440 12776
rect 13035 12736 13584 12764
rect 35347 12736 35440 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 2041 12699 2099 12705
rect 2041 12696 2053 12699
rect 1412 12668 2053 12696
rect 2041 12665 2053 12668
rect 2087 12696 2099 12699
rect 11330 12696 11336 12708
rect 2087 12668 11336 12696
rect 2087 12665 2099 12668
rect 2041 12659 2099 12665
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2639 12631 2697 12637
rect 2639 12628 2651 12631
rect 2004 12600 2651 12628
rect 2004 12588 2010 12600
rect 2639 12597 2651 12600
rect 2685 12597 2697 12631
rect 2639 12591 2697 12597
rect 2777 12631 2835 12637
rect 2777 12597 2789 12631
rect 2823 12628 2835 12631
rect 3053 12631 3111 12637
rect 3053 12628 3065 12631
rect 2823 12600 3065 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3053 12597 3065 12600
rect 3099 12628 3111 12631
rect 3694 12628 3700 12640
rect 3099 12600 3700 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 5031 12631 5089 12637
rect 5031 12597 5043 12631
rect 5077 12628 5089 12631
rect 5258 12628 5264 12640
rect 5077 12600 5264 12628
rect 5077 12597 5089 12600
rect 5031 12591 5089 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5442 12628 5448 12640
rect 5403 12600 5448 12628
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 13170 12628 13176 12640
rect 13131 12600 13176 12628
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 13556 12637 13584 12736
rect 35434 12724 35440 12736
rect 35492 12764 35498 12776
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35492 12736 36001 12764
rect 35492 12724 35498 12736
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 13541 12631 13599 12637
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 18414 12628 18420 12640
rect 13587 12600 18420 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1486 12384 1492 12436
rect 1544 12424 1550 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1544 12396 1593 12424
rect 1544 12384 1550 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1670 12288 1676 12300
rect 1443 12260 1676 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12288 2559 12291
rect 2866 12288 2872 12300
rect 2547 12260 2872 12288
rect 2547 12257 2559 12260
rect 2501 12251 2559 12257
rect 2866 12248 2872 12260
rect 2924 12288 2930 12300
rect 3970 12288 3976 12300
rect 2924 12260 3976 12288
rect 2924 12248 2930 12260
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 4132 12291 4190 12297
rect 4132 12257 4144 12291
rect 4178 12288 4190 12291
rect 4246 12288 4252 12300
rect 4178 12260 4252 12288
rect 4178 12257 4190 12260
rect 4132 12251 4190 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 5902 12248 5908 12300
rect 5960 12297 5966 12300
rect 5960 12291 5998 12297
rect 5986 12257 5998 12291
rect 5960 12251 5998 12257
rect 5960 12248 5966 12251
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 11330 12297 11336 12300
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 10100 12260 10241 12288
rect 10100 12248 10106 12260
rect 10229 12257 10241 12260
rect 10275 12257 10287 12291
rect 10229 12251 10287 12257
rect 11308 12291 11336 12297
rect 11308 12257 11320 12291
rect 11388 12288 11394 12300
rect 12158 12288 12164 12300
rect 11388 12260 12164 12288
rect 11308 12251 11336 12257
rect 11330 12248 11336 12251
rect 11388 12248 11394 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13446 12288 13452 12300
rect 13127 12260 13452 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 2038 12084 2044 12096
rect 1999 12056 2044 12084
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 2406 12084 2412 12096
rect 2367 12056 2412 12084
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 2682 12084 2688 12096
rect 2643 12056 2688 12084
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 4154 12044 4160 12096
rect 4212 12093 4218 12096
rect 4212 12087 4261 12093
rect 4212 12053 4215 12087
rect 4249 12053 4261 12087
rect 4212 12047 4261 12053
rect 6043 12087 6101 12093
rect 6043 12053 6055 12087
rect 6089 12084 6101 12087
rect 6730 12084 6736 12096
rect 6089 12056 6736 12084
rect 6089 12053 6101 12056
rect 6043 12047 6101 12053
rect 4212 12044 4218 12047
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 10410 12084 10416 12096
rect 10371 12056 10416 12084
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 11379 12087 11437 12093
rect 11379 12053 11391 12087
rect 11425 12084 11437 12087
rect 11790 12084 11796 12096
rect 11425 12056 11796 12084
rect 11425 12053 11437 12056
rect 11379 12047 11437 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13998 12084 14004 12096
rect 13311 12056 14004 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 14274 12084 14280 12096
rect 14235 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 14826 11744 14832 11756
rect 14292 11716 14832 11744
rect 14292 11688 14320 11716
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 2038 11676 2044 11688
rect 1999 11648 2044 11676
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2406 11676 2412 11688
rect 2367 11648 2412 11676
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3344 11648 3433 11676
rect 2590 11608 2596 11620
rect 2551 11580 2596 11608
rect 2590 11568 2596 11580
rect 2648 11568 2654 11620
rect 3344 11552 3372 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 4890 11636 4896 11688
rect 4948 11685 4954 11688
rect 4948 11679 4986 11685
rect 4974 11676 4986 11679
rect 5353 11679 5411 11685
rect 5353 11676 5365 11679
rect 4974 11648 5365 11676
rect 4974 11645 4986 11648
rect 4948 11639 4986 11645
rect 5353 11645 5365 11648
rect 5399 11645 5411 11679
rect 5353 11639 5411 11645
rect 6892 11679 6950 11685
rect 6892 11645 6904 11679
rect 6938 11676 6950 11679
rect 7006 11676 7012 11688
rect 6938 11648 7012 11676
rect 6938 11645 6950 11648
rect 6892 11639 6950 11645
rect 4948 11636 4954 11639
rect 7006 11636 7012 11648
rect 7064 11676 7070 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 7064 11648 7297 11676
rect 7064 11636 7070 11648
rect 7285 11645 7297 11648
rect 7331 11676 7343 11679
rect 8110 11676 8116 11688
rect 7331 11648 8116 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10502 11676 10508 11688
rect 10275 11648 10508 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10560 11648 11069 11676
rect 10560 11636 10566 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11238 11636 11244 11688
rect 11296 11685 11302 11688
rect 11296 11679 11334 11685
rect 11322 11676 11334 11679
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11322 11648 11713 11676
rect 11322 11645 11334 11648
rect 11296 11639 11334 11645
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 14274 11676 14280 11688
rect 14235 11648 14280 11676
rect 11701 11639 11759 11645
rect 11296 11636 11302 11639
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14737 11679 14795 11685
rect 14737 11645 14749 11679
rect 14783 11645 14795 11679
rect 14737 11639 14795 11645
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4246 11608 4252 11620
rect 4203 11580 4252 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4246 11568 4252 11580
rect 4304 11608 4310 11620
rect 5442 11608 5448 11620
rect 4304 11580 5448 11608
rect 4304 11568 4310 11580
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 10042 11568 10048 11620
rect 10100 11608 10106 11620
rect 10689 11611 10747 11617
rect 10689 11608 10701 11611
rect 10100 11580 10701 11608
rect 10100 11568 10106 11580
rect 10689 11577 10701 11580
rect 10735 11577 10747 11611
rect 14752 11608 14780 11639
rect 18322 11636 18328 11688
rect 18380 11676 18386 11688
rect 18452 11679 18510 11685
rect 18452 11676 18464 11679
rect 18380 11648 18464 11676
rect 18380 11636 18386 11648
rect 18452 11645 18464 11648
rect 18498 11676 18510 11679
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18498 11648 18889 11676
rect 18498 11645 18510 11648
rect 18452 11639 18510 11645
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 19740 11679 19798 11685
rect 19740 11676 19752 11679
rect 19484 11648 19752 11676
rect 19484 11636 19490 11648
rect 19740 11645 19752 11648
rect 19786 11676 19798 11679
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 19786 11648 20177 11676
rect 19786 11645 19798 11648
rect 19740 11639 19798 11645
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 15010 11608 15016 11620
rect 10689 11571 10747 11577
rect 14108 11580 14780 11608
rect 14971 11580 15016 11608
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 3326 11540 3332 11552
rect 3287 11512 3332 11540
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 3602 11540 3608 11552
rect 3563 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 4982 11500 4988 11552
rect 5040 11549 5046 11552
rect 5040 11543 5089 11549
rect 5040 11509 5043 11543
rect 5077 11509 5089 11543
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5040 11503 5089 11509
rect 5040 11500 5046 11503
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6914 11500 6920 11552
rect 6972 11549 6978 11552
rect 6972 11543 7021 11549
rect 6972 11509 6975 11543
rect 7009 11509 7021 11543
rect 10410 11540 10416 11552
rect 10371 11512 10416 11540
rect 6972 11503 7021 11509
rect 6972 11500 6978 11503
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11422 11549 11428 11552
rect 11379 11543 11428 11549
rect 11379 11509 11391 11543
rect 11425 11509 11428 11543
rect 11379 11503 11428 11509
rect 11422 11500 11428 11503
rect 11480 11500 11486 11552
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12710 11540 12716 11552
rect 12483 11512 12716 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13446 11540 13452 11552
rect 13219 11512 13452 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 14108 11549 14136 11580
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 14056 11512 14105 11540
rect 14056 11500 14062 11512
rect 14093 11509 14105 11512
rect 14139 11509 14151 11543
rect 14093 11503 14151 11509
rect 18555 11543 18613 11549
rect 18555 11509 18567 11543
rect 18601 11540 18613 11543
rect 18782 11540 18788 11552
rect 18601 11512 18788 11540
rect 18601 11509 18613 11512
rect 18555 11503 18613 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19843 11543 19901 11549
rect 19843 11509 19855 11543
rect 19889 11540 19901 11543
rect 20070 11540 20076 11552
rect 19889 11512 20076 11540
rect 19889 11509 19901 11512
rect 19843 11503 19901 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 17034 11345 17040 11348
rect 16991 11339 17040 11345
rect 16991 11305 17003 11339
rect 17037 11305 17040 11339
rect 16991 11299 17040 11305
rect 17034 11296 17040 11299
rect 17092 11296 17098 11348
rect 35618 11336 35624 11348
rect 35579 11308 35624 11336
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 4132 11203 4190 11209
rect 4132 11169 4144 11203
rect 4178 11200 4190 11203
rect 4246 11200 4252 11212
rect 4178 11172 4252 11200
rect 4178 11169 4190 11172
rect 4132 11163 4190 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 5166 11209 5172 11212
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5144 11203 5172 11209
rect 5144 11200 5156 11203
rect 4663 11172 5156 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 5144 11169 5156 11172
rect 5144 11163 5172 11169
rect 5166 11160 5172 11163
rect 5224 11160 5230 11212
rect 6178 11209 6184 11212
rect 6156 11203 6184 11209
rect 6156 11169 6168 11203
rect 6156 11163 6184 11169
rect 6178 11160 6184 11163
rect 6236 11160 6242 11212
rect 7098 11160 7104 11212
rect 7156 11209 7162 11212
rect 8202 11209 8208 11212
rect 7156 11203 7194 11209
rect 7182 11169 7194 11203
rect 7156 11163 7194 11169
rect 8180 11203 8208 11209
rect 8180 11169 8192 11203
rect 8180 11163 8208 11169
rect 7156 11160 7162 11163
rect 8202 11160 8208 11163
rect 8260 11160 8266 11212
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 10756 11203 10814 11209
rect 10756 11169 10768 11203
rect 10802 11200 10814 11203
rect 10802 11169 10824 11200
rect 10756 11163 10824 11169
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2280 11104 2329 11132
rect 2280 11092 2286 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10796 11132 10824 11163
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11756 11172 11805 11200
rect 11756 11160 11762 11172
rect 11793 11169 11805 11172
rect 11839 11169 11851 11203
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 11793 11163 11851 11169
rect 13464 11172 13645 11200
rect 9640 11104 11100 11132
rect 9640 11092 9646 11104
rect 4203 11067 4261 11073
rect 4203 11064 4215 11067
rect 4080 11036 4215 11064
rect 1765 10999 1823 11005
rect 1765 10965 1777 10999
rect 1811 10996 1823 10999
rect 1854 10996 1860 11008
rect 1811 10968 1860 10996
rect 1811 10965 1823 10968
rect 1765 10959 1823 10965
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 4080 10996 4108 11036
rect 4203 11033 4215 11036
rect 4249 11033 4261 11067
rect 4203 11027 4261 11033
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 5215 11067 5273 11073
rect 5215 11064 5227 11067
rect 4764 11036 5227 11064
rect 4764 11024 4770 11036
rect 5215 11033 5227 11036
rect 5261 11033 5273 11067
rect 5215 11027 5273 11033
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 6227 11067 6285 11073
rect 6227 11064 6239 11067
rect 5500 11036 6239 11064
rect 5500 11024 5506 11036
rect 6227 11033 6239 11036
rect 6273 11033 6285 11067
rect 6227 11027 6285 11033
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 7239 11067 7297 11073
rect 7239 11064 7251 11067
rect 6420 11036 7251 11064
rect 6420 11024 6426 11036
rect 7239 11033 7251 11036
rect 7285 11033 7297 11067
rect 9858 11064 9864 11076
rect 9819 11036 9864 11064
rect 7239 11027 7297 11033
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 10827 11067 10885 11073
rect 10827 11033 10839 11067
rect 10873 11064 10885 11067
rect 10962 11064 10968 11076
rect 10873 11036 10968 11064
rect 10873 11033 10885 11036
rect 10827 11027 10885 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 3568 10968 4108 10996
rect 3568 10956 3574 10968
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 8251 10999 8309 11005
rect 8251 10996 8263 10999
rect 7524 10968 8263 10996
rect 7524 10956 7530 10968
rect 8251 10965 8263 10968
rect 8297 10965 8309 10999
rect 11072 10996 11100 11104
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12492 11104 12537 11132
rect 12492 11092 12498 11104
rect 11238 10996 11244 11008
rect 11072 10968 11244 10996
rect 8251 10959 8309 10965
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13464 11005 13492 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 14056 11172 14105 11200
rect 14056 11160 14062 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 18506 11209 18512 11212
rect 16888 11203 16946 11209
rect 16888 11200 16900 11203
rect 16724 11172 16900 11200
rect 16724 11160 16730 11172
rect 16888 11169 16900 11172
rect 16934 11169 16946 11203
rect 16888 11163 16946 11169
rect 18484 11203 18512 11209
rect 18484 11169 18496 11203
rect 18484 11163 18512 11169
rect 18506 11160 18512 11163
rect 18564 11160 18570 11212
rect 19518 11209 19524 11212
rect 19496 11203 19524 11209
rect 19496 11169 19508 11203
rect 19496 11163 19524 11169
rect 19518 11160 19524 11163
rect 19576 11160 19582 11212
rect 22094 11209 22100 11212
rect 22072 11203 22100 11209
rect 22072 11169 22084 11203
rect 22072 11163 22100 11169
rect 22094 11160 22100 11163
rect 22152 11160 22158 11212
rect 26602 11160 26608 11212
rect 26660 11209 26666 11212
rect 26660 11203 26698 11209
rect 26686 11169 26698 11203
rect 26660 11163 26698 11169
rect 26660 11160 26666 11163
rect 34146 11160 34152 11212
rect 34204 11200 34210 11212
rect 34368 11203 34426 11209
rect 34368 11200 34380 11203
rect 34204 11172 34380 11200
rect 34204 11160 34210 11172
rect 34368 11169 34380 11172
rect 34414 11169 34426 11203
rect 34368 11163 34426 11169
rect 35250 11160 35256 11212
rect 35308 11200 35314 11212
rect 35437 11203 35495 11209
rect 35437 11200 35449 11203
rect 35308 11172 35449 11200
rect 35308 11160 35314 11172
rect 35437 11169 35449 11172
rect 35483 11169 35495 11203
rect 35437 11163 35495 11169
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 14918 11132 14924 11144
rect 14415 11104 14924 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15654 11132 15660 11144
rect 15615 11104 15660 11132
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 18598 11073 18604 11076
rect 18555 11067 18604 11073
rect 18555 11033 18567 11067
rect 18601 11033 18604 11067
rect 18555 11027 18604 11033
rect 18598 11024 18604 11027
rect 18656 11024 18662 11076
rect 19610 11073 19616 11076
rect 19567 11067 19616 11073
rect 19567 11033 19579 11067
rect 19613 11033 19616 11067
rect 19567 11027 19616 11033
rect 19610 11024 19616 11027
rect 19668 11024 19674 11076
rect 22143 11067 22201 11073
rect 22143 11033 22155 11067
rect 22189 11064 22201 11067
rect 24302 11064 24308 11076
rect 22189 11036 24308 11064
rect 22189 11033 22201 11036
rect 22143 11027 22201 11033
rect 24302 11024 24308 11036
rect 24360 11024 24366 11076
rect 26743 11067 26801 11073
rect 26743 11033 26755 11067
rect 26789 11064 26801 11067
rect 27522 11064 27528 11076
rect 26789 11036 27528 11064
rect 26789 11033 26801 11036
rect 26743 11027 26801 11033
rect 27522 11024 27528 11036
rect 27580 11024 27586 11076
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 13412 10968 13461 10996
rect 13412 10956 13418 10968
rect 13449 10965 13461 10968
rect 13495 10965 13507 10999
rect 13449 10959 13507 10965
rect 34054 10956 34060 11008
rect 34112 10996 34118 11008
rect 34471 10999 34529 11005
rect 34471 10996 34483 10999
rect 34112 10968 34483 10996
rect 34112 10956 34118 10968
rect 34471 10965 34483 10968
rect 34517 10965 34529 10999
rect 34471 10959 34529 10965
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1452 10764 1593 10792
rect 1452 10752 1458 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4120 10764 4537 10792
rect 4120 10752 4126 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 5859 10795 5917 10801
rect 5859 10761 5871 10795
rect 5905 10792 5917 10795
rect 6638 10792 6644 10804
rect 5905 10764 6644 10792
rect 5905 10761 5917 10764
rect 5859 10755 5917 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7156 10764 7481 10792
rect 7156 10752 7162 10764
rect 7469 10761 7481 10764
rect 7515 10792 7527 10795
rect 8018 10792 8024 10804
rect 7515 10764 8024 10792
rect 7515 10761 7527 10764
rect 7469 10755 7527 10761
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 8352 10764 8585 10792
rect 8352 10752 8358 10764
rect 8573 10761 8585 10764
rect 8619 10792 8631 10795
rect 9582 10792 9588 10804
rect 8619 10764 9588 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 18506 10792 18512 10804
rect 18467 10764 18512 10792
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 26234 10792 26240 10804
rect 26195 10764 26240 10792
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 35618 10792 35624 10804
rect 35579 10764 35624 10792
rect 35618 10752 35624 10764
rect 35676 10752 35682 10804
rect 2038 10684 2044 10736
rect 2096 10724 2102 10736
rect 2593 10727 2651 10733
rect 2593 10724 2605 10727
rect 2096 10696 2605 10724
rect 2096 10684 2102 10696
rect 2593 10693 2605 10696
rect 2639 10693 2651 10727
rect 2593 10687 2651 10693
rect 2608 10656 2636 10687
rect 2608 10628 3372 10656
rect 3344 10600 3372 10628
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4157 10659 4215 10665
rect 4157 10656 4169 10659
rect 4120 10628 4169 10656
rect 4120 10616 4126 10628
rect 4157 10625 4169 10628
rect 4203 10656 4215 10659
rect 4246 10656 4252 10668
rect 4203 10628 4252 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 13633 10659 13691 10665
rect 13633 10656 13645 10659
rect 11572 10628 13645 10656
rect 11572 10616 11578 10628
rect 13633 10625 13645 10628
rect 13679 10656 13691 10659
rect 13998 10656 14004 10668
rect 13679 10628 14004 10656
rect 13679 10625 13691 10628
rect 13633 10619 13691 10625
rect 13998 10616 14004 10628
rect 14056 10656 14062 10668
rect 15749 10659 15807 10665
rect 14056 10628 14596 10656
rect 14056 10616 14062 10628
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1443 10560 2084 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2056 10464 2084 10560
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 2777 10591 2835 10597
rect 2777 10588 2789 10591
rect 2556 10560 2789 10588
rect 2556 10548 2562 10560
rect 2777 10557 2789 10560
rect 2823 10557 2835 10591
rect 3326 10588 3332 10600
rect 3287 10560 3332 10588
rect 2777 10551 2835 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 5166 10588 5172 10600
rect 4387 10560 5172 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5810 10597 5816 10600
rect 5788 10591 5816 10597
rect 5788 10557 5800 10591
rect 5868 10588 5874 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 5868 10560 6561 10588
rect 5788 10551 5816 10557
rect 5810 10548 5816 10551
rect 5868 10548 5874 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 8067 10560 8677 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8665 10557 8677 10560
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 10318 10548 10324 10600
rect 10376 10597 10382 10600
rect 10376 10591 10414 10597
rect 10402 10588 10414 10591
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10402 10560 10793 10588
rect 10402 10557 10414 10560
rect 10376 10551 10414 10557
rect 10781 10557 10793 10560
rect 10827 10588 10839 10591
rect 11368 10591 11426 10597
rect 11368 10588 11380 10591
rect 10827 10560 11380 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11368 10557 11380 10560
rect 11414 10588 11426 10591
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11414 10560 11805 10588
rect 11414 10557 11426 10560
rect 11368 10551 11426 10557
rect 11793 10557 11805 10560
rect 11839 10588 11851 10591
rect 11882 10588 11888 10600
rect 11839 10560 11888 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 10376 10548 10382 10551
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12299 10560 12541 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12529 10557 12541 10560
rect 12575 10588 12587 10591
rect 12986 10588 12992 10600
rect 12575 10560 12992 10588
rect 12575 10557 12587 10560
rect 12529 10551 12587 10557
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 14090 10588 14096 10600
rect 14051 10560 14096 10588
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 14568 10597 14596 10628
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 19518 10656 19524 10668
rect 15795 10628 16344 10656
rect 19479 10628 19524 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16316 10600 16344 10628
rect 19518 10616 19524 10628
rect 19576 10656 19582 10668
rect 26252 10656 26280 10752
rect 19576 10628 21404 10656
rect 19576 10616 19582 10628
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15841 10591 15899 10597
rect 15841 10588 15853 10591
rect 15344 10560 15853 10588
rect 15344 10548 15350 10560
rect 15841 10557 15853 10560
rect 15887 10557 15899 10591
rect 16298 10588 16304 10600
rect 16259 10560 16304 10588
rect 15841 10551 15899 10557
rect 3513 10523 3571 10529
rect 3513 10489 3525 10523
rect 3559 10520 3571 10523
rect 3970 10520 3976 10532
rect 3559 10492 3976 10520
rect 3559 10489 3571 10492
rect 3513 10483 3571 10489
rect 3970 10480 3976 10492
rect 4028 10480 4034 10532
rect 8570 10480 8576 10532
rect 8628 10520 8634 10532
rect 9309 10523 9367 10529
rect 9309 10520 9321 10523
rect 8628 10492 9321 10520
rect 8628 10480 8634 10492
rect 9309 10489 9321 10492
rect 9355 10489 9367 10523
rect 9309 10483 9367 10489
rect 11471 10523 11529 10529
rect 11471 10489 11483 10523
rect 11517 10520 11529 10523
rect 12066 10520 12072 10532
rect 11517 10492 12072 10520
rect 11517 10489 11529 10492
rect 11471 10483 11529 10489
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 14829 10523 14887 10529
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 15102 10520 15108 10532
rect 14875 10492 15108 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 15856 10520 15884 10551
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 18046 10548 18052 10600
rect 18104 10597 18110 10600
rect 18104 10591 18142 10597
rect 18130 10588 18142 10591
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18130 10560 18889 10588
rect 18130 10557 18142 10560
rect 18104 10551 18142 10557
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 18104 10548 18110 10551
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19096 10591 19154 10597
rect 19096 10588 19108 10591
rect 19024 10560 19108 10588
rect 19024 10548 19030 10560
rect 19096 10557 19108 10560
rect 19142 10588 19154 10591
rect 19889 10591 19947 10597
rect 19889 10588 19901 10591
rect 19142 10560 19901 10588
rect 19142 10557 19154 10560
rect 19096 10551 19154 10557
rect 19889 10557 19901 10560
rect 19935 10588 19947 10591
rect 19978 10588 19984 10600
rect 19935 10560 19984 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 20844 10591 20902 10597
rect 20844 10588 20856 10591
rect 20772 10560 20856 10588
rect 20772 10548 20778 10560
rect 20844 10557 20856 10560
rect 20890 10588 20902 10591
rect 21269 10591 21327 10597
rect 21269 10588 21281 10591
rect 20890 10560 21281 10588
rect 20890 10557 20902 10560
rect 20844 10551 20902 10557
rect 21269 10557 21281 10560
rect 21315 10557 21327 10591
rect 21376 10588 21404 10628
rect 25700 10628 26280 10656
rect 25700 10600 25728 10628
rect 21856 10591 21914 10597
rect 21856 10588 21868 10591
rect 21376 10560 21868 10588
rect 21269 10551 21327 10557
rect 21856 10557 21868 10560
rect 21902 10588 21914 10591
rect 22370 10588 22376 10600
rect 21902 10560 22376 10588
rect 21902 10557 21914 10560
rect 21856 10551 21914 10557
rect 16482 10520 16488 10532
rect 15856 10492 16488 10520
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 5166 10452 5172 10464
rect 5127 10424 5172 10452
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 7282 10452 7288 10464
rect 7055 10424 7288 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8665 10455 8723 10461
rect 8665 10421 8677 10455
rect 8711 10452 8723 10455
rect 8941 10455 8999 10461
rect 8941 10452 8953 10455
rect 8711 10424 8953 10452
rect 8711 10421 8723 10424
rect 8665 10415 8723 10421
rect 8941 10421 8953 10424
rect 8987 10452 8999 10455
rect 9398 10452 9404 10464
rect 8987 10424 9404 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 9766 10452 9772 10464
rect 9727 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10459 10455 10517 10461
rect 10459 10421 10471 10455
rect 10505 10452 10517 10455
rect 10686 10452 10692 10464
rect 10505 10424 10692 10452
rect 10505 10421 10517 10424
rect 10459 10415 10517 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11238 10452 11244 10464
rect 11199 10424 11244 10452
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16206 10452 16212 10464
rect 16163 10424 16212 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16724 10424 16865 10452
rect 16724 10412 16730 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18187 10455 18245 10461
rect 18187 10452 18199 10455
rect 17920 10424 18199 10452
rect 17920 10412 17926 10424
rect 18187 10421 18199 10424
rect 18233 10421 18245 10455
rect 18187 10415 18245 10421
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19199 10455 19257 10461
rect 19199 10452 19211 10455
rect 19116 10424 19211 10452
rect 19116 10412 19122 10424
rect 19199 10421 19211 10424
rect 19245 10421 19257 10455
rect 19199 10415 19257 10421
rect 20714 10412 20720 10464
rect 20772 10452 20778 10464
rect 20947 10455 21005 10461
rect 20947 10452 20959 10455
rect 20772 10424 20959 10452
rect 20772 10412 20778 10424
rect 20947 10421 20959 10424
rect 20993 10421 21005 10455
rect 21284 10452 21312 10551
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 25682 10588 25688 10600
rect 25740 10597 25746 10600
rect 25740 10591 25778 10597
rect 25595 10560 25688 10588
rect 25682 10548 25688 10560
rect 25766 10557 25778 10591
rect 25740 10551 25778 10557
rect 25823 10591 25881 10597
rect 25823 10557 25835 10591
rect 25869 10588 25881 10591
rect 26142 10588 26148 10600
rect 25869 10560 26148 10588
rect 25869 10557 25881 10560
rect 25823 10551 25881 10557
rect 25740 10548 25746 10551
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 26694 10548 26700 10600
rect 26752 10597 26758 10600
rect 26752 10591 26790 10597
rect 26778 10588 26790 10591
rect 27154 10588 27160 10600
rect 26778 10560 27160 10588
rect 26778 10557 26790 10560
rect 26752 10551 26790 10557
rect 26752 10548 26758 10551
rect 27154 10548 27160 10560
rect 27212 10548 27218 10600
rect 27776 10591 27834 10597
rect 27776 10557 27788 10591
rect 27822 10588 27834 10591
rect 28166 10588 28172 10600
rect 27822 10560 28172 10588
rect 27822 10557 27834 10560
rect 27776 10551 27834 10557
rect 28166 10548 28172 10560
rect 28224 10548 28230 10600
rect 33296 10591 33354 10597
rect 33296 10557 33308 10591
rect 33342 10588 33354 10591
rect 33342 10557 33364 10588
rect 33296 10551 33364 10557
rect 21726 10480 21732 10532
rect 21784 10520 21790 10532
rect 22094 10520 22100 10532
rect 21784 10492 22100 10520
rect 21784 10480 21790 10492
rect 22094 10480 22100 10492
rect 22152 10520 22158 10532
rect 22649 10523 22707 10529
rect 22649 10520 22661 10523
rect 22152 10492 22661 10520
rect 22152 10480 22158 10492
rect 22649 10489 22661 10492
rect 22695 10489 22707 10523
rect 22649 10483 22707 10489
rect 26835 10523 26893 10529
rect 26835 10489 26847 10523
rect 26881 10520 26893 10523
rect 27982 10520 27988 10532
rect 26881 10492 27988 10520
rect 26881 10489 26893 10492
rect 26835 10483 26893 10489
rect 27982 10480 27988 10492
rect 28040 10480 28046 10532
rect 33336 10520 33364 10551
rect 33410 10548 33416 10600
rect 33468 10588 33474 10600
rect 35250 10588 35256 10600
rect 33468 10560 35256 10588
rect 33468 10548 33474 10560
rect 35250 10548 35256 10560
rect 35308 10548 35314 10600
rect 35434 10588 35440 10600
rect 35395 10560 35440 10588
rect 35434 10548 35440 10560
rect 35492 10588 35498 10600
rect 35989 10591 36047 10597
rect 35989 10588 36001 10591
rect 35492 10560 36001 10588
rect 35492 10548 35498 10560
rect 35989 10557 36001 10560
rect 36035 10557 36047 10591
rect 35989 10551 36047 10557
rect 33336 10492 33824 10520
rect 33796 10464 33824 10492
rect 21818 10452 21824 10464
rect 21284 10424 21824 10452
rect 20947 10415 21005 10421
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 22002 10461 22008 10464
rect 21959 10455 22008 10461
rect 21959 10421 21971 10455
rect 22005 10421 22008 10455
rect 21959 10415 22008 10421
rect 22002 10412 22008 10415
rect 22060 10412 22066 10464
rect 22370 10452 22376 10464
rect 22331 10424 22376 10452
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 27246 10412 27252 10464
rect 27304 10452 27310 10464
rect 27847 10455 27905 10461
rect 27847 10452 27859 10455
rect 27304 10424 27859 10452
rect 27304 10412 27310 10424
rect 27847 10421 27859 10424
rect 27893 10421 27905 10455
rect 27847 10415 27905 10421
rect 33367 10455 33425 10461
rect 33367 10421 33379 10455
rect 33413 10452 33425 10455
rect 33594 10452 33600 10464
rect 33413 10424 33600 10452
rect 33413 10421 33425 10424
rect 33367 10415 33425 10421
rect 33594 10412 33600 10424
rect 33652 10412 33658 10464
rect 33778 10452 33784 10464
rect 33739 10424 33784 10452
rect 33778 10412 33784 10424
rect 33836 10412 33842 10464
rect 34146 10412 34152 10464
rect 34204 10452 34210 10464
rect 34425 10455 34483 10461
rect 34425 10452 34437 10455
rect 34204 10424 34437 10452
rect 34204 10412 34210 10424
rect 34425 10421 34437 10424
rect 34471 10452 34483 10455
rect 34790 10452 34796 10464
rect 34471 10424 34796 10452
rect 34471 10421 34483 10424
rect 34425 10415 34483 10421
rect 34790 10412 34796 10424
rect 34848 10412 34854 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 3510 10248 3516 10260
rect 3471 10220 3516 10248
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6880 10220 6929 10248
rect 6880 10208 6886 10220
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 10778 10248 10784 10260
rect 10739 10220 10784 10248
rect 6917 10211 6975 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 13446 10248 13452 10260
rect 13407 10220 13452 10248
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 14056 10220 14105 10248
rect 14056 10208 14062 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 27157 10251 27215 10257
rect 27157 10217 27169 10251
rect 27203 10248 27215 10251
rect 27246 10248 27252 10260
rect 27203 10220 27252 10248
rect 27203 10217 27215 10220
rect 27157 10211 27215 10217
rect 27246 10208 27252 10220
rect 27304 10208 27310 10260
rect 35621 10251 35679 10257
rect 35621 10217 35633 10251
rect 35667 10248 35679 10251
rect 35710 10248 35716 10260
rect 35667 10220 35716 10248
rect 35667 10217 35679 10220
rect 35621 10211 35679 10217
rect 35710 10208 35716 10220
rect 35768 10208 35774 10260
rect 2424 10180 2452 10208
rect 2774 10180 2780 10192
rect 2424 10152 2780 10180
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 27430 10180 27436 10192
rect 27391 10152 27436 10180
rect 27430 10140 27436 10152
rect 27488 10140 27494 10192
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1854 10112 1860 10124
rect 1767 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10112 1918 10124
rect 2314 10112 2320 10124
rect 1912 10084 2320 10112
rect 1912 10072 1918 10084
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 3050 10121 3056 10124
rect 3028 10115 3056 10121
rect 3028 10081 3040 10115
rect 3028 10075 3056 10081
rect 3050 10072 3056 10075
rect 3108 10072 3114 10124
rect 4246 10112 4252 10124
rect 4207 10084 4252 10112
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5718 10121 5724 10124
rect 5696 10115 5724 10121
rect 5696 10081 5708 10115
rect 5696 10075 5724 10081
rect 5718 10072 5724 10075
rect 5776 10072 5782 10124
rect 6638 10112 6644 10124
rect 6599 10084 6644 10112
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6972 10084 7113 10112
rect 6972 10072 6978 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 8640 10115 8698 10121
rect 8640 10081 8652 10115
rect 8686 10112 8698 10115
rect 9030 10112 9036 10124
rect 8686 10084 9036 10112
rect 8686 10081 8698 10084
rect 8640 10075 8698 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 9824 10084 10517 10112
rect 9824 10072 9830 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11514 10112 11520 10124
rect 11103 10084 11520 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 13722 10112 13728 10124
rect 12851 10084 13728 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15841 10115 15899 10121
rect 15841 10112 15853 10115
rect 15436 10084 15853 10112
rect 15436 10072 15442 10084
rect 15841 10081 15853 10084
rect 15887 10081 15899 10115
rect 16298 10112 16304 10124
rect 16259 10084 16304 10112
rect 15841 10075 15899 10081
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 17954 10112 17960 10124
rect 17915 10084 17960 10112
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18230 10112 18236 10124
rect 18191 10084 18236 10112
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 19334 10072 19340 10124
rect 19392 10121 19398 10124
rect 19392 10115 19430 10121
rect 19418 10081 19430 10115
rect 20936 10115 20994 10121
rect 20936 10112 20948 10115
rect 19392 10075 19430 10081
rect 20824 10084 20948 10112
rect 19392 10072 19398 10075
rect 20824 10056 20852 10084
rect 20936 10081 20948 10084
rect 20982 10081 20994 10115
rect 21948 10115 22006 10121
rect 21948 10112 21960 10115
rect 20936 10075 20994 10081
rect 21284 10084 21960 10112
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 4614 10044 4620 10056
rect 4575 10016 4620 10044
rect 1949 10007 2007 10013
rect 1854 9936 1860 9988
rect 1912 9976 1918 9988
rect 1964 9976 1992 10007
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12618 10044 12624 10056
rect 12492 10016 12624 10044
rect 12492 10004 12498 10016
rect 12618 10004 12624 10016
rect 12676 10044 12682 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12676 10016 13185 10044
rect 12676 10004 12682 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 16390 10044 16396 10056
rect 16351 10016 16396 10044
rect 13173 10007 13231 10013
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 18322 10044 18328 10056
rect 18283 10016 18328 10044
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 20806 10004 20812 10056
rect 20864 10004 20870 10056
rect 1912 9948 1992 9976
rect 1912 9936 1918 9948
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12943 9979 13001 9985
rect 12943 9976 12955 9979
rect 12860 9948 12955 9976
rect 12860 9936 12866 9948
rect 12943 9945 12955 9948
rect 12989 9945 13001 9979
rect 12943 9939 13001 9945
rect 20622 9936 20628 9988
rect 20680 9976 20686 9988
rect 21284 9976 21312 10084
rect 21948 10081 21960 10084
rect 21994 10112 22006 10115
rect 22922 10112 22928 10124
rect 21994 10081 22023 10112
rect 22883 10084 22928 10112
rect 21948 10075 22023 10081
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10044 21511 10047
rect 21542 10044 21548 10056
rect 21499 10016 21548 10044
rect 21499 10013 21511 10016
rect 21453 10007 21511 10013
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 21995 10044 22023 10075
rect 22922 10072 22928 10084
rect 22980 10072 22986 10124
rect 24118 10072 24124 10124
rect 24176 10112 24182 10124
rect 25498 10121 25504 10124
rect 24397 10115 24455 10121
rect 24397 10112 24409 10115
rect 24176 10084 24409 10112
rect 24176 10072 24182 10084
rect 24397 10081 24409 10084
rect 24443 10081 24455 10115
rect 24397 10075 24455 10081
rect 25476 10115 25504 10121
rect 25476 10081 25488 10115
rect 25476 10075 25504 10081
rect 25498 10072 25504 10075
rect 25556 10072 25562 10124
rect 28902 10121 28908 10124
rect 28880 10115 28908 10121
rect 28880 10081 28892 10115
rect 28880 10075 28908 10081
rect 28902 10072 28908 10075
rect 28960 10072 28966 10124
rect 33410 10072 33416 10124
rect 33468 10121 33474 10124
rect 33468 10115 33506 10121
rect 33494 10081 33506 10115
rect 33468 10075 33506 10081
rect 34492 10115 34550 10121
rect 34492 10081 34504 10115
rect 34538 10112 34550 10115
rect 34698 10112 34704 10124
rect 34538 10084 34704 10112
rect 34538 10081 34550 10084
rect 34492 10075 34550 10081
rect 33468 10072 33474 10075
rect 34698 10072 34704 10084
rect 34756 10072 34762 10124
rect 35437 10115 35495 10121
rect 35437 10081 35449 10115
rect 35483 10112 35495 10115
rect 35802 10112 35808 10124
rect 35483 10084 35808 10112
rect 35483 10081 35495 10084
rect 35437 10075 35495 10081
rect 35802 10072 35808 10084
rect 35860 10072 35866 10124
rect 36262 10072 36268 10124
rect 36320 10112 36326 10124
rect 36608 10115 36666 10121
rect 36608 10112 36620 10115
rect 36320 10084 36620 10112
rect 36320 10072 36326 10084
rect 36608 10081 36620 10084
rect 36654 10112 36666 10115
rect 37182 10112 37188 10124
rect 36654 10084 37188 10112
rect 36654 10081 36666 10084
rect 36608 10075 36666 10081
rect 37182 10072 37188 10084
rect 37240 10072 37246 10124
rect 22462 10044 22468 10056
rect 21995 10016 22468 10044
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 27341 10047 27399 10053
rect 27341 10013 27353 10047
rect 27387 10044 27399 10047
rect 27522 10044 27528 10056
rect 27387 10016 27528 10044
rect 27387 10013 27399 10016
rect 27341 10007 27399 10013
rect 27522 10004 27528 10016
rect 27580 10004 27586 10056
rect 27985 10047 28043 10053
rect 27985 10013 27997 10047
rect 28031 10044 28043 10047
rect 29178 10044 29184 10056
rect 28031 10016 29184 10044
rect 28031 10013 28043 10016
rect 27985 10007 28043 10013
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 20680 9948 21312 9976
rect 20680 9936 20686 9948
rect 21634 9936 21640 9988
rect 21692 9976 21698 9988
rect 22051 9979 22109 9985
rect 22051 9976 22063 9979
rect 21692 9948 22063 9976
rect 21692 9936 21698 9948
rect 22051 9945 22063 9948
rect 22097 9945 22109 9979
rect 22051 9939 22109 9945
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 2777 9911 2835 9917
rect 2777 9908 2789 9911
rect 2556 9880 2789 9908
rect 2556 9868 2562 9880
rect 2777 9877 2789 9880
rect 2823 9877 2835 9911
rect 2777 9871 2835 9877
rect 3099 9911 3157 9917
rect 3099 9877 3111 9911
rect 3145 9908 3157 9911
rect 3234 9908 3240 9920
rect 3145 9880 3240 9908
rect 3145 9877 3157 9880
rect 3099 9871 3157 9877
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5767 9911 5825 9917
rect 5767 9908 5779 9911
rect 5592 9880 5779 9908
rect 5592 9868 5598 9880
rect 5767 9877 5779 9880
rect 5813 9877 5825 9911
rect 5767 9871 5825 9877
rect 8711 9911 8769 9917
rect 8711 9877 8723 9911
rect 8757 9908 8769 9911
rect 9582 9908 9588 9920
rect 8757 9880 9588 9908
rect 8757 9877 8769 9880
rect 8711 9871 8769 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 11698 9908 11704 9920
rect 11659 9880 11704 9908
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13170 9908 13176 9920
rect 13127 9880 13176 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 14148 9880 14473 9908
rect 14148 9868 14154 9880
rect 14461 9877 14473 9880
rect 14507 9877 14519 9911
rect 14461 9871 14519 9877
rect 19475 9911 19533 9917
rect 19475 9877 19487 9911
rect 19521 9908 19533 9911
rect 19702 9908 19708 9920
rect 19521 9880 19708 9908
rect 19521 9877 19533 9880
rect 19475 9871 19533 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 19886 9908 19892 9920
rect 19847 9880 19892 9908
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 21039 9911 21097 9917
rect 21039 9877 21051 9911
rect 21085 9908 21097 9911
rect 21266 9908 21272 9920
rect 21085 9880 21272 9908
rect 21085 9877 21097 9880
rect 21039 9871 21097 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 21729 9911 21787 9917
rect 21729 9908 21741 9911
rect 21508 9880 21741 9908
rect 21508 9868 21514 9880
rect 21729 9877 21741 9880
rect 21775 9877 21787 9911
rect 21729 9871 21787 9877
rect 23109 9911 23167 9917
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23750 9908 23756 9920
rect 23155 9880 23756 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23750 9868 23756 9880
rect 23808 9908 23814 9920
rect 24121 9911 24179 9917
rect 24121 9908 24133 9911
rect 23808 9880 24133 9908
rect 23808 9868 23814 9880
rect 24121 9877 24133 9880
rect 24167 9908 24179 9911
rect 24486 9908 24492 9920
rect 24167 9880 24492 9908
rect 24167 9877 24179 9880
rect 24121 9871 24179 9877
rect 24486 9868 24492 9880
rect 24544 9868 24550 9920
rect 24578 9868 24584 9920
rect 24636 9908 24642 9920
rect 25547 9911 25605 9917
rect 24636 9880 24681 9908
rect 24636 9868 24642 9880
rect 25547 9877 25559 9911
rect 25593 9908 25605 9911
rect 25958 9908 25964 9920
rect 25593 9880 25964 9908
rect 25593 9877 25605 9880
rect 25547 9871 25605 9877
rect 25958 9868 25964 9880
rect 26016 9868 26022 9920
rect 28442 9868 28448 9920
rect 28500 9908 28506 9920
rect 28951 9911 29009 9917
rect 28951 9908 28963 9911
rect 28500 9880 28963 9908
rect 28500 9868 28506 9880
rect 28951 9877 28963 9880
rect 28997 9877 29009 9911
rect 28951 9871 29009 9877
rect 33551 9911 33609 9917
rect 33551 9877 33563 9911
rect 33597 9908 33609 9911
rect 34146 9908 34152 9920
rect 33597 9880 34152 9908
rect 33597 9877 33609 9880
rect 33551 9871 33609 9877
rect 34146 9868 34152 9880
rect 34204 9868 34210 9920
rect 34563 9911 34621 9917
rect 34563 9877 34575 9911
rect 34609 9908 34621 9911
rect 35250 9908 35256 9920
rect 34609 9880 35256 9908
rect 34609 9877 34621 9880
rect 34563 9871 34621 9877
rect 35250 9868 35256 9880
rect 35308 9868 35314 9920
rect 35342 9868 35348 9920
rect 35400 9908 35406 9920
rect 36679 9911 36737 9917
rect 36679 9908 36691 9911
rect 35400 9880 36691 9908
rect 35400 9868 35406 9880
rect 36679 9877 36691 9880
rect 36725 9877 36737 9911
rect 36679 9871 36737 9877
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 2869 9707 2927 9713
rect 2869 9673 2881 9707
rect 2915 9704 2927 9707
rect 3050 9704 3056 9716
rect 2915 9676 3056 9704
rect 2915 9673 2927 9676
rect 2869 9667 2927 9673
rect 3050 9664 3056 9676
rect 3108 9704 3114 9716
rect 3326 9704 3332 9716
rect 3108 9676 3332 9704
rect 3108 9664 3114 9676
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 4522 9704 4528 9716
rect 4172 9676 4528 9704
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 2832 9608 3985 9636
rect 2832 9596 2838 9608
rect 3973 9605 3985 9608
rect 4019 9636 4031 9639
rect 4172 9636 4200 9676
rect 4522 9664 4528 9676
rect 4580 9704 4586 9716
rect 6273 9707 6331 9713
rect 4580 9676 5488 9704
rect 4580 9664 4586 9676
rect 4019 9608 4200 9636
rect 5460 9636 5488 9676
rect 6273 9673 6285 9707
rect 6319 9704 6331 9707
rect 6638 9704 6644 9716
rect 6319 9676 6644 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 8202 9704 8208 9716
rect 6932 9676 8208 9704
rect 6932 9648 6960 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 9824 9676 10241 9704
rect 9824 9664 9830 9676
rect 10229 9673 10241 9676
rect 10275 9673 10287 9707
rect 11514 9704 11520 9716
rect 11475 9676 11520 9704
rect 10229 9667 10287 9673
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 13078 9704 13084 9716
rect 12860 9676 13084 9704
rect 12860 9664 12866 9676
rect 13078 9664 13084 9676
rect 13136 9704 13142 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13136 9676 13461 9704
rect 13136 9664 13142 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 13449 9667 13507 9673
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 17954 9704 17960 9716
rect 17880 9676 17960 9704
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 5460 9608 6561 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 6549 9605 6561 9608
rect 6595 9636 6607 9639
rect 6914 9636 6920 9648
rect 6595 9608 6920 9636
rect 6595 9605 6607 9608
rect 6549 9599 6607 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 8220 9636 8248 9664
rect 11790 9636 11796 9648
rect 8220 9608 8524 9636
rect 11751 9608 11796 9636
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3510 9568 3516 9580
rect 3099 9540 3516 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 5868 9540 7205 9568
rect 5868 9528 5874 9540
rect 7193 9537 7205 9540
rect 7239 9568 7251 9571
rect 7558 9568 7564 9580
rect 7239 9540 7564 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 1670 9500 1676 9512
rect 1583 9472 1676 9500
rect 1670 9460 1676 9472
rect 1728 9500 1734 9512
rect 1949 9503 2007 9509
rect 1728 9472 1808 9500
rect 1728 9460 1734 9472
rect 1780 9364 1808 9472
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2406 9500 2412 9512
rect 1995 9472 2412 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4479 9472 4629 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4617 9469 4629 9472
rect 4663 9500 4675 9503
rect 5166 9500 5172 9512
rect 4663 9472 5172 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 8386 9500 8392 9512
rect 8347 9472 8392 9500
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8496 9500 8524 9608
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12452 9608 13216 9636
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 12452 9568 12480 9608
rect 13188 9580 13216 9608
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13780 9608 13829 9636
rect 13780 9596 13786 9608
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 15286 9596 15292 9648
rect 15344 9636 15350 9648
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 15344 9608 15853 9636
rect 15344 9596 15350 9608
rect 15841 9605 15853 9608
rect 15887 9636 15899 9639
rect 16298 9636 16304 9648
rect 15887 9608 16304 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 17880 9636 17908 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 19334 9704 19340 9716
rect 19295 9676 19340 9704
rect 19334 9664 19340 9676
rect 19392 9704 19398 9716
rect 20806 9704 20812 9716
rect 19392 9676 20812 9704
rect 19392 9664 19398 9676
rect 20806 9664 20812 9676
rect 20864 9704 20870 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20864 9676 20913 9704
rect 20864 9664 20870 9676
rect 20901 9673 20913 9676
rect 20947 9673 20959 9707
rect 25498 9704 25504 9716
rect 25459 9676 25504 9704
rect 20901 9667 20959 9673
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 33410 9704 33416 9716
rect 33371 9676 33416 9704
rect 33410 9664 33416 9676
rect 33468 9664 33474 9716
rect 17420 9608 17908 9636
rect 12299 9540 12480 9568
rect 12529 9571 12587 9577
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12802 9568 12808 9580
rect 12575 9540 12808 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 13906 9568 13912 9580
rect 13228 9540 13912 9568
rect 13228 9528 13234 9540
rect 13906 9528 13912 9540
rect 13964 9568 13970 9580
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 13964 9540 14381 9568
rect 13964 9528 13970 9540
rect 14369 9537 14381 9540
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15712 9540 16037 9568
rect 15712 9528 15718 9540
rect 16025 9537 16037 9540
rect 16071 9568 16083 9571
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 16071 9540 16957 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 8662 9500 8668 9512
rect 8496 9472 8668 9500
rect 8662 9460 8668 9472
rect 8720 9500 8726 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8720 9472 8861 9500
rect 8720 9460 8726 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 10502 9500 10508 9512
rect 10463 9472 10508 9500
rect 8849 9463 8907 9469
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10928 9472 10977 9500
rect 10928 9460 10934 9472
rect 10965 9469 10977 9472
rect 11011 9500 11023 9503
rect 11514 9500 11520 9512
rect 11011 9472 11520 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14323 9472 14473 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 14461 9469 14473 9472
rect 14507 9500 14519 9503
rect 14642 9500 14648 9512
rect 14507 9472 14648 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 2038 9392 2044 9444
rect 2096 9432 2102 9444
rect 2133 9435 2191 9441
rect 2133 9432 2145 9435
rect 2096 9404 2145 9432
rect 2096 9392 2102 9404
rect 2133 9401 2145 9404
rect 2179 9401 2191 9435
rect 2133 9395 2191 9401
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3510 9432 3516 9444
rect 3191 9404 3516 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3694 9432 3700 9444
rect 3655 9404 3700 9432
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 6270 9432 6276 9444
rect 5307 9404 6276 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 6917 9435 6975 9441
rect 6917 9401 6929 9435
rect 6963 9401 6975 9435
rect 6917 9395 6975 9401
rect 2498 9364 2504 9376
rect 1780 9336 2504 9364
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 5718 9364 5724 9376
rect 5679 9336 5724 9364
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 6932 9364 6960 9395
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 9953 9435 10011 9441
rect 7064 9404 7109 9432
rect 7064 9392 7070 9404
rect 9953 9401 9965 9435
rect 9999 9432 10011 9435
rect 10888 9432 10916 9460
rect 9999 9404 10916 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 12621 9435 12679 9441
rect 12621 9432 12633 9435
rect 12584 9404 12633 9432
rect 12584 9392 12590 9404
rect 12621 9401 12633 9404
rect 12667 9401 12679 9435
rect 12621 9395 12679 9401
rect 13173 9435 13231 9441
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 13538 9432 13544 9444
rect 13219 9404 13544 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 16666 9432 16672 9444
rect 16172 9404 16217 9432
rect 16627 9404 16672 9432
rect 16172 9392 16178 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 7098 9364 7104 9376
rect 6932 9336 7104 9364
rect 7098 9324 7104 9336
rect 7156 9364 7162 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7156 9336 7849 9364
rect 7156 9324 7162 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 8352 9336 8493 9364
rect 8352 9324 8358 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 8481 9327 8539 9333
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9088 9336 9413 9364
rect 9088 9324 9094 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 10502 9364 10508 9376
rect 10463 9336 10508 9364
rect 9401 9327 9459 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 12802 9364 12808 9376
rect 11848 9336 12808 9364
rect 11848 9324 11854 9336
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 13814 9364 13820 9376
rect 13320 9336 13820 9364
rect 13320 9324 13326 9336
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17420 9373 17448 9608
rect 26602 9596 26608 9648
rect 26660 9636 26666 9648
rect 28626 9636 28632 9648
rect 26660 9608 28632 9636
rect 26660 9596 26666 9608
rect 28626 9596 28632 9608
rect 28684 9596 28690 9648
rect 32306 9636 32312 9648
rect 32267 9608 32312 9636
rect 32306 9596 32312 9608
rect 32364 9596 32370 9648
rect 35526 9636 35532 9648
rect 35487 9608 35532 9636
rect 35526 9596 35532 9608
rect 35584 9596 35590 9648
rect 36630 9636 36636 9648
rect 36591 9608 36636 9636
rect 36630 9596 36636 9608
rect 36688 9596 36694 9648
rect 20530 9528 20536 9580
rect 20588 9568 20594 9580
rect 21729 9571 21787 9577
rect 21729 9568 21741 9571
rect 20588 9540 21741 9568
rect 20588 9528 20594 9540
rect 21729 9537 21741 9540
rect 21775 9568 21787 9571
rect 21910 9568 21916 9580
rect 21775 9540 21916 9568
rect 21775 9537 21787 9540
rect 21729 9531 21787 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 24762 9568 24768 9580
rect 24723 9540 24768 9568
rect 24762 9528 24768 9540
rect 24820 9528 24826 9580
rect 27246 9528 27252 9580
rect 27304 9568 27310 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 27304 9540 27445 9568
rect 27304 9528 27310 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 18012 9472 18061 9500
rect 18012 9460 18018 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18506 9500 18512 9512
rect 18467 9472 18512 9500
rect 18049 9463 18107 9469
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 19518 9460 19524 9512
rect 19576 9500 19582 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19576 9472 19625 9500
rect 19576 9460 19582 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19886 9460 19892 9512
rect 19944 9500 19950 9512
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19944 9472 20085 9500
rect 19944 9460 19950 9472
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 22462 9500 22468 9512
rect 22423 9472 22468 9500
rect 20073 9463 20131 9469
rect 22462 9460 22468 9472
rect 22520 9460 22526 9512
rect 24397 9503 24455 9509
rect 24397 9469 24409 9503
rect 24443 9469 24455 9503
rect 24397 9463 24455 9469
rect 18230 9432 18236 9444
rect 17880 9404 18236 9432
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17092 9336 17417 9364
rect 17092 9324 17098 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17405 9327 17463 9333
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17736 9336 17785 9364
rect 17736 9324 17742 9336
rect 17773 9333 17785 9336
rect 17819 9364 17831 9367
rect 17880 9364 17908 9404
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 21450 9432 21456 9444
rect 21411 9404 21456 9432
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 21542 9392 21548 9444
rect 21600 9432 21606 9444
rect 21600 9404 21645 9432
rect 21600 9392 21606 9404
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 22922 9432 22928 9444
rect 22152 9404 22928 9432
rect 22152 9392 22158 9404
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 24026 9432 24032 9444
rect 23939 9404 24032 9432
rect 24026 9392 24032 9404
rect 24084 9432 24090 9444
rect 24412 9432 24440 9463
rect 24486 9460 24492 9512
rect 24544 9500 24550 9512
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 24544 9472 24593 9500
rect 24544 9460 24550 9472
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 26234 9460 26240 9512
rect 26292 9500 26298 9512
rect 26396 9503 26454 9509
rect 26396 9500 26408 9503
rect 26292 9472 26408 9500
rect 26292 9460 26298 9472
rect 26396 9469 26408 9472
rect 26442 9500 26454 9503
rect 29340 9503 29398 9509
rect 26442 9472 26924 9500
rect 26442 9469 26454 9472
rect 26396 9463 26454 9469
rect 24854 9432 24860 9444
rect 24084 9404 24860 9432
rect 24084 9392 24090 9404
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 26896 9376 26924 9472
rect 29340 9469 29352 9503
rect 29386 9500 29398 9503
rect 29386 9472 29868 9500
rect 29386 9469 29398 9472
rect 29340 9463 29398 9469
rect 27249 9435 27307 9441
rect 27249 9401 27261 9435
rect 27295 9432 27307 9435
rect 27430 9432 27436 9444
rect 27295 9404 27436 9432
rect 27295 9401 27307 9404
rect 27249 9395 27307 9401
rect 27430 9392 27436 9404
rect 27488 9432 27494 9444
rect 27525 9435 27583 9441
rect 27525 9432 27537 9435
rect 27488 9404 27537 9432
rect 27488 9392 27494 9404
rect 27525 9401 27537 9404
rect 27571 9401 27583 9435
rect 28074 9432 28080 9444
rect 28035 9404 28080 9432
rect 27525 9395 27583 9401
rect 18138 9364 18144 9376
rect 17819 9336 17908 9364
rect 18099 9336 18144 9364
rect 17819 9333 17831 9336
rect 17773 9327 17831 9333
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 19886 9364 19892 9376
rect 19847 9336 19892 9364
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 26467 9367 26525 9373
rect 26467 9333 26479 9367
rect 26513 9364 26525 9367
rect 26694 9364 26700 9376
rect 26513 9336 26700 9364
rect 26513 9333 26525 9336
rect 26467 9327 26525 9333
rect 26694 9324 26700 9336
rect 26752 9324 26758 9376
rect 26878 9364 26884 9376
rect 26839 9336 26884 9364
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 27540 9364 27568 9395
rect 28074 9392 28080 9404
rect 28132 9392 28138 9444
rect 29840 9376 29868 9472
rect 30190 9460 30196 9512
rect 30248 9500 30254 9512
rect 30285 9503 30343 9509
rect 30285 9500 30297 9503
rect 30248 9472 30297 9500
rect 30248 9460 30254 9472
rect 30285 9469 30297 9472
rect 30331 9500 30343 9503
rect 30745 9503 30803 9509
rect 30745 9500 30757 9503
rect 30331 9472 30757 9500
rect 30331 9469 30343 9472
rect 30285 9463 30343 9469
rect 30745 9469 30757 9472
rect 30791 9469 30803 9503
rect 30745 9463 30803 9469
rect 31824 9503 31882 9509
rect 31824 9469 31836 9503
rect 31870 9500 31882 9503
rect 32324 9500 32352 9596
rect 32582 9568 32588 9580
rect 32543 9540 32588 9568
rect 32582 9528 32588 9540
rect 32640 9528 32646 9580
rect 35158 9568 35164 9580
rect 35119 9540 35164 9568
rect 35158 9528 35164 9540
rect 35216 9528 35222 9580
rect 31870 9472 32352 9500
rect 32600 9500 32628 9528
rect 32804 9503 32862 9509
rect 32804 9500 32816 9503
rect 32600 9472 32816 9500
rect 31870 9469 31882 9472
rect 31824 9463 31882 9469
rect 32804 9469 32816 9472
rect 32850 9469 32862 9503
rect 32804 9463 32862 9469
rect 33686 9460 33692 9512
rect 33744 9500 33750 9512
rect 33848 9503 33906 9509
rect 33848 9500 33860 9503
rect 33744 9472 33860 9500
rect 33744 9460 33750 9472
rect 33848 9469 33860 9472
rect 33894 9500 33906 9503
rect 35176 9500 35204 9528
rect 35345 9503 35403 9509
rect 35345 9500 35357 9503
rect 33894 9472 34376 9500
rect 35176 9472 35357 9500
rect 33894 9469 33906 9472
rect 33848 9463 33906 9469
rect 34348 9441 34376 9472
rect 35345 9469 35357 9472
rect 35391 9469 35403 9503
rect 36446 9500 36452 9512
rect 36407 9472 36452 9500
rect 35345 9463 35403 9469
rect 36446 9460 36452 9472
rect 36504 9500 36510 9512
rect 37001 9503 37059 9509
rect 37001 9500 37013 9503
rect 36504 9472 37013 9500
rect 36504 9460 36510 9472
rect 37001 9469 37013 9472
rect 37047 9469 37059 9503
rect 37001 9463 37059 9469
rect 34333 9435 34391 9441
rect 34333 9401 34345 9435
rect 34379 9432 34391 9435
rect 36078 9432 36084 9444
rect 34379 9404 36084 9432
rect 34379 9401 34391 9404
rect 34333 9395 34391 9401
rect 36078 9392 36084 9404
rect 36136 9392 36142 9444
rect 28353 9367 28411 9373
rect 28353 9364 28365 9367
rect 27540 9336 28365 9364
rect 28353 9333 28365 9336
rect 28399 9333 28411 9367
rect 28353 9327 28411 9333
rect 28718 9324 28724 9376
rect 28776 9364 28782 9376
rect 28813 9367 28871 9373
rect 28813 9364 28825 9367
rect 28776 9336 28825 9364
rect 28776 9324 28782 9336
rect 28813 9333 28825 9336
rect 28859 9364 28871 9367
rect 28902 9364 28908 9376
rect 28859 9336 28908 9364
rect 28859 9333 28871 9336
rect 28813 9327 28871 9333
rect 28902 9324 28908 9336
rect 28960 9324 28966 9376
rect 29086 9324 29092 9376
rect 29144 9364 29150 9376
rect 29411 9367 29469 9373
rect 29411 9364 29423 9367
rect 29144 9336 29423 9364
rect 29144 9324 29150 9336
rect 29411 9333 29423 9336
rect 29457 9333 29469 9367
rect 29822 9364 29828 9376
rect 29783 9336 29828 9364
rect 29411 9327 29469 9333
rect 29822 9324 29828 9336
rect 29880 9324 29886 9376
rect 30466 9364 30472 9376
rect 30427 9336 30472 9364
rect 30466 9324 30472 9336
rect 30524 9324 30530 9376
rect 31895 9367 31953 9373
rect 31895 9333 31907 9367
rect 31941 9364 31953 9367
rect 32674 9364 32680 9376
rect 31941 9336 32680 9364
rect 31941 9333 31953 9336
rect 31895 9327 31953 9333
rect 32674 9324 32680 9336
rect 32732 9324 32738 9376
rect 32907 9367 32965 9373
rect 32907 9333 32919 9367
rect 32953 9364 32965 9367
rect 33318 9364 33324 9376
rect 32953 9336 33324 9364
rect 32953 9333 32965 9336
rect 32907 9327 32965 9333
rect 33318 9324 33324 9336
rect 33376 9324 33382 9376
rect 33502 9324 33508 9376
rect 33560 9364 33566 9376
rect 33919 9367 33977 9373
rect 33919 9364 33931 9367
rect 33560 9336 33931 9364
rect 33560 9324 33566 9336
rect 33919 9333 33931 9336
rect 33965 9333 33977 9367
rect 34698 9364 34704 9376
rect 34611 9336 34704 9364
rect 33919 9327 33977 9333
rect 34698 9324 34704 9336
rect 34756 9364 34762 9376
rect 35158 9364 35164 9376
rect 34756 9336 35164 9364
rect 34756 9324 34762 9336
rect 35158 9324 35164 9336
rect 35216 9324 35222 9376
rect 35894 9364 35900 9376
rect 35855 9336 35900 9364
rect 35894 9324 35900 9336
rect 35952 9324 35958 9376
rect 37274 9324 37280 9376
rect 37332 9364 37338 9376
rect 37369 9367 37427 9373
rect 37369 9364 37381 9367
rect 37332 9336 37381 9364
rect 37332 9324 37338 9336
rect 37369 9333 37381 9336
rect 37415 9333 37427 9367
rect 37369 9327 37427 9333
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2498 9160 2504 9172
rect 1995 9132 2504 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 10652 9132 11069 9160
rect 10652 9120 10658 9132
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11422 9160 11428 9172
rect 11383 9132 11428 9160
rect 11057 9123 11115 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 12676 9132 12817 9160
rect 12676 9120 12682 9132
rect 12805 9129 12817 9132
rect 12851 9160 12863 9163
rect 13170 9160 13176 9172
rect 12851 9132 13176 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 16172 9132 16221 9160
rect 16172 9120 16178 9132
rect 16209 9129 16221 9132
rect 16255 9160 16267 9163
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16255 9132 16497 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 16485 9123 16543 9129
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 18012 9132 18061 9160
rect 18012 9120 18018 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18690 9160 18696 9172
rect 18651 9132 18696 9160
rect 18049 9123 18107 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 20070 9160 20076 9172
rect 19983 9132 20076 9160
rect 20070 9120 20076 9132
rect 20128 9160 20134 9172
rect 20622 9160 20628 9172
rect 20128 9132 20628 9160
rect 20128 9120 20134 9132
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 21818 9120 21824 9172
rect 21876 9160 21882 9172
rect 22186 9160 22192 9172
rect 21876 9132 22192 9160
rect 21876 9120 21882 9132
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 23891 9163 23949 9169
rect 23891 9160 23903 9163
rect 23532 9132 23903 9160
rect 23532 9120 23538 9132
rect 23891 9129 23903 9132
rect 23937 9129 23949 9163
rect 23891 9123 23949 9129
rect 26694 9120 26700 9172
rect 26752 9160 26758 9172
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 26752 9132 28273 9160
rect 26752 9120 26758 9132
rect 27724 9104 27752 9132
rect 28261 9129 28273 9132
rect 28307 9129 28319 9163
rect 28261 9123 28319 9129
rect 28445 9163 28503 9169
rect 28445 9129 28457 9163
rect 28491 9160 28503 9163
rect 28902 9160 28908 9172
rect 28491 9132 28908 9160
rect 28491 9129 28503 9132
rect 28445 9123 28503 9129
rect 28902 9120 28908 9132
rect 28960 9120 28966 9172
rect 33594 9160 33600 9172
rect 33555 9132 33600 9160
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 2593 9095 2651 9101
rect 2593 9061 2605 9095
rect 2639 9092 2651 9095
rect 2866 9092 2872 9104
rect 2639 9064 2872 9092
rect 2639 9061 2651 9064
rect 2593 9055 2651 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3694 9092 3700 9104
rect 3191 9064 3700 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3694 9052 3700 9064
rect 3752 9052 3758 9104
rect 4246 9092 4252 9104
rect 4207 9064 4252 9092
rect 4246 9052 4252 9064
rect 4304 9052 4310 9104
rect 7374 9092 7380 9104
rect 7335 9064 7380 9092
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 11793 9095 11851 9101
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 11882 9092 11888 9104
rect 11839 9064 11888 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 11882 9052 11888 9064
rect 11940 9092 11946 9104
rect 13357 9095 13415 9101
rect 13357 9092 13369 9095
rect 11940 9064 13369 9092
rect 11940 9052 11946 9064
rect 13357 9061 13369 9064
rect 13403 9092 13415 9095
rect 13446 9092 13452 9104
rect 13403 9064 13452 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15610 9095 15668 9101
rect 15610 9092 15622 9095
rect 15436 9064 15622 9092
rect 15436 9052 15442 9064
rect 15610 9061 15622 9064
rect 15656 9061 15668 9095
rect 17218 9092 17224 9104
rect 17179 9064 17224 9092
rect 15610 9055 15668 9061
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 18506 9092 18512 9104
rect 18419 9064 18512 9092
rect 18506 9052 18512 9064
rect 18564 9092 18570 9104
rect 21266 9092 21272 9104
rect 18564 9064 19196 9092
rect 21227 9064 21272 9092
rect 18564 9052 18570 9064
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 9024 1522 9027
rect 1670 9024 1676 9036
rect 1510 8996 1676 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 5626 9024 5632 9036
rect 5587 8996 5632 9024
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 6270 9024 6276 9036
rect 5951 8996 6276 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 10192 8996 10517 9024
rect 10192 8984 10198 8996
rect 10505 8993 10517 8996
rect 10551 9024 10563 9027
rect 10870 9024 10876 9036
rect 10551 8996 10876 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15252 8996 15301 9024
rect 15252 8984 15258 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 18230 8984 18236 9036
rect 18288 9024 18294 9036
rect 19168 9033 19196 9064
rect 21266 9052 21272 9064
rect 21324 9052 21330 9104
rect 21358 9052 21364 9104
rect 21416 9092 21422 9104
rect 21416 9064 21461 9092
rect 21416 9052 21422 9064
rect 24578 9052 24584 9104
rect 24636 9092 24642 9104
rect 24636 9064 24992 9092
rect 24636 9052 24642 9064
rect 24964 9036 24992 9064
rect 26970 9052 26976 9104
rect 27028 9092 27034 9104
rect 27433 9095 27491 9101
rect 27433 9092 27445 9095
rect 27028 9064 27445 9092
rect 27028 9052 27034 9064
rect 27433 9061 27445 9064
rect 27479 9061 27491 9095
rect 27433 9055 27491 9061
rect 27706 9052 27712 9104
rect 27764 9052 27770 9104
rect 27982 9052 27988 9104
rect 28040 9092 28046 9104
rect 28629 9095 28687 9101
rect 28629 9092 28641 9095
rect 28040 9064 28641 9092
rect 28040 9052 28046 9064
rect 28629 9061 28641 9064
rect 28675 9061 28687 9095
rect 28994 9092 29000 9104
rect 28955 9064 29000 9092
rect 28629 9055 28687 9061
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 18288 8996 18613 9024
rect 18288 8984 18294 8996
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 9024 19211 9027
rect 19794 9024 19800 9036
rect 19199 8996 19800 9024
rect 19199 8993 19211 8996
rect 19153 8987 19211 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2682 8956 2688 8968
rect 2547 8928 2688 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4430 8956 4436 8968
rect 4391 8928 4436 8956
rect 4157 8919 4215 8925
rect 4172 8888 4200 8919
rect 4430 8916 4436 8928
rect 4488 8956 4494 8968
rect 5074 8956 5080 8968
rect 4488 8928 5080 8956
rect 4488 8916 4494 8928
rect 5074 8916 5080 8928
rect 5132 8956 5138 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5132 8928 5181 8956
rect 5132 8916 5138 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 5169 8919 5227 8925
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7558 8956 7564 8968
rect 7519 8928 7564 8956
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 11698 8956 11704 8968
rect 11659 8928 11704 8956
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13538 8916 13544 8928
rect 13596 8956 13602 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 13596 8928 16865 8956
rect 13596 8916 13602 8928
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 16899 8928 17141 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8925 17463 8959
rect 18616 8956 18644 8987
rect 19794 8984 19800 8996
rect 19852 9024 19858 9036
rect 20806 9024 20812 9036
rect 19852 8996 20812 9024
rect 19852 8984 19858 8996
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 22830 9033 22836 9036
rect 22808 9027 22836 9033
rect 22808 8993 22820 9027
rect 22808 8987 22836 8993
rect 22823 8984 22836 8987
rect 22888 8984 22894 9036
rect 23820 9027 23878 9033
rect 23820 8993 23832 9027
rect 23866 9024 23878 9027
rect 23934 9024 23940 9036
rect 23866 8996 23940 9024
rect 23866 8993 23878 8996
rect 23820 8987 23878 8993
rect 23934 8984 23940 8996
rect 23992 9024 23998 9036
rect 24854 9024 24860 9036
rect 23992 8996 24716 9024
rect 24767 8996 24860 9024
rect 23992 8984 23998 8996
rect 19242 8956 19248 8968
rect 18616 8928 19248 8956
rect 17405 8919 17463 8925
rect 4522 8888 4528 8900
rect 4172 8860 4528 8888
rect 4522 8848 4528 8860
rect 4580 8888 4586 8900
rect 5442 8888 5448 8900
rect 4580 8860 5448 8888
rect 4580 8848 4586 8860
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 5721 8891 5779 8897
rect 5721 8857 5733 8891
rect 5767 8888 5779 8891
rect 5994 8888 6000 8900
rect 5767 8860 6000 8888
rect 5767 8857 5779 8860
rect 5721 8851 5779 8857
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 8444 8860 8493 8888
rect 8444 8848 8450 8860
rect 8481 8857 8493 8860
rect 8527 8888 8539 8891
rect 8754 8888 8760 8900
rect 8527 8860 8760 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 12250 8888 12256 8900
rect 12211 8860 12256 8888
rect 12250 8848 12256 8860
rect 12308 8848 12314 8900
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 17420 8888 17448 8919
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 22823 8956 22851 8984
rect 19392 8928 22851 8956
rect 19392 8916 19398 8928
rect 21818 8888 21824 8900
rect 16724 8860 17448 8888
rect 21779 8860 21824 8888
rect 16724 8848 16730 8860
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 24688 8888 24716 8996
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 24946 8984 24952 9036
rect 25004 9024 25010 9036
rect 25317 9027 25375 9033
rect 25317 9024 25329 9027
rect 25004 8996 25329 9024
rect 25004 8984 25010 8996
rect 25317 8993 25329 8996
rect 25363 8993 25375 9027
rect 25317 8987 25375 8993
rect 24872 8956 24900 8984
rect 25406 8956 25412 8968
rect 24872 8928 25412 8956
rect 25406 8916 25412 8928
rect 25464 8916 25470 8968
rect 25590 8956 25596 8968
rect 25551 8928 25596 8956
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 27341 8959 27399 8965
rect 27341 8925 27353 8959
rect 27387 8956 27399 8959
rect 27614 8956 27620 8968
rect 27387 8928 27620 8956
rect 27387 8925 27399 8928
rect 27341 8919 27399 8925
rect 27614 8916 27620 8928
rect 27672 8916 27678 8968
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8956 28043 8959
rect 28074 8956 28080 8968
rect 28031 8928 28080 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 28074 8916 28080 8928
rect 28132 8956 28138 8968
rect 28534 8956 28540 8968
rect 28132 8928 28540 8956
rect 28132 8916 28138 8928
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 28644 8956 28672 9055
rect 28994 9052 29000 9064
rect 29052 9052 29058 9104
rect 34054 9092 34060 9104
rect 34015 9064 34060 9092
rect 34054 9052 34060 9064
rect 34112 9052 34118 9104
rect 35618 9092 35624 9104
rect 35579 9064 35624 9092
rect 35618 9052 35624 9064
rect 35676 9052 35682 9104
rect 30374 8984 30380 9036
rect 30432 9033 30438 9036
rect 30432 9027 30470 9033
rect 30458 8993 30470 9027
rect 32306 9024 32312 9036
rect 32267 8996 32312 9024
rect 30432 8987 30470 8993
rect 30432 8984 30438 8987
rect 32306 8984 32312 8996
rect 32364 8984 32370 9036
rect 32677 9027 32735 9033
rect 32677 8993 32689 9027
rect 32723 9024 32735 9027
rect 32766 9024 32772 9036
rect 32723 8996 32772 9024
rect 32723 8993 32735 8996
rect 32677 8987 32735 8993
rect 32766 8984 32772 8996
rect 32824 8984 32830 9036
rect 28905 8959 28963 8965
rect 28905 8956 28917 8959
rect 28644 8928 28917 8956
rect 28905 8925 28917 8928
rect 28951 8925 28963 8959
rect 29178 8956 29184 8968
rect 29139 8928 29184 8956
rect 28905 8919 28963 8925
rect 29178 8916 29184 8928
rect 29236 8916 29242 8968
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 32950 8956 32956 8968
rect 32907 8928 32956 8956
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 32950 8916 32956 8928
rect 33008 8916 33014 8968
rect 33318 8916 33324 8968
rect 33376 8956 33382 8968
rect 33965 8959 34023 8965
rect 33965 8956 33977 8959
rect 33376 8928 33977 8956
rect 33376 8916 33382 8928
rect 33965 8925 33977 8928
rect 34011 8956 34023 8959
rect 34146 8956 34152 8968
rect 34011 8928 34152 8956
rect 34011 8925 34023 8928
rect 33965 8919 34023 8925
rect 34146 8916 34152 8928
rect 34204 8916 34210 8968
rect 34241 8959 34299 8965
rect 34241 8925 34253 8959
rect 34287 8925 34299 8959
rect 34241 8919 34299 8925
rect 29822 8888 29828 8900
rect 24688 8860 29828 8888
rect 29822 8848 29828 8860
rect 29880 8848 29886 8900
rect 33870 8848 33876 8900
rect 33928 8888 33934 8900
rect 34256 8888 34284 8919
rect 34330 8916 34336 8968
rect 34388 8956 34394 8968
rect 35529 8959 35587 8965
rect 35529 8956 35541 8959
rect 34388 8928 35541 8956
rect 34388 8916 34394 8928
rect 35529 8925 35541 8928
rect 35575 8956 35587 8959
rect 36262 8956 36268 8968
rect 35575 8928 36268 8956
rect 35575 8925 35587 8928
rect 35529 8919 35587 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 33928 8860 34284 8888
rect 36081 8891 36139 8897
rect 33928 8848 33934 8860
rect 36081 8857 36093 8891
rect 36127 8888 36139 8891
rect 36722 8888 36728 8900
rect 36127 8860 36728 8888
rect 36127 8857 36139 8860
rect 36081 8851 36139 8857
rect 36722 8848 36728 8860
rect 36780 8848 36786 8900
rect 1486 8780 1492 8832
rect 1544 8829 1550 8832
rect 1544 8823 1593 8829
rect 1544 8789 1547 8823
rect 1581 8789 1593 8823
rect 2314 8820 2320 8832
rect 2275 8792 2320 8820
rect 1544 8783 1593 8789
rect 1544 8780 1550 8783
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 3510 8820 3516 8832
rect 3471 8792 3516 8820
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8846 8820 8852 8832
rect 8807 8792 8852 8820
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19705 8823 19763 8829
rect 19705 8820 19717 8823
rect 19576 8792 19717 8820
rect 19576 8780 19582 8792
rect 19705 8789 19717 8792
rect 19751 8820 19763 8823
rect 19794 8820 19800 8832
rect 19751 8792 19800 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 21450 8780 21456 8832
rect 21508 8820 21514 8832
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 21508 8792 22293 8820
rect 21508 8780 21514 8792
rect 22281 8789 22293 8792
rect 22327 8820 22339 8823
rect 22879 8823 22937 8829
rect 22879 8820 22891 8823
rect 22327 8792 22891 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 22879 8789 22891 8792
rect 22925 8789 22937 8823
rect 22879 8783 22937 8789
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 24397 8823 24455 8829
rect 24397 8820 24409 8823
rect 24176 8792 24409 8820
rect 24176 8780 24182 8792
rect 24397 8789 24409 8792
rect 24443 8789 24455 8823
rect 24397 8783 24455 8789
rect 27157 8823 27215 8829
rect 27157 8789 27169 8823
rect 27203 8820 27215 8823
rect 27522 8820 27528 8832
rect 27203 8792 27528 8820
rect 27203 8789 27215 8792
rect 27157 8783 27215 8789
rect 27522 8780 27528 8792
rect 27580 8780 27586 8832
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 28074 8820 28080 8832
rect 27672 8792 28080 8820
rect 27672 8780 27678 8792
rect 28074 8780 28080 8792
rect 28132 8820 28138 8832
rect 30558 8829 30564 8832
rect 28445 8823 28503 8829
rect 28445 8820 28457 8823
rect 28132 8792 28457 8820
rect 28132 8780 28138 8792
rect 28445 8789 28457 8792
rect 28491 8789 28503 8823
rect 28445 8783 28503 8789
rect 30515 8823 30564 8829
rect 30515 8789 30527 8823
rect 30561 8789 30564 8823
rect 30515 8783 30564 8789
rect 30558 8780 30564 8783
rect 30616 8780 30622 8832
rect 31297 8823 31355 8829
rect 31297 8789 31309 8823
rect 31343 8820 31355 8823
rect 31386 8820 31392 8832
rect 31343 8792 31392 8820
rect 31343 8789 31355 8792
rect 31297 8783 31355 8789
rect 31386 8780 31392 8792
rect 31444 8780 31450 8832
rect 33318 8820 33324 8832
rect 33279 8792 33324 8820
rect 33318 8780 33324 8792
rect 33376 8780 33382 8832
rect 34974 8820 34980 8832
rect 34935 8792 34980 8820
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 3200 8588 4169 8616
rect 3200 8576 3206 8588
rect 4157 8585 4169 8588
rect 4203 8616 4215 8619
rect 4246 8616 4252 8628
rect 4203 8588 4252 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 4522 8616 4528 8628
rect 4483 8588 4528 8616
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 5684 8588 6193 8616
rect 5684 8576 5690 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6181 8579 6239 8585
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 8018 8616 8024 8628
rect 7432 8588 8024 8616
rect 7432 8576 7438 8588
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12894 8616 12900 8628
rect 12676 8588 12900 8616
rect 12676 8576 12682 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 17126 8625 17132 8628
rect 17083 8619 17132 8625
rect 17083 8585 17095 8619
rect 17129 8585 17132 8619
rect 17083 8579 17132 8585
rect 17126 8576 17132 8579
rect 17184 8576 17190 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18506 8616 18512 8628
rect 17911 8588 18512 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 19242 8616 19248 8628
rect 19203 8588 19248 8616
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 21324 8588 22385 8616
rect 21324 8576 21330 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22830 8616 22836 8628
rect 22791 8588 22836 8616
rect 22373 8579 22431 8585
rect 22830 8576 22836 8588
rect 22888 8576 22894 8628
rect 23934 8616 23940 8628
rect 23895 8588 23940 8616
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 26789 8619 26847 8625
rect 26789 8585 26801 8619
rect 26835 8616 26847 8619
rect 27798 8616 27804 8628
rect 26835 8588 27804 8616
rect 26835 8585 26847 8588
rect 26789 8579 26847 8585
rect 27798 8576 27804 8588
rect 27856 8616 27862 8628
rect 28721 8619 28779 8625
rect 28721 8616 28733 8619
rect 27856 8588 28733 8616
rect 27856 8576 27862 8588
rect 28721 8585 28733 8588
rect 28767 8616 28779 8619
rect 28994 8616 29000 8628
rect 28767 8588 29000 8616
rect 28767 8585 28779 8588
rect 28721 8579 28779 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 34054 8576 34060 8628
rect 34112 8616 34118 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 34112 8588 34253 8616
rect 34112 8576 34118 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 34425 8619 34483 8625
rect 34425 8585 34437 8619
rect 34471 8616 34483 8619
rect 35618 8616 35624 8628
rect 34471 8588 35624 8616
rect 34471 8585 34483 8588
rect 34425 8579 34483 8585
rect 35618 8576 35624 8588
rect 35676 8616 35682 8628
rect 35897 8619 35955 8625
rect 35897 8616 35909 8619
rect 35676 8588 35909 8616
rect 35676 8576 35682 8588
rect 35897 8585 35909 8588
rect 35943 8585 35955 8619
rect 36262 8616 36268 8628
rect 36223 8588 36268 8616
rect 35897 8579 35955 8585
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 36630 8616 36636 8628
rect 36591 8588 36636 8616
rect 36630 8576 36636 8588
rect 36688 8576 36694 8628
rect 2406 8548 2412 8560
rect 2367 8520 2412 8548
rect 2406 8508 2412 8520
rect 2464 8548 2470 8560
rect 3878 8548 3884 8560
rect 2464 8520 3884 8548
rect 2464 8508 2470 8520
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 4985 8551 5043 8557
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5810 8548 5816 8560
rect 5031 8520 5672 8548
rect 5771 8520 5816 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 1946 8480 1952 8492
rect 1535 8452 1952 8480
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 5132 8452 5273 8480
rect 5132 8440 5138 8452
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5644 8480 5672 8520
rect 5810 8508 5816 8520
rect 5868 8508 5874 8560
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 8297 8551 8355 8557
rect 8297 8548 8309 8551
rect 7340 8520 8309 8548
rect 7340 8508 7346 8520
rect 8297 8517 8309 8520
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 5994 8480 6000 8492
rect 5644 8452 6000 8480
rect 5261 8443 5319 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 8680 8480 8708 8576
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 10413 8551 10471 8557
rect 10413 8548 10425 8551
rect 10100 8520 10425 8548
rect 10100 8508 10106 8520
rect 10413 8517 10425 8520
rect 10459 8517 10471 8551
rect 10413 8511 10471 8517
rect 11425 8551 11483 8557
rect 11425 8517 11437 8551
rect 11471 8548 11483 8551
rect 12250 8548 12256 8560
rect 11471 8520 12256 8548
rect 11471 8517 11483 8520
rect 11425 8511 11483 8517
rect 12250 8508 12256 8520
rect 12308 8548 12314 8560
rect 12308 8520 12848 8548
rect 12308 8508 12314 8520
rect 10873 8483 10931 8489
rect 8680 8452 9352 8480
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7147 8384 8156 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2866 8344 2872 8356
rect 1627 8316 2872 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 3200 8316 3245 8344
rect 3200 8304 3206 8316
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 7422 8347 7480 8353
rect 7422 8344 7434 8347
rect 5408 8316 5453 8344
rect 7300 8316 7434 8344
rect 5408 8304 5414 8316
rect 7300 8288 7328 8316
rect 7422 8313 7434 8316
rect 7468 8313 7480 8347
rect 8128 8344 8156 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 8846 8412 8852 8424
rect 8720 8384 8852 8412
rect 8720 8372 8726 8384
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9324 8421 9352 8452
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11330 8480 11336 8492
rect 10919 8452 11336 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12820 8489 12848 8520
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13320 8520 13829 8548
rect 13320 8508 13326 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 15105 8551 15163 8557
rect 15105 8517 15117 8551
rect 15151 8548 15163 8551
rect 15378 8548 15384 8560
rect 15151 8520 15384 8548
rect 15151 8517 15163 8520
rect 15105 8511 15163 8517
rect 15378 8508 15384 8520
rect 15436 8548 15442 8560
rect 16485 8551 16543 8557
rect 16485 8548 16497 8551
rect 15436 8520 16497 8548
rect 15436 8508 15442 8520
rect 16485 8517 16497 8520
rect 16531 8548 16543 8551
rect 16942 8548 16948 8560
rect 16531 8520 16948 8548
rect 16531 8517 16543 8520
rect 16485 8511 16543 8517
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 18877 8551 18935 8557
rect 18877 8548 18889 8551
rect 18012 8520 18889 8548
rect 18012 8508 18018 8520
rect 18877 8517 18889 8520
rect 18923 8548 18935 8551
rect 18966 8548 18972 8560
rect 18923 8520 18972 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 18966 8508 18972 8520
rect 19024 8508 19030 8560
rect 19260 8548 19288 8576
rect 23566 8548 23572 8560
rect 19260 8520 23572 8548
rect 23566 8508 23572 8520
rect 23624 8508 23630 8560
rect 29178 8508 29184 8560
rect 29236 8548 29242 8560
rect 33870 8548 33876 8560
rect 29236 8520 29684 8548
rect 33831 8520 33876 8548
rect 29236 8508 29242 8520
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13722 8480 13728 8492
rect 12851 8452 13728 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14700 8452 14872 8480
rect 14700 8440 14706 8452
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 14052 8415 14110 8421
rect 14052 8381 14064 8415
rect 14098 8412 14110 8415
rect 14553 8415 14611 8421
rect 14553 8412 14565 8415
rect 14098 8384 14565 8412
rect 14098 8381 14110 8384
rect 14052 8375 14110 8381
rect 14553 8381 14565 8384
rect 14599 8412 14611 8415
rect 14734 8412 14740 8424
rect 14599 8384 14740 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 10962 8344 10968 8356
rect 8128 8316 8984 8344
rect 10923 8316 10968 8344
rect 7422 8307 7480 8313
rect 8956 8288 8984 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11882 8344 11888 8356
rect 11843 8316 11888 8344
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8344 12679 8347
rect 14139 8347 14197 8353
rect 12667 8316 12701 8344
rect 12667 8313 12679 8316
rect 12621 8307 12679 8313
rect 14139 8313 14151 8347
rect 14185 8344 14197 8347
rect 14642 8344 14648 8356
rect 14185 8316 14648 8344
rect 14185 8313 14197 8316
rect 14139 8307 14197 8313
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3786 8276 3792 8288
rect 2832 8248 3792 8276
rect 2832 8236 2838 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 7282 8276 7288 8288
rect 6687 8248 7288 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8938 8276 8944 8288
rect 8899 8248 8944 8276
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12636 8276 12664 8307
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 14844 8344 14872 8452
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 15197 8483 15255 8489
rect 15197 8480 15209 8483
rect 14976 8452 15209 8480
rect 14976 8440 14982 8452
rect 15197 8449 15209 8452
rect 15243 8480 15255 8483
rect 16761 8483 16819 8489
rect 16761 8480 16773 8483
rect 15243 8452 16773 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 16761 8449 16773 8452
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 19702 8480 19708 8492
rect 18371 8452 19708 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20070 8480 20076 8492
rect 19935 8452 20076 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 21450 8480 21456 8492
rect 21411 8452 21456 8480
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 21818 8480 21824 8492
rect 21779 8452 21824 8480
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 27706 8480 27712 8492
rect 27667 8452 27712 8480
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8480 29423 8483
rect 29454 8480 29460 8492
rect 29411 8452 29460 8480
rect 29411 8449 29423 8452
rect 29365 8443 29423 8449
rect 29454 8440 29460 8452
rect 29512 8440 29518 8492
rect 29656 8489 29684 8520
rect 33870 8508 33876 8520
rect 33928 8548 33934 8560
rect 35526 8548 35532 8560
rect 33928 8520 35532 8548
rect 33928 8508 33934 8520
rect 35526 8508 35532 8520
rect 35584 8508 35590 8560
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8449 29699 8483
rect 29641 8443 29699 8449
rect 33321 8483 33379 8489
rect 33321 8449 33333 8483
rect 33367 8480 33379 8483
rect 33594 8480 33600 8492
rect 33367 8452 33600 8480
rect 33367 8449 33379 8452
rect 33321 8443 33379 8449
rect 33594 8440 33600 8452
rect 33652 8440 33658 8492
rect 34974 8480 34980 8492
rect 34887 8452 34980 8480
rect 34974 8440 34980 8452
rect 35032 8480 35038 8492
rect 37691 8483 37749 8489
rect 37691 8480 37703 8483
rect 35032 8452 37703 8480
rect 35032 8440 35038 8452
rect 37691 8449 37703 8452
rect 37737 8449 37749 8483
rect 37691 8443 37749 8449
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 16980 8415 17038 8421
rect 16980 8412 16992 8415
rect 16908 8384 16992 8412
rect 16908 8372 16914 8384
rect 16980 8381 16992 8384
rect 17026 8381 17038 8415
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 16980 8375 17038 8381
rect 20640 8384 21189 8412
rect 14918 8344 14924 8356
rect 14844 8316 14924 8344
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 15518 8347 15576 8353
rect 15518 8344 15530 8347
rect 15436 8316 15530 8344
rect 15436 8304 15442 8316
rect 15518 8313 15530 8316
rect 15564 8313 15576 8347
rect 17218 8344 17224 8356
rect 15518 8307 15576 8313
rect 16592 8316 17224 8344
rect 12894 8276 12900 8288
rect 12299 8248 12900 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 16114 8276 16120 8288
rect 16075 8248 16120 8276
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 16482 8236 16488 8288
rect 16540 8276 16546 8288
rect 16592 8276 16620 8316
rect 17218 8304 17224 8316
rect 17276 8344 17282 8356
rect 17405 8347 17463 8353
rect 17405 8344 17417 8347
rect 17276 8316 17417 8344
rect 17276 8304 17282 8316
rect 17405 8313 17417 8316
rect 17451 8313 17463 8347
rect 17405 8307 17463 8313
rect 18417 8347 18475 8353
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 18506 8344 18512 8356
rect 18463 8316 18512 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 19613 8347 19671 8353
rect 19613 8344 19625 8347
rect 19392 8316 19625 8344
rect 19392 8304 19398 8316
rect 19613 8313 19625 8316
rect 19659 8344 19671 8347
rect 19981 8347 20039 8353
rect 19981 8344 19993 8347
rect 19659 8316 19993 8344
rect 19659 8313 19671 8316
rect 19613 8307 19671 8313
rect 19981 8313 19993 8316
rect 20027 8344 20039 8347
rect 20027 8316 20484 8344
rect 20027 8313 20039 8316
rect 19981 8307 20039 8313
rect 16540 8248 16620 8276
rect 20456 8276 20484 8316
rect 20640 8276 20668 8384
rect 21177 8381 21189 8384
rect 21223 8412 21235 8415
rect 21266 8412 21272 8424
rect 21223 8384 21272 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 24394 8412 24400 8424
rect 24355 8384 24400 8412
rect 24394 8372 24400 8384
rect 24452 8372 24458 8424
rect 24857 8415 24915 8421
rect 24857 8381 24869 8415
rect 24903 8412 24915 8415
rect 24946 8412 24952 8424
rect 24903 8384 24952 8412
rect 24903 8381 24915 8384
rect 24857 8375 24915 8381
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 20809 8347 20867 8353
rect 20809 8344 20821 8347
rect 20772 8316 20821 8344
rect 20772 8304 20778 8316
rect 20809 8313 20821 8316
rect 20855 8344 20867 8347
rect 21542 8344 21548 8356
rect 20855 8316 21548 8344
rect 20855 8313 20867 8316
rect 20809 8307 20867 8313
rect 21542 8304 21548 8316
rect 21600 8304 21606 8356
rect 23477 8347 23535 8353
rect 23477 8313 23489 8347
rect 23523 8344 23535 8347
rect 24872 8344 24900 8375
rect 24946 8372 24952 8384
rect 25004 8372 25010 8424
rect 25041 8415 25099 8421
rect 25041 8381 25053 8415
rect 25087 8412 25099 8415
rect 25866 8412 25872 8424
rect 25087 8384 25872 8412
rect 25087 8381 25099 8384
rect 25041 8375 25099 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8412 31263 8415
rect 31386 8412 31392 8424
rect 31251 8384 31392 8412
rect 31251 8381 31263 8384
rect 31205 8375 31263 8381
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 32125 8415 32183 8421
rect 32125 8381 32137 8415
rect 32171 8412 32183 8415
rect 32171 8384 33180 8412
rect 32171 8381 32183 8384
rect 32125 8375 32183 8381
rect 25406 8344 25412 8356
rect 23523 8316 24900 8344
rect 25367 8316 25412 8344
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 25406 8304 25412 8316
rect 25464 8304 25470 8356
rect 26231 8347 26289 8353
rect 26231 8313 26243 8347
rect 26277 8313 26289 8347
rect 27798 8344 27804 8356
rect 27759 8316 27804 8344
rect 26231 8307 26289 8313
rect 20456 8248 20668 8276
rect 25777 8279 25835 8285
rect 16540 8236 16546 8248
rect 25777 8245 25789 8279
rect 25823 8276 25835 8279
rect 26252 8276 26280 8307
rect 27798 8304 27804 8316
rect 27856 8344 27862 8356
rect 27982 8344 27988 8356
rect 27856 8316 27988 8344
rect 27856 8304 27862 8316
rect 27982 8304 27988 8316
rect 28040 8304 28046 8356
rect 28353 8347 28411 8353
rect 28353 8313 28365 8347
rect 28399 8344 28411 8347
rect 28534 8344 28540 8356
rect 28399 8316 28540 8344
rect 28399 8313 28411 8316
rect 28353 8307 28411 8313
rect 28534 8304 28540 8316
rect 28592 8304 28598 8356
rect 28997 8347 29055 8353
rect 28997 8344 29009 8347
rect 28828 8316 29009 8344
rect 26786 8276 26792 8288
rect 25823 8248 26792 8276
rect 25823 8245 25835 8248
rect 25777 8239 25835 8245
rect 26786 8236 26792 8248
rect 26844 8236 26850 8288
rect 26970 8236 26976 8288
rect 27028 8276 27034 8288
rect 27249 8279 27307 8285
rect 27249 8276 27261 8279
rect 27028 8248 27261 8276
rect 27028 8236 27034 8248
rect 27249 8245 27261 8248
rect 27295 8276 27307 8279
rect 28828 8276 28856 8316
rect 28997 8313 29009 8316
rect 29043 8344 29055 8347
rect 29457 8347 29515 8353
rect 29457 8344 29469 8347
rect 29043 8316 29469 8344
rect 29043 8313 29055 8316
rect 28997 8307 29055 8313
rect 29457 8313 29469 8316
rect 29503 8313 29515 8347
rect 30374 8344 30380 8356
rect 30335 8316 30380 8344
rect 29457 8307 29515 8313
rect 30374 8304 30380 8316
rect 30432 8304 30438 8356
rect 31526 8347 31584 8353
rect 31526 8313 31538 8347
rect 31572 8344 31584 8347
rect 31572 8316 31606 8344
rect 31572 8313 31584 8316
rect 31526 8307 31584 8313
rect 27295 8248 28856 8276
rect 31113 8279 31171 8285
rect 27295 8245 27307 8248
rect 27249 8239 27307 8245
rect 31113 8245 31125 8279
rect 31159 8276 31171 8279
rect 31541 8276 31569 8307
rect 32306 8304 32312 8356
rect 32364 8344 32370 8356
rect 32401 8347 32459 8353
rect 32401 8344 32413 8347
rect 32364 8316 32413 8344
rect 32364 8304 32370 8316
rect 32401 8313 32413 8316
rect 32447 8313 32459 8347
rect 32766 8344 32772 8356
rect 32727 8316 32772 8344
rect 32401 8307 32459 8313
rect 32766 8304 32772 8316
rect 32824 8304 32830 8356
rect 33152 8344 33180 8384
rect 36262 8372 36268 8424
rect 36320 8412 36326 8424
rect 36449 8415 36507 8421
rect 36449 8412 36461 8415
rect 36320 8384 36461 8412
rect 36320 8372 36326 8384
rect 36449 8381 36461 8384
rect 36495 8412 36507 8415
rect 37001 8415 37059 8421
rect 37001 8412 37013 8415
rect 36495 8384 37013 8412
rect 36495 8381 36507 8384
rect 36449 8375 36507 8381
rect 37001 8381 37013 8384
rect 37047 8381 37059 8415
rect 37588 8415 37646 8421
rect 37588 8412 37600 8415
rect 37001 8375 37059 8381
rect 37108 8384 37600 8412
rect 33318 8344 33324 8356
rect 33152 8316 33324 8344
rect 33318 8304 33324 8316
rect 33376 8344 33382 8356
rect 33413 8347 33471 8353
rect 33413 8344 33425 8347
rect 33376 8316 33425 8344
rect 33376 8304 33382 8316
rect 33413 8313 33425 8316
rect 33459 8344 33471 8347
rect 34425 8347 34483 8353
rect 34425 8344 34437 8347
rect 33459 8316 34437 8344
rect 33459 8313 33471 8316
rect 33413 8307 33471 8313
rect 34425 8313 34437 8316
rect 34471 8313 34483 8347
rect 34425 8307 34483 8313
rect 34606 8304 34612 8356
rect 34664 8344 34670 8356
rect 34701 8347 34759 8353
rect 34701 8344 34713 8347
rect 34664 8316 34713 8344
rect 34664 8304 34670 8316
rect 34701 8313 34713 8316
rect 34747 8344 34759 8347
rect 35069 8347 35127 8353
rect 35069 8344 35081 8347
rect 34747 8316 35081 8344
rect 34747 8313 34759 8316
rect 34701 8307 34759 8313
rect 35069 8313 35081 8316
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 32214 8276 32220 8288
rect 31159 8248 32220 8276
rect 31159 8245 31171 8248
rect 31113 8239 31171 8245
rect 32214 8236 32220 8248
rect 32272 8236 32278 8288
rect 33962 8236 33968 8288
rect 34020 8276 34026 8288
rect 37108 8276 37136 8384
rect 37588 8381 37600 8384
rect 37634 8412 37646 8415
rect 38010 8412 38016 8424
rect 37634 8384 38016 8412
rect 37634 8381 37646 8384
rect 37588 8375 37646 8381
rect 38010 8372 38016 8384
rect 38068 8372 38074 8424
rect 34020 8248 37136 8276
rect 34020 8236 34026 8248
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 2682 8072 2688 8084
rect 2087 8044 2688 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3142 8072 3148 8084
rect 3099 8044 3148 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3142 8032 3148 8044
rect 3200 8072 3206 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 3200 8044 3341 8072
rect 3200 8032 3206 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3329 8035 3387 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 6822 8072 6828 8084
rect 6687 8044 6828 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 2498 8013 2504 8016
rect 2495 8004 2504 8013
rect 2459 7976 2504 8004
rect 2495 7967 2504 7976
rect 2498 7964 2504 7967
rect 2556 7964 2562 8016
rect 4154 8004 4160 8016
rect 4115 7976 4160 8004
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 4246 7964 4252 8016
rect 4304 8004 4310 8016
rect 4801 8007 4859 8013
rect 4304 7976 4349 8004
rect 4304 7964 4310 7976
rect 4801 7973 4813 8007
rect 4847 8004 4859 8007
rect 5074 8004 5080 8016
rect 4847 7976 5080 8004
rect 4847 7973 4859 7976
rect 4801 7967 4859 7973
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2222 7936 2228 7948
rect 2179 7908 2228 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5629 7939 5687 7945
rect 5629 7936 5641 7939
rect 5500 7908 5641 7936
rect 5500 7896 5506 7908
rect 5629 7905 5641 7908
rect 5675 7936 5687 7939
rect 6454 7936 6460 7948
rect 5675 7908 6460 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 6748 7945 6776 8044
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 6972 8044 7665 8072
rect 6972 8032 6978 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 7653 8035 7711 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8938 8072 8944 8084
rect 8435 8044 8944 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10594 8072 10600 8084
rect 10551 8044 10600 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 10962 8072 10968 8084
rect 10919 8044 10968 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 10962 8032 10968 8044
rect 11020 8072 11026 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11020 8044 11897 8072
rect 11020 8032 11026 8044
rect 11885 8041 11897 8044
rect 11931 8072 11943 8075
rect 12342 8072 12348 8084
rect 11931 8044 12348 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 16209 8075 16267 8081
rect 15436 8044 15694 8072
rect 15436 8032 15442 8044
rect 7095 8007 7153 8013
rect 7095 7973 7107 8007
rect 7141 8004 7153 8007
rect 7282 8004 7288 8016
rect 7141 7976 7288 8004
rect 7141 7973 7153 7976
rect 7095 7967 7153 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 8444 7908 8493 7936
rect 8444 7896 8450 7908
rect 8481 7905 8493 7908
rect 8527 7905 8539 7939
rect 8481 7899 8539 7905
rect 9950 7896 9956 7948
rect 10008 7945 10014 7948
rect 10008 7939 10046 7945
rect 10034 7905 10046 7939
rect 10612 7936 10640 8032
rect 11327 8007 11385 8013
rect 11327 7973 11339 8007
rect 11373 8004 11385 8007
rect 11974 8004 11980 8016
rect 11373 7976 11980 8004
rect 11373 7973 11385 7976
rect 11327 7967 11385 7973
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 12894 8004 12900 8016
rect 12855 7976 12900 8004
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 15666 8013 15694 8044
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16482 8072 16488 8084
rect 16255 8044 16488 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19760 8044 19809 8072
rect 19760 8032 19766 8044
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 19797 8035 19855 8041
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 22097 8075 22155 8081
rect 22097 8072 22109 8075
rect 22060 8044 22109 8072
rect 22060 8032 22066 8044
rect 22097 8041 22109 8044
rect 22143 8041 22155 8075
rect 23658 8072 23664 8084
rect 23619 8044 23664 8072
rect 22097 8035 22155 8041
rect 23658 8032 23664 8044
rect 23716 8032 23722 8084
rect 25866 8072 25872 8084
rect 25827 8044 25872 8072
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 27430 8072 27436 8084
rect 27391 8044 27436 8072
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 27801 8075 27859 8081
rect 27801 8041 27813 8075
rect 27847 8072 27859 8075
rect 27982 8072 27988 8084
rect 27847 8044 27988 8072
rect 27847 8041 27859 8044
rect 27801 8035 27859 8041
rect 27982 8032 27988 8044
rect 28040 8032 28046 8084
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 33413 8075 33471 8081
rect 28132 8044 28177 8072
rect 28132 8032 28138 8044
rect 33413 8041 33425 8075
rect 33459 8072 33471 8075
rect 33502 8072 33508 8084
rect 33459 8044 33508 8072
rect 33459 8041 33471 8044
rect 33413 8035 33471 8041
rect 33502 8032 33508 8044
rect 33560 8032 33566 8084
rect 34146 8032 34152 8084
rect 34204 8072 34210 8084
rect 34333 8075 34391 8081
rect 34333 8072 34345 8075
rect 34204 8044 34345 8072
rect 34204 8032 34210 8044
rect 34333 8041 34345 8044
rect 34379 8041 34391 8075
rect 34333 8035 34391 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35897 8075 35955 8081
rect 35897 8072 35909 8075
rect 35584 8044 35909 8072
rect 35584 8032 35590 8044
rect 35897 8041 35909 8044
rect 35943 8041 35955 8075
rect 36630 8072 36636 8084
rect 36591 8044 36636 8072
rect 35897 8035 35955 8041
rect 36630 8032 36636 8044
rect 36688 8032 36694 8084
rect 15630 8007 15694 8013
rect 15630 7973 15642 8007
rect 15676 7976 15694 8007
rect 15676 7973 15688 7976
rect 15630 7967 15688 7973
rect 17126 7964 17132 8016
rect 17184 8004 17190 8016
rect 17221 8007 17279 8013
rect 17221 8004 17233 8007
rect 17184 7976 17233 8004
rect 17184 7964 17190 7976
rect 17221 7973 17233 7976
rect 17267 7973 17279 8007
rect 17221 7967 17279 7973
rect 17773 8007 17831 8013
rect 17773 7973 17785 8007
rect 17819 8004 17831 8007
rect 17954 8004 17960 8016
rect 17819 7976 17960 8004
rect 17819 7973 17831 7976
rect 17773 7967 17831 7973
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 18963 8007 19021 8013
rect 18963 7973 18975 8007
rect 19009 8004 19021 8007
rect 19150 8004 19156 8016
rect 19009 7976 19156 8004
rect 19009 7973 19021 7976
rect 18963 7967 19021 7973
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 21266 8004 21272 8016
rect 21227 7976 21272 8004
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 21818 8004 21824 8016
rect 21779 7976 21824 8004
rect 21818 7964 21824 7976
rect 21876 7964 21882 8016
rect 22830 8004 22836 8016
rect 22791 7976 22836 8004
rect 22830 7964 22836 7976
rect 22888 7964 22894 8016
rect 26786 7964 26792 8016
rect 26844 8013 26850 8016
rect 26844 8007 26892 8013
rect 26844 7973 26846 8007
rect 26880 7973 26892 8007
rect 28626 8004 28632 8016
rect 28587 7976 28632 8004
rect 26844 7967 26892 7973
rect 26844 7964 26850 7967
rect 28626 7964 28632 7976
rect 28684 7964 28690 8016
rect 32214 7964 32220 8016
rect 32272 8004 32278 8016
rect 32446 8007 32504 8013
rect 32446 8004 32458 8007
rect 32272 7976 32458 8004
rect 32272 7964 32278 7976
rect 32446 7973 32458 7976
rect 32492 7973 32504 8007
rect 34054 8004 34060 8016
rect 32446 7967 32504 7973
rect 33060 7976 34060 8004
rect 33060 7948 33088 7976
rect 34054 7964 34060 7976
rect 34112 7964 34118 8016
rect 34698 7964 34704 8016
rect 34756 8004 34762 8016
rect 35069 8007 35127 8013
rect 35069 8004 35081 8007
rect 34756 7976 35081 8004
rect 34756 7964 34762 7976
rect 35069 7973 35081 7976
rect 35115 7973 35127 8007
rect 35069 7967 35127 7973
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 10612 7908 10977 7936
rect 10008 7899 10046 7905
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 10008 7896 10014 7899
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 15252 7908 15301 7936
rect 15252 7896 15258 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 18601 7939 18659 7945
rect 18601 7905 18613 7939
rect 18647 7936 18659 7939
rect 18690 7936 18696 7948
rect 18647 7908 18696 7936
rect 18647 7905 18659 7908
rect 18601 7899 18659 7905
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 20714 7936 20720 7948
rect 19567 7908 20720 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 24854 7936 24860 7948
rect 24815 7908 24860 7936
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 25314 7936 25320 7948
rect 25275 7908 25320 7936
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 30742 7936 30748 7948
rect 30703 7908 30748 7936
rect 30742 7896 30748 7908
rect 30800 7896 30806 7948
rect 31021 7939 31079 7945
rect 31021 7905 31033 7939
rect 31067 7936 31079 7939
rect 31294 7936 31300 7948
rect 31067 7908 31300 7936
rect 31067 7905 31079 7908
rect 31021 7899 31079 7905
rect 31294 7896 31300 7908
rect 31352 7896 31358 7948
rect 33042 7936 33048 7948
rect 32955 7908 33048 7936
rect 33042 7896 33048 7908
rect 33100 7896 33106 7948
rect 33870 7896 33876 7948
rect 33928 7945 33934 7948
rect 33928 7939 33966 7945
rect 33954 7905 33966 7939
rect 36446 7936 36452 7948
rect 36407 7908 36452 7936
rect 33928 7899 33966 7905
rect 33928 7896 33934 7899
rect 36446 7896 36452 7908
rect 36504 7896 36510 7948
rect 6270 7868 6276 7880
rect 6231 7840 6276 7868
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 10091 7871 10149 7877
rect 10091 7837 10103 7871
rect 10137 7868 10149 7871
rect 11698 7868 11704 7880
rect 10137 7840 11704 7868
rect 10137 7837 10149 7840
rect 10091 7831 10149 7837
rect 11698 7828 11704 7840
rect 11756 7868 11762 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11756 7840 12173 7868
rect 11756 7828 11762 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12161 7831 12219 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13538 7868 13544 7880
rect 13495 7840 13544 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 16482 7868 16488 7880
rect 16443 7840 16488 7868
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 17494 7868 17500 7880
rect 17175 7840 17500 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 17494 7828 17500 7840
rect 17552 7868 17558 7880
rect 17862 7868 17868 7880
rect 17552 7840 17868 7868
rect 17552 7828 17558 7840
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20732 7840 21189 7868
rect 566 7760 572 7812
rect 624 7800 630 7812
rect 20732 7809 20760 7840
rect 21177 7837 21189 7840
rect 21223 7868 21235 7871
rect 21634 7868 21640 7880
rect 21223 7840 21640 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 22462 7828 22468 7880
rect 22520 7868 22526 7880
rect 22741 7871 22799 7877
rect 22741 7868 22753 7871
rect 22520 7840 22753 7868
rect 22520 7828 22526 7840
rect 22741 7837 22753 7840
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 24026 7868 24032 7880
rect 23431 7840 24032 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 24946 7868 24952 7880
rect 24811 7840 24952 7868
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 24946 7828 24952 7840
rect 25004 7868 25010 7880
rect 25332 7868 25360 7896
rect 25004 7840 25360 7868
rect 25593 7871 25651 7877
rect 25004 7828 25010 7840
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 26513 7871 26571 7877
rect 26513 7868 26525 7871
rect 25639 7840 26525 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 26513 7837 26525 7840
rect 26559 7868 26571 7871
rect 27614 7868 27620 7880
rect 26559 7840 27620 7868
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 28534 7868 28540 7880
rect 28495 7840 28540 7868
rect 28534 7828 28540 7840
rect 28592 7828 28598 7880
rect 29181 7871 29239 7877
rect 29181 7837 29193 7871
rect 29227 7868 29239 7871
rect 29638 7868 29644 7880
rect 29227 7840 29644 7868
rect 29227 7837 29239 7840
rect 29181 7831 29239 7837
rect 29638 7828 29644 7840
rect 29696 7828 29702 7880
rect 31205 7871 31263 7877
rect 31205 7837 31217 7871
rect 31251 7868 31263 7871
rect 32122 7868 32128 7880
rect 31251 7840 32128 7868
rect 31251 7837 31263 7840
rect 31205 7831 31263 7837
rect 32122 7828 32128 7840
rect 32180 7828 32186 7880
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7837 35035 7871
rect 35618 7868 35624 7880
rect 35579 7840 35624 7868
rect 34977 7831 35035 7837
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 624 7772 5825 7800
rect 624 7760 630 7772
rect 5813 7769 5825 7772
rect 5859 7769 5871 7803
rect 5813 7763 5871 7769
rect 20717 7803 20775 7809
rect 20717 7769 20729 7803
rect 20763 7769 20775 7803
rect 34790 7800 34796 7812
rect 34703 7772 34796 7800
rect 20717 7763 20775 7769
rect 34790 7760 34796 7772
rect 34848 7800 34854 7812
rect 34992 7800 35020 7831
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 36722 7800 36728 7812
rect 34848 7772 36728 7800
rect 34848 7760 34854 7772
rect 36722 7760 36728 7772
rect 36780 7760 36786 7812
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 5350 7732 5356 7744
rect 5307 7704 5356 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 8662 7732 8668 7744
rect 8623 7704 8668 7732
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 16850 7732 16856 7744
rect 16811 7704 16856 7732
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18506 7732 18512 7744
rect 18371 7704 18512 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18506 7692 18512 7704
rect 18564 7732 18570 7744
rect 18874 7732 18880 7744
rect 18564 7704 18880 7732
rect 18564 7692 18570 7704
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 23566 7692 23572 7744
rect 23624 7732 23630 7744
rect 24394 7732 24400 7744
rect 23624 7704 24400 7732
rect 23624 7692 23630 7704
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 29454 7732 29460 7744
rect 29415 7704 29460 7732
rect 29454 7692 29460 7704
rect 29512 7692 29518 7744
rect 34011 7735 34069 7741
rect 34011 7701 34023 7735
rect 34057 7732 34069 7735
rect 34146 7732 34152 7744
rect 34057 7704 34152 7732
rect 34057 7701 34069 7704
rect 34011 7695 34069 7701
rect 34146 7692 34152 7704
rect 34204 7692 34210 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3510 7528 3516 7540
rect 3191 7500 3516 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3510 7488 3516 7500
rect 3568 7528 3574 7540
rect 4246 7528 4252 7540
rect 3568 7500 4252 7528
rect 3568 7488 3574 7500
rect 4246 7488 4252 7500
rect 4304 7528 4310 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4304 7500 4905 7528
rect 4304 7488 4310 7500
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 4893 7491 4951 7497
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6454 7528 6460 7540
rect 6319 7500 6460 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 6972 7500 7757 7528
rect 6972 7488 6978 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 12860 7500 13829 7528
rect 12860 7488 12866 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 15378 7528 15384 7540
rect 15339 7500 15384 7528
rect 13817 7491 13875 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 18969 7531 19027 7537
rect 18969 7497 18981 7531
rect 19015 7528 19027 7531
rect 19242 7528 19248 7540
rect 19015 7500 19248 7528
rect 19015 7497 19027 7500
rect 18969 7491 19027 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 20901 7531 20959 7537
rect 20901 7497 20913 7531
rect 20947 7528 20959 7531
rect 21266 7528 21272 7540
rect 20947 7500 21272 7528
rect 20947 7497 20959 7500
rect 20901 7491 20959 7497
rect 21266 7488 21272 7500
rect 21324 7528 21330 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 21324 7500 21465 7528
rect 21324 7488 21330 7500
rect 21453 7497 21465 7500
rect 21499 7528 21511 7531
rect 21545 7531 21603 7537
rect 21545 7528 21557 7531
rect 21499 7500 21557 7528
rect 21499 7497 21511 7500
rect 21453 7491 21511 7497
rect 21545 7497 21557 7500
rect 21591 7497 21603 7531
rect 26970 7528 26976 7540
rect 26931 7500 26976 7528
rect 21545 7491 21603 7497
rect 26970 7488 26976 7500
rect 27028 7488 27034 7540
rect 27614 7528 27620 7540
rect 27575 7500 27620 7528
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 28626 7528 28632 7540
rect 28587 7500 28632 7528
rect 28626 7488 28632 7500
rect 28684 7488 28690 7540
rect 32122 7488 32128 7540
rect 32180 7528 32186 7540
rect 32493 7531 32551 7537
rect 32493 7528 32505 7531
rect 32180 7500 32505 7528
rect 32180 7488 32186 7500
rect 32493 7497 32505 7500
rect 32539 7497 32551 7531
rect 33042 7528 33048 7540
rect 33003 7500 33048 7528
rect 32493 7491 32551 7497
rect 33042 7488 33048 7500
rect 33100 7488 33106 7540
rect 33870 7488 33876 7540
rect 33928 7528 33934 7540
rect 34241 7531 34299 7537
rect 34241 7528 34253 7531
rect 33928 7500 34253 7528
rect 33928 7488 33934 7500
rect 34241 7497 34253 7500
rect 34287 7528 34299 7531
rect 36265 7531 36323 7537
rect 36265 7528 36277 7531
rect 34287 7500 36277 7528
rect 34287 7497 34299 7500
rect 34241 7491 34299 7497
rect 36265 7497 36277 7500
rect 36311 7528 36323 7531
rect 36446 7528 36452 7540
rect 36311 7500 36452 7528
rect 36311 7497 36323 7500
rect 36265 7491 36323 7497
rect 36446 7488 36452 7500
rect 36504 7488 36510 7540
rect 2314 7420 2320 7472
rect 2372 7460 2378 7472
rect 3789 7463 3847 7469
rect 3789 7460 3801 7463
rect 2372 7432 3801 7460
rect 2372 7420 2378 7432
rect 3789 7429 3801 7432
rect 3835 7429 3847 7463
rect 3789 7423 3847 7429
rect 4157 7463 4215 7469
rect 4157 7429 4169 7463
rect 4203 7460 4215 7463
rect 4338 7460 4344 7472
rect 4203 7432 4344 7460
rect 4203 7429 4215 7432
rect 4157 7423 4215 7429
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 7190 7420 7196 7472
rect 7248 7460 7254 7472
rect 8021 7463 8079 7469
rect 8021 7460 8033 7463
rect 7248 7432 8033 7460
rect 7248 7420 7254 7432
rect 8021 7429 8033 7432
rect 8067 7429 8079 7463
rect 8021 7423 8079 7429
rect 11517 7463 11575 7469
rect 11517 7429 11529 7463
rect 11563 7460 11575 7463
rect 12894 7460 12900 7472
rect 11563 7432 12900 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7392 2283 7395
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2271 7364 3525 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 3513 7361 3525 7364
rect 3559 7392 3571 7395
rect 4614 7392 4620 7404
rect 3559 7364 4620 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 5040 7364 5273 7392
rect 5040 7352 5046 7364
rect 5261 7361 5273 7364
rect 5307 7392 5319 7395
rect 5534 7392 5540 7404
rect 5307 7364 5540 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 6822 7392 6828 7404
rect 5684 7364 5729 7392
rect 6783 7364 6828 7392
rect 5684 7352 5690 7364
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 1728 7296 3985 7324
rect 1728 7284 1734 7296
rect 3973 7293 3985 7296
rect 4019 7324 4031 7327
rect 4522 7324 4528 7336
rect 4019 7296 4528 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 8036 7324 8064 7423
rect 12894 7420 12900 7432
rect 12952 7460 12958 7472
rect 13449 7463 13507 7469
rect 13449 7460 13461 7463
rect 12952 7432 13461 7460
rect 12952 7420 12958 7432
rect 13449 7429 13461 7432
rect 13495 7429 13507 7463
rect 13449 7423 13507 7429
rect 21910 7420 21916 7472
rect 21968 7460 21974 7472
rect 22462 7460 22468 7472
rect 21968 7432 22468 7460
rect 21968 7420 21974 7432
rect 22462 7420 22468 7432
rect 22520 7420 22526 7472
rect 23658 7420 23664 7472
rect 23716 7420 23722 7472
rect 27522 7420 27528 7472
rect 27580 7460 27586 7472
rect 27939 7463 27997 7469
rect 27939 7460 27951 7463
rect 27580 7432 27951 7460
rect 27580 7420 27586 7432
rect 27939 7429 27951 7432
rect 27985 7429 27997 7463
rect 35526 7460 35532 7472
rect 27939 7423 27997 7429
rect 34992 7432 35532 7460
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10560 7364 10609 7392
rect 10560 7352 10566 7364
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 15286 7392 15292 7404
rect 14323 7364 15292 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8036 7296 8585 7324
rect 8573 7293 8585 7296
rect 8619 7324 8631 7327
rect 8754 7324 8760 7336
rect 8619 7296 8760 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 8846 7284 8852 7336
rect 8904 7324 8910 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8904 7296 9045 7324
rect 8904 7284 8910 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 9033 7287 9091 7293
rect 12158 7284 12164 7296
rect 12216 7324 12222 7336
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 12216 7296 12541 7324
rect 12216 7284 12222 7296
rect 12529 7293 12541 7296
rect 12575 7293 12587 7327
rect 14550 7324 14556 7336
rect 14511 7296 14556 7324
rect 12529 7287 12587 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 14936 7333 14964 7364
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 16482 7392 16488 7404
rect 16071 7364 16488 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16666 7392 16672 7404
rect 16627 7364 16672 7392
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7392 18107 7395
rect 18138 7392 18144 7404
rect 18095 7364 18144 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19944 7364 19993 7392
rect 19944 7352 19950 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 22002 7392 22008 7404
rect 21867 7364 22008 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 23676 7392 23704 7420
rect 23753 7395 23811 7401
rect 23753 7392 23765 7395
rect 23676 7364 23765 7392
rect 23753 7361 23765 7364
rect 23799 7361 23811 7395
rect 24026 7392 24032 7404
rect 23987 7364 24032 7392
rect 23753 7355 23811 7361
rect 24026 7352 24032 7364
rect 24084 7392 24090 7404
rect 24486 7392 24492 7404
rect 24084 7364 24492 7392
rect 24084 7352 24090 7364
rect 24486 7352 24492 7364
rect 24544 7352 24550 7404
rect 25590 7352 25596 7404
rect 25648 7392 25654 7404
rect 26050 7392 26056 7404
rect 25648 7364 26056 7392
rect 25648 7352 25654 7364
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 29365 7395 29423 7401
rect 29365 7392 29377 7395
rect 29236 7364 29377 7392
rect 29236 7352 29242 7364
rect 29365 7361 29377 7364
rect 29411 7361 29423 7395
rect 29638 7392 29644 7404
rect 29599 7364 29644 7392
rect 29365 7355 29423 7361
rect 29638 7352 29644 7364
rect 29696 7352 29702 7404
rect 31386 7392 31392 7404
rect 31347 7364 31392 7392
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 33321 7395 33379 7401
rect 33321 7361 33333 7395
rect 33367 7392 33379 7395
rect 33502 7392 33508 7404
rect 33367 7364 33508 7392
rect 33367 7361 33379 7364
rect 33321 7355 33379 7361
rect 33502 7352 33508 7364
rect 33560 7352 33566 7404
rect 33965 7395 34023 7401
rect 33965 7361 33977 7395
rect 34011 7392 34023 7395
rect 34790 7392 34796 7404
rect 34011 7364 34796 7392
rect 34011 7361 34023 7364
rect 33965 7355 34023 7361
rect 34790 7352 34796 7364
rect 34848 7352 34854 7404
rect 34992 7401 35020 7432
rect 35526 7420 35532 7432
rect 35584 7420 35590 7472
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7361 35035 7395
rect 35618 7392 35624 7404
rect 35579 7364 35624 7392
rect 34977 7355 35035 7361
rect 35618 7352 35624 7364
rect 35676 7352 35682 7404
rect 36538 7392 36544 7404
rect 36499 7364 36544 7392
rect 36538 7352 36544 7364
rect 36596 7352 36602 7404
rect 36722 7352 36728 7404
rect 36780 7392 36786 7404
rect 36817 7395 36875 7401
rect 36817 7392 36829 7395
rect 36780 7364 36829 7392
rect 36780 7352 36786 7364
rect 36817 7361 36829 7364
rect 36863 7361 36875 7395
rect 36817 7355 36875 7361
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7293 14979 7327
rect 14921 7287 14979 7293
rect 27868 7327 27926 7333
rect 27868 7293 27880 7327
rect 27914 7324 27926 7327
rect 28258 7324 28264 7336
rect 27914 7296 28264 7324
rect 27914 7293 27926 7296
rect 27868 7287 27926 7293
rect 28258 7284 28264 7296
rect 28316 7284 28322 7336
rect 30837 7327 30895 7333
rect 30837 7293 30849 7327
rect 30883 7293 30895 7327
rect 31294 7324 31300 7336
rect 31255 7296 31300 7324
rect 30837 7287 30895 7293
rect 2498 7256 2504 7268
rect 2148 7228 2504 7256
rect 2148 7200 2176 7228
rect 2498 7216 2504 7228
rect 2556 7265 2562 7268
rect 2556 7259 2604 7265
rect 2556 7225 2558 7259
rect 2592 7225 2604 7259
rect 2556 7219 2604 7225
rect 2556 7216 2562 7219
rect 5350 7216 5356 7268
rect 5408 7256 5414 7268
rect 6641 7259 6699 7265
rect 5408 7228 5453 7256
rect 5408 7216 5414 7228
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 7187 7259 7245 7265
rect 7187 7256 7199 7259
rect 6687 7228 7199 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 7187 7225 7199 7228
rect 7233 7256 7245 7259
rect 7282 7256 7288 7268
rect 7233 7228 7288 7256
rect 7233 7225 7245 7228
rect 7187 7219 7245 7225
rect 7282 7216 7288 7228
rect 7340 7256 7346 7268
rect 10505 7259 10563 7265
rect 10505 7256 10517 7259
rect 7340 7228 10517 7256
rect 7340 7216 7346 7228
rect 10505 7225 10517 7228
rect 10551 7256 10563 7259
rect 10959 7259 11017 7265
rect 10959 7256 10971 7259
rect 10551 7228 10971 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10959 7225 10971 7228
rect 11005 7256 11017 7259
rect 11005 7228 11928 7256
rect 11005 7225 11017 7228
rect 10959 7219 11017 7225
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 2130 7188 2136 7200
rect 1811 7160 2136 7188
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 8386 7188 8392 7200
rect 8347 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8478 7148 8484 7200
rect 8536 7188 8542 7200
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8536 7160 8677 7188
rect 8536 7148 8542 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 8665 7151 8723 7157
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 11900 7197 11928 7228
rect 11885 7191 11943 7197
rect 11885 7157 11897 7191
rect 11931 7188 11943 7191
rect 11974 7188 11980 7200
rect 11931 7160 11980 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 14568 7188 14596 7284
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 15286 7256 15292 7268
rect 15151 7228 15292 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 16114 7216 16120 7268
rect 16172 7256 16178 7268
rect 17862 7256 17868 7268
rect 16172 7228 16217 7256
rect 17775 7228 17868 7256
rect 16172 7216 16178 7228
rect 17862 7216 17868 7228
rect 17920 7256 17926 7268
rect 18411 7259 18469 7265
rect 18411 7256 18423 7259
rect 17920 7228 18423 7256
rect 17920 7216 17926 7228
rect 18411 7225 18423 7228
rect 18457 7256 18469 7259
rect 20302 7259 20360 7265
rect 20302 7256 20314 7259
rect 18457 7228 19196 7256
rect 18457 7225 18469 7228
rect 18411 7219 18469 7225
rect 14734 7188 14740 7200
rect 14568 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16132 7188 16160 7216
rect 19168 7200 19196 7228
rect 19812 7228 20314 7256
rect 17126 7188 17132 7200
rect 15887 7160 16160 7188
rect 17087 7160 17132 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19812 7197 19840 7228
rect 20302 7225 20314 7228
rect 20348 7256 20360 7259
rect 20622 7256 20628 7268
rect 20348 7228 20628 7256
rect 20348 7225 20360 7228
rect 20302 7219 20360 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 21913 7259 21971 7265
rect 21913 7225 21925 7259
rect 21959 7225 21971 7259
rect 22462 7256 22468 7268
rect 22423 7228 22468 7256
rect 21913 7219 21971 7225
rect 19245 7191 19303 7197
rect 19245 7188 19257 7191
rect 19208 7160 19257 7188
rect 19208 7148 19214 7160
rect 19245 7157 19257 7160
rect 19291 7188 19303 7191
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 19291 7160 19809 7188
rect 19291 7157 19303 7160
rect 19245 7151 19303 7157
rect 19797 7157 19809 7160
rect 19843 7157 19855 7191
rect 19797 7151 19855 7157
rect 21453 7191 21511 7197
rect 21453 7157 21465 7191
rect 21499 7188 21511 7191
rect 21928 7188 21956 7219
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 23845 7259 23903 7265
rect 23845 7225 23857 7259
rect 23891 7225 23903 7259
rect 24854 7256 24860 7268
rect 24815 7228 24860 7256
rect 23845 7219 23903 7225
rect 22830 7188 22836 7200
rect 21499 7160 21956 7188
rect 22791 7160 22836 7188
rect 21499 7157 21511 7160
rect 21453 7151 21511 7157
rect 22830 7148 22836 7160
rect 22888 7148 22894 7200
rect 23474 7188 23480 7200
rect 23435 7160 23480 7188
rect 23474 7148 23480 7160
rect 23532 7188 23538 7200
rect 23860 7188 23888 7219
rect 24854 7216 24860 7228
rect 24912 7216 24918 7268
rect 25958 7256 25964 7268
rect 25871 7228 25964 7256
rect 25958 7216 25964 7228
rect 26016 7256 26022 7268
rect 26415 7259 26473 7265
rect 26415 7256 26427 7259
rect 26016 7228 26427 7256
rect 26016 7216 26022 7228
rect 26415 7225 26427 7228
rect 26461 7256 26473 7259
rect 26786 7256 26792 7268
rect 26461 7228 26792 7256
rect 26461 7225 26473 7228
rect 26415 7219 26473 7225
rect 26786 7216 26792 7228
rect 26844 7256 26850 7268
rect 26844 7228 27384 7256
rect 26844 7216 26850 7228
rect 25314 7188 25320 7200
rect 23532 7160 23888 7188
rect 25275 7160 25320 7188
rect 23532 7148 23538 7160
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 27356 7197 27384 7228
rect 29454 7216 29460 7268
rect 29512 7256 29518 7268
rect 29512 7228 29557 7256
rect 29512 7216 29518 7228
rect 29822 7216 29828 7268
rect 29880 7256 29886 7268
rect 30653 7259 30711 7265
rect 30653 7256 30665 7259
rect 29880 7228 30665 7256
rect 29880 7216 29886 7228
rect 30653 7225 30665 7228
rect 30699 7256 30711 7259
rect 30852 7256 30880 7287
rect 31294 7284 31300 7296
rect 31352 7284 31358 7336
rect 30699 7228 30880 7256
rect 30699 7225 30711 7228
rect 30653 7219 30711 7225
rect 33042 7216 33048 7268
rect 33100 7256 33106 7268
rect 33413 7259 33471 7265
rect 33413 7256 33425 7259
rect 33100 7228 33425 7256
rect 33100 7216 33106 7228
rect 33413 7225 33425 7228
rect 33459 7225 33471 7259
rect 33413 7219 33471 7225
rect 35069 7259 35127 7265
rect 35069 7225 35081 7259
rect 35115 7225 35127 7259
rect 36633 7259 36691 7265
rect 36633 7256 36645 7259
rect 35069 7219 35127 7225
rect 35912 7228 36645 7256
rect 27341 7191 27399 7197
rect 27341 7157 27353 7191
rect 27387 7188 27399 7191
rect 27522 7188 27528 7200
rect 27387 7160 27528 7188
rect 27387 7157 27399 7160
rect 27341 7151 27399 7157
rect 27522 7148 27528 7160
rect 27580 7148 27586 7200
rect 29089 7191 29147 7197
rect 29089 7157 29101 7191
rect 29135 7188 29147 7191
rect 29472 7188 29500 7216
rect 29135 7160 29500 7188
rect 30377 7191 30435 7197
rect 29135 7157 29147 7160
rect 29089 7151 29147 7157
rect 30377 7157 30389 7191
rect 30423 7188 30435 7191
rect 30742 7188 30748 7200
rect 30423 7160 30748 7188
rect 30423 7157 30435 7160
rect 30377 7151 30435 7157
rect 30742 7148 30748 7160
rect 30800 7148 30806 7200
rect 32214 7188 32220 7200
rect 32175 7160 32220 7188
rect 32214 7148 32220 7160
rect 32272 7148 32278 7200
rect 34698 7188 34704 7200
rect 34659 7160 34704 7188
rect 34698 7148 34704 7160
rect 34756 7148 34762 7200
rect 34790 7148 34796 7200
rect 34848 7188 34854 7200
rect 35084 7188 35112 7219
rect 35912 7200 35940 7228
rect 36633 7225 36645 7228
rect 36679 7225 36691 7259
rect 36633 7219 36691 7225
rect 35894 7188 35900 7200
rect 34848 7160 35112 7188
rect 35855 7160 35900 7188
rect 34848 7148 34854 7160
rect 35894 7148 35900 7160
rect 35952 7148 35958 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 4249 6987 4307 6993
rect 4249 6984 4261 6987
rect 4212 6956 4261 6984
rect 4212 6944 4218 6956
rect 4249 6953 4261 6956
rect 4295 6953 4307 6987
rect 4249 6947 4307 6953
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10560 6956 10609 6984
rect 10560 6944 10566 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 10597 6947 10655 6953
rect 11974 6944 11980 6996
rect 12032 6944 12038 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 14148 6956 14473 6984
rect 14148 6944 14154 6956
rect 14461 6953 14473 6956
rect 14507 6984 14519 6987
rect 14734 6984 14740 6996
rect 14507 6956 14740 6984
rect 14507 6953 14519 6956
rect 14461 6947 14519 6953
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15749 6987 15807 6993
rect 15749 6984 15761 6987
rect 15252 6956 15761 6984
rect 15252 6944 15258 6956
rect 15749 6953 15761 6956
rect 15795 6953 15807 6987
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 15749 6947 15807 6953
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18601 6987 18659 6993
rect 18601 6953 18613 6987
rect 18647 6984 18659 6987
rect 18690 6984 18696 6996
rect 18647 6956 18696 6984
rect 18647 6953 18659 6956
rect 18601 6947 18659 6953
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 19886 6944 19892 6996
rect 19944 6984 19950 6996
rect 19981 6987 20039 6993
rect 19981 6984 19993 6987
rect 19944 6956 19993 6984
rect 19944 6944 19950 6956
rect 19981 6953 19993 6956
rect 20027 6953 20039 6987
rect 19981 6947 20039 6953
rect 20806 6944 20812 6996
rect 20864 6984 20870 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 20864 6956 21833 6984
rect 20864 6944 20870 6956
rect 21821 6953 21833 6956
rect 21867 6984 21879 6987
rect 21910 6984 21916 6996
rect 21867 6956 21916 6984
rect 21867 6953 21879 6956
rect 21821 6947 21879 6953
rect 21910 6944 21916 6956
rect 21968 6944 21974 6996
rect 22462 6944 22468 6996
rect 22520 6984 22526 6996
rect 23569 6987 23627 6993
rect 23569 6984 23581 6987
rect 22520 6956 23581 6984
rect 22520 6944 22526 6956
rect 23569 6953 23581 6956
rect 23615 6953 23627 6987
rect 26050 6984 26056 6996
rect 26011 6956 26056 6984
rect 23569 6947 23627 6953
rect 26050 6944 26056 6956
rect 26108 6944 26114 6996
rect 27709 6987 27767 6993
rect 27709 6953 27721 6987
rect 27755 6984 27767 6987
rect 28534 6984 28540 6996
rect 27755 6956 28540 6984
rect 27755 6953 27767 6956
rect 27709 6947 27767 6953
rect 28534 6944 28540 6956
rect 28592 6944 28598 6996
rect 28626 6944 28632 6996
rect 28684 6984 28690 6996
rect 28721 6987 28779 6993
rect 28721 6984 28733 6987
rect 28684 6956 28733 6984
rect 28684 6944 28690 6956
rect 28721 6953 28733 6956
rect 28767 6953 28779 6987
rect 28721 6947 28779 6953
rect 29178 6944 29184 6996
rect 29236 6984 29242 6996
rect 29273 6987 29331 6993
rect 29273 6984 29285 6987
rect 29236 6956 29285 6984
rect 29236 6944 29242 6956
rect 29273 6953 29285 6956
rect 29319 6953 29331 6987
rect 29273 6947 29331 6953
rect 29454 6944 29460 6996
rect 29512 6984 29518 6996
rect 30469 6987 30527 6993
rect 30469 6984 30481 6987
rect 29512 6956 30481 6984
rect 29512 6944 29518 6956
rect 30469 6953 30481 6956
rect 30515 6953 30527 6987
rect 30469 6947 30527 6953
rect 36538 6944 36544 6996
rect 36596 6984 36602 6996
rect 36725 6987 36783 6993
rect 36725 6984 36737 6987
rect 36596 6956 36737 6984
rect 36596 6944 36602 6956
rect 36725 6953 36737 6956
rect 36771 6953 36783 6987
rect 36725 6947 36783 6953
rect 2498 6876 2504 6928
rect 2556 6925 2562 6928
rect 2556 6919 2604 6925
rect 2556 6885 2558 6919
rect 2592 6885 2604 6919
rect 2556 6879 2604 6885
rect 2556 6876 2562 6879
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 4801 6919 4859 6925
rect 4801 6916 4813 6919
rect 4764 6888 4813 6916
rect 4764 6876 4770 6888
rect 4801 6885 4813 6888
rect 4847 6885 4859 6919
rect 4801 6879 4859 6885
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 6365 6919 6423 6925
rect 6365 6916 6377 6919
rect 6328 6888 6377 6916
rect 6328 6876 6334 6888
rect 6365 6885 6377 6888
rect 6411 6885 6423 6919
rect 6365 6879 6423 6885
rect 7929 6919 7987 6925
rect 7929 6885 7941 6919
rect 7975 6916 7987 6919
rect 8018 6916 8024 6928
rect 7975 6888 8024 6916
rect 7975 6885 7987 6888
rect 7929 6879 7987 6885
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 11419 6919 11477 6925
rect 11419 6885 11431 6919
rect 11465 6916 11477 6919
rect 11992 6916 12020 6944
rect 11465 6888 12020 6916
rect 11465 6885 11477 6888
rect 11419 6879 11477 6885
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 12989 6919 13047 6925
rect 12989 6916 13001 6919
rect 12952 6888 13001 6916
rect 12952 6876 12958 6888
rect 12989 6885 13001 6888
rect 13035 6885 13047 6919
rect 12989 6879 13047 6885
rect 16826 6919 16884 6925
rect 16826 6885 16838 6919
rect 16872 6916 16884 6919
rect 16942 6916 16948 6928
rect 16872 6888 16948 6916
rect 16872 6885 16884 6888
rect 16826 6879 16884 6885
rect 16942 6876 16948 6888
rect 17000 6916 17006 6928
rect 17862 6916 17868 6928
rect 17000 6888 17868 6916
rect 17000 6876 17006 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 18874 6916 18880 6928
rect 18835 6888 18880 6916
rect 18874 6876 18880 6888
rect 18932 6876 18938 6928
rect 20622 6876 20628 6928
rect 20680 6916 20686 6928
rect 22643 6919 22701 6925
rect 20680 6888 22140 6916
rect 20680 6876 20686 6888
rect 2038 6848 2044 6860
rect 1999 6820 2044 6848
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 2924 6820 3157 6848
rect 2924 6808 2930 6820
rect 3145 6817 3157 6820
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5408 6820 5641 6848
rect 5408 6808 5414 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9712 6851 9770 6857
rect 9712 6848 9724 6851
rect 9640 6820 9724 6848
rect 9640 6808 9646 6820
rect 9712 6817 9724 6820
rect 9758 6817 9770 6851
rect 9712 6811 9770 6817
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10836 6820 11069 6848
rect 10836 6808 10842 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11940 6820 11989 6848
rect 11940 6808 11946 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15746 6848 15752 6860
rect 15335 6820 15752 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16390 6848 16396 6860
rect 16347 6820 16396 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20128 6820 20913 6848
rect 20128 6808 20134 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6848 21143 6851
rect 21266 6848 21272 6860
rect 21131 6820 21272 6848
rect 21131 6817 21143 6820
rect 21085 6811 21143 6817
rect 21266 6808 21272 6820
rect 21324 6808 21330 6860
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6848 21511 6851
rect 22002 6848 22008 6860
rect 21499 6820 22008 6848
rect 21499 6817 21511 6820
rect 21453 6811 21511 6817
rect 22002 6808 22008 6820
rect 22060 6808 22066 6860
rect 22112 6848 22140 6888
rect 22643 6885 22655 6919
rect 22689 6885 22701 6919
rect 23474 6916 23480 6928
rect 22643 6879 22701 6885
rect 23400 6888 23480 6916
rect 22664 6848 22692 6879
rect 22922 6848 22928 6860
rect 22112 6820 22928 6848
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 23201 6851 23259 6857
rect 23201 6817 23213 6851
rect 23247 6848 23259 6851
rect 23400 6848 23428 6888
rect 23474 6876 23480 6888
rect 23532 6876 23538 6928
rect 34146 6925 34152 6928
rect 24391 6919 24449 6925
rect 24391 6885 24403 6919
rect 24437 6885 24449 6919
rect 24391 6879 24449 6885
rect 28163 6919 28221 6925
rect 28163 6885 28175 6919
rect 28209 6885 28221 6919
rect 28163 6879 28221 6885
rect 29911 6919 29969 6925
rect 29911 6885 29923 6919
rect 29957 6916 29969 6919
rect 32861 6919 32919 6925
rect 29957 6888 29991 6916
rect 29957 6885 29969 6888
rect 29911 6879 29969 6885
rect 32861 6885 32873 6919
rect 32907 6916 32919 6919
rect 34143 6916 34152 6925
rect 32907 6888 33088 6916
rect 34107 6888 34152 6916
rect 32907 6885 32919 6888
rect 32861 6879 32919 6885
rect 23247 6820 23428 6848
rect 24412 6848 24440 6879
rect 24670 6848 24676 6860
rect 24412 6820 24676 6848
rect 23247 6817 23259 6820
rect 23201 6811 23259 6817
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 24946 6848 24952 6860
rect 24907 6820 24952 6848
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 26786 6808 26792 6860
rect 26844 6857 26850 6860
rect 26844 6851 26882 6857
rect 26870 6817 26882 6851
rect 26844 6811 26882 6817
rect 26927 6851 26985 6857
rect 26927 6817 26939 6851
rect 26973 6848 26985 6851
rect 27430 6848 27436 6860
rect 26973 6820 27436 6848
rect 26973 6817 26985 6820
rect 26927 6811 26985 6817
rect 26844 6808 26850 6811
rect 27430 6808 27436 6820
rect 27488 6808 27494 6860
rect 27522 6808 27528 6860
rect 27580 6848 27586 6860
rect 28074 6848 28080 6860
rect 27580 6820 28080 6848
rect 27580 6808 27586 6820
rect 28074 6808 28080 6820
rect 28132 6848 28138 6860
rect 28184 6848 28212 6879
rect 29926 6848 29954 6879
rect 30374 6848 30380 6860
rect 28132 6820 30380 6848
rect 28132 6808 28138 6820
rect 30374 6808 30380 6820
rect 30432 6808 30438 6860
rect 30466 6808 30472 6860
rect 30524 6848 30530 6860
rect 31113 6851 31171 6857
rect 31113 6848 31125 6851
rect 30524 6820 31125 6848
rect 30524 6808 30530 6820
rect 31113 6817 31125 6820
rect 31159 6848 31171 6851
rect 31570 6848 31576 6860
rect 31159 6820 31576 6848
rect 31159 6817 31171 6820
rect 31113 6811 31171 6817
rect 31570 6808 31576 6820
rect 31628 6808 31634 6860
rect 32122 6848 32128 6860
rect 32083 6820 32128 6848
rect 32122 6808 32128 6820
rect 32180 6808 32186 6860
rect 32585 6851 32643 6857
rect 32585 6817 32597 6851
rect 32631 6848 32643 6851
rect 32766 6848 32772 6860
rect 32631 6820 32772 6848
rect 32631 6817 32643 6820
rect 32585 6811 32643 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1946 6780 1952 6792
rect 1719 6752 1952 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2590 6780 2596 6792
rect 2271 6752 2596 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 3108 6752 3433 6780
rect 3108 6740 3114 6752
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4798 6780 4804 6792
rect 4755 6752 4804 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5592 6752 6009 6780
rect 5592 6740 5598 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 6362 6780 6368 6792
rect 6319 6752 6368 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7466 6780 7472 6792
rect 6972 6752 7472 6780
rect 6972 6740 6978 6752
rect 7466 6740 7472 6752
rect 7524 6780 7530 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7524 6752 7849 6780
rect 7524 6740 7530 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5626 6712 5632 6724
rect 5307 6684 5632 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 6564 6712 6592 6740
rect 8128 6712 8156 6743
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12768 6752 12909 6780
rect 12768 6740 12774 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 13170 6780 13176 6792
rect 13131 6752 13176 6780
rect 12897 6743 12955 6749
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 16485 6783 16543 6789
rect 16485 6780 16497 6783
rect 16264 6752 16497 6780
rect 16264 6740 16270 6752
rect 16485 6749 16497 6752
rect 16531 6749 16543 6783
rect 18782 6780 18788 6792
rect 18743 6752 18788 6780
rect 16485 6743 16543 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 22281 6783 22339 6789
rect 22281 6749 22293 6783
rect 22327 6780 22339 6783
rect 22370 6780 22376 6792
rect 22327 6752 22376 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 22370 6740 22376 6752
rect 22428 6740 22434 6792
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6749 24087 6783
rect 27798 6780 27804 6792
rect 27759 6752 27804 6780
rect 24029 6743 24087 6749
rect 8202 6712 8208 6724
rect 6564 6684 8208 6712
rect 8202 6672 8208 6684
rect 8260 6712 8266 6724
rect 9125 6715 9183 6721
rect 9125 6712 9137 6715
rect 8260 6684 9137 6712
rect 8260 6672 8266 6684
rect 9125 6681 9137 6684
rect 9171 6681 9183 6715
rect 9125 6675 9183 6681
rect 18598 6672 18604 6724
rect 18656 6712 18662 6724
rect 20349 6715 20407 6721
rect 20349 6712 20361 6715
rect 18656 6684 20361 6712
rect 18656 6672 18662 6684
rect 20349 6681 20361 6684
rect 20395 6681 20407 6715
rect 20349 6675 20407 6681
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 8110 6644 8116 6656
rect 7699 6616 8116 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8846 6644 8852 6656
rect 8807 6616 8852 6644
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9766 6604 9772 6656
rect 9824 6653 9830 6656
rect 9824 6647 9873 6653
rect 9824 6613 9827 6647
rect 9861 6613 9873 6647
rect 10134 6644 10140 6656
rect 10095 6616 10140 6644
rect 9824 6607 9873 6613
rect 9824 6604 9830 6607
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 15470 6644 15476 6656
rect 15431 6616 15476 6644
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 17126 6604 17132 6656
rect 17184 6644 17190 6656
rect 17405 6647 17463 6653
rect 17405 6644 17417 6647
rect 17184 6616 17417 6644
rect 17184 6604 17190 6616
rect 17405 6613 17417 6616
rect 17451 6644 17463 6647
rect 17862 6644 17868 6656
rect 17451 6616 17868 6644
rect 17451 6613 17463 6616
rect 17405 6607 17463 6613
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 23842 6644 23848 6656
rect 23803 6616 23848 6644
rect 23842 6604 23848 6616
rect 23900 6644 23906 6656
rect 24044 6644 24072 6743
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 29546 6780 29552 6792
rect 29507 6752 29552 6780
rect 29546 6740 29552 6752
rect 29604 6740 29610 6792
rect 32600 6780 32628 6811
rect 32766 6808 32772 6820
rect 32824 6808 32830 6860
rect 33060 6848 33088 6888
rect 34143 6879 34152 6888
rect 34146 6876 34152 6879
rect 34204 6876 34210 6928
rect 34698 6876 34704 6928
rect 34756 6916 34762 6928
rect 35894 6925 35900 6928
rect 35891 6916 35900 6925
rect 34756 6888 35756 6916
rect 35855 6888 35900 6916
rect 34756 6876 34762 6888
rect 33686 6848 33692 6860
rect 33060 6820 33692 6848
rect 33686 6808 33692 6820
rect 33744 6848 33750 6860
rect 33781 6851 33839 6857
rect 33781 6848 33793 6851
rect 33744 6820 33793 6848
rect 33744 6808 33750 6820
rect 33781 6817 33793 6820
rect 33827 6817 33839 6851
rect 35342 6848 35348 6860
rect 35303 6820 35348 6848
rect 33781 6811 33839 6817
rect 35342 6808 35348 6820
rect 35400 6808 35406 6860
rect 35728 6848 35756 6888
rect 35891 6879 35900 6888
rect 35894 6876 35900 6879
rect 35952 6876 35958 6928
rect 36449 6851 36507 6857
rect 36449 6848 36461 6851
rect 35728 6820 36461 6848
rect 36449 6817 36461 6820
rect 36495 6817 36507 6851
rect 36449 6811 36507 6817
rect 31496 6752 32628 6780
rect 23900 6616 24072 6644
rect 23900 6604 23906 6616
rect 27062 6604 27068 6656
rect 27120 6644 27126 6656
rect 27249 6647 27307 6653
rect 27249 6644 27261 6647
rect 27120 6616 27261 6644
rect 27120 6604 27126 6616
rect 27249 6613 27261 6616
rect 27295 6613 27307 6647
rect 27249 6607 27307 6613
rect 30837 6647 30895 6653
rect 30837 6613 30849 6647
rect 30883 6644 30895 6647
rect 30926 6644 30932 6656
rect 30883 6616 30932 6644
rect 30883 6613 30895 6616
rect 30837 6607 30895 6613
rect 30926 6604 30932 6616
rect 30984 6644 30990 6656
rect 31294 6644 31300 6656
rect 30984 6616 31300 6644
rect 30984 6604 30990 6616
rect 31294 6604 31300 6616
rect 31352 6644 31358 6656
rect 31496 6653 31524 6752
rect 35434 6740 35440 6792
rect 35492 6780 35498 6792
rect 35529 6783 35587 6789
rect 35529 6780 35541 6783
rect 35492 6752 35541 6780
rect 35492 6740 35498 6752
rect 35529 6749 35541 6752
rect 35575 6749 35587 6783
rect 35529 6743 35587 6749
rect 34606 6672 34612 6724
rect 34664 6712 34670 6724
rect 34701 6715 34759 6721
rect 34701 6712 34713 6715
rect 34664 6684 34713 6712
rect 34664 6672 34670 6684
rect 34701 6681 34713 6684
rect 34747 6712 34759 6715
rect 35802 6712 35808 6724
rect 34747 6684 35808 6712
rect 34747 6681 34759 6684
rect 34701 6675 34759 6681
rect 35802 6672 35808 6684
rect 35860 6672 35866 6724
rect 31481 6647 31539 6653
rect 31481 6644 31493 6647
rect 31352 6616 31493 6644
rect 31352 6604 31358 6616
rect 31481 6613 31493 6616
rect 31527 6613 31539 6647
rect 33318 6644 33324 6656
rect 33279 6616 33324 6644
rect 31481 6607 31539 6613
rect 33318 6604 33324 6616
rect 33376 6604 33382 6656
rect 34790 6604 34796 6656
rect 34848 6644 34854 6656
rect 34977 6647 35035 6653
rect 34977 6644 34989 6647
rect 34848 6616 34989 6644
rect 34848 6604 34854 6616
rect 34977 6613 34989 6616
rect 35023 6613 35035 6647
rect 34977 6607 35035 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 2590 6400 2596 6452
rect 2648 6440 2654 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 2648 6412 3617 6440
rect 2648 6400 2654 6412
rect 3605 6409 3617 6412
rect 3651 6409 3663 6443
rect 3605 6403 3663 6409
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 5442 6440 5448 6452
rect 4387 6412 5448 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 3856 6239 3914 6245
rect 3856 6205 3868 6239
rect 3902 6236 3914 6239
rect 4356 6236 4384 6403
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6420 6412 6561 6440
rect 6420 6400 6426 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9125 6443 9183 6449
rect 9125 6440 9137 6443
rect 8812 6412 9137 6440
rect 8812 6400 8818 6412
rect 9125 6409 9137 6412
rect 9171 6409 9183 6443
rect 9582 6440 9588 6452
rect 9543 6412 9588 6440
rect 9125 6403 9183 6409
rect 4614 6332 4620 6384
rect 4672 6372 4678 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 4672 6344 6193 6372
rect 4672 6332 4678 6344
rect 6181 6341 6193 6344
rect 6227 6372 6239 6375
rect 6270 6372 6276 6384
rect 6227 6344 6276 6372
rect 6227 6341 6239 6344
rect 6181 6335 6239 6341
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 5258 6304 5264 6316
rect 5219 6276 5264 6304
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6546 6304 6552 6316
rect 5951 6276 6552 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 8202 6304 8208 6316
rect 8163 6276 8208 6304
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 3902 6208 4384 6236
rect 6892 6239 6950 6245
rect 3902 6205 3914 6208
rect 3856 6199 3914 6205
rect 6892 6205 6904 6239
rect 6938 6236 6950 6239
rect 7006 6236 7012 6248
rect 6938 6208 7012 6236
rect 6938 6205 6950 6208
rect 6892 6199 6950 6205
rect 7006 6196 7012 6208
rect 7064 6236 7070 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7064 6208 7297 6236
rect 7064 6196 7070 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 9140 6236 9168 6403
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 10778 6440 10784 6452
rect 10739 6412 10784 6440
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11974 6440 11980 6452
rect 11195 6412 11980 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 12802 6440 12808 6452
rect 12676 6412 12808 6440
rect 12676 6400 12682 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 12952 6412 13461 6440
rect 12952 6400 12958 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 15749 6443 15807 6449
rect 15749 6409 15761 6443
rect 15795 6440 15807 6443
rect 16206 6440 16212 6452
rect 15795 6412 16212 6440
rect 15795 6409 15807 6412
rect 15749 6403 15807 6409
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 17129 6443 17187 6449
rect 17129 6409 17141 6443
rect 17175 6440 17187 6443
rect 18509 6443 18567 6449
rect 18509 6440 18521 6443
rect 17175 6412 18521 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 18509 6409 18521 6412
rect 18555 6440 18567 6443
rect 18874 6440 18880 6452
rect 18555 6412 18880 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19668 6412 19717 6440
rect 19668 6400 19674 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 21266 6440 21272 6452
rect 21227 6412 21272 6440
rect 19705 6403 19763 6409
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 9692 6344 11529 6372
rect 9692 6245 9720 6344
rect 11517 6341 11529 6344
rect 11563 6372 11575 6375
rect 11698 6372 11704 6384
rect 11563 6344 11704 6372
rect 11563 6341 11575 6344
rect 11517 6335 11575 6341
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 13081 6375 13139 6381
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13170 6372 13176 6384
rect 13127 6344 13176 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6372 17555 6375
rect 18782 6372 18788 6384
rect 17543 6344 18788 6372
rect 17543 6341 17555 6344
rect 17497 6335 17555 6341
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 12526 6304 12532 6316
rect 12487 6276 12532 6304
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 16209 6307 16267 6313
rect 12676 6276 13952 6304
rect 12676 6264 12682 6276
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 9140 6208 9689 6236
rect 7285 6199 7343 6205
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 10134 6236 10140 6248
rect 10095 6208 10140 6236
rect 9677 6199 9735 6205
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 13924 6245 13952 6276
rect 16209 6273 16221 6307
rect 16255 6304 16267 6307
rect 16390 6304 16396 6316
rect 16255 6276 16396 6304
rect 16255 6273 16267 6276
rect 16209 6267 16267 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 19720 6304 19748 6403
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 28074 6440 28080 6452
rect 28035 6412 28080 6440
rect 28074 6400 28080 6412
rect 28132 6400 28138 6452
rect 30834 6400 30840 6452
rect 30892 6440 30898 6452
rect 30929 6443 30987 6449
rect 30929 6440 30941 6443
rect 30892 6412 30941 6440
rect 30892 6400 30898 6412
rect 30929 6409 30941 6412
rect 30975 6440 30987 6443
rect 32122 6440 32128 6452
rect 30975 6412 32128 6440
rect 30975 6409 30987 6412
rect 30929 6403 30987 6409
rect 20070 6372 20076 6384
rect 20031 6344 20076 6372
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 21818 6332 21824 6384
rect 21876 6372 21882 6384
rect 26786 6372 26792 6384
rect 21876 6344 26792 6372
rect 21876 6332 21882 6344
rect 26786 6332 26792 6344
rect 26844 6372 26850 6384
rect 27430 6372 27436 6384
rect 26844 6344 27436 6372
rect 26844 6332 26850 6344
rect 27430 6332 27436 6344
rect 27488 6332 27494 6384
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 19720 6276 20361 6304
rect 20349 6273 20361 6276
rect 20395 6273 20407 6307
rect 22370 6304 22376 6316
rect 22331 6276 22376 6304
rect 20349 6267 20407 6273
rect 22370 6264 22376 6276
rect 22428 6264 22434 6316
rect 22922 6304 22928 6316
rect 22835 6276 22928 6304
rect 22922 6264 22928 6276
rect 22980 6304 22986 6316
rect 24670 6304 24676 6316
rect 22980 6276 24676 6304
rect 22980 6264 22986 6276
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 25222 6304 25228 6316
rect 24912 6276 25228 6304
rect 24912 6264 24918 6276
rect 25222 6264 25228 6276
rect 25280 6264 25286 6316
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 27341 6307 27399 6313
rect 27341 6304 27353 6307
rect 27304 6276 27353 6304
rect 27304 6264 27310 6276
rect 27341 6273 27353 6276
rect 27387 6273 27399 6307
rect 28994 6304 29000 6316
rect 28955 6276 29000 6304
rect 27341 6267 27399 6273
rect 28994 6264 29000 6276
rect 29052 6304 29058 6316
rect 29052 6276 29316 6304
rect 29052 6264 29058 6276
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6205 11391 6239
rect 11333 6199 11391 6205
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13955 6208 14105 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 14093 6199 14151 6205
rect 21652 6208 21833 6236
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 2130 6168 2136 6180
rect 1995 6140 2136 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 2130 6128 2136 6140
rect 2188 6168 2194 6180
rect 2403 6171 2461 6177
rect 2403 6168 2415 6171
rect 2188 6140 2415 6168
rect 2188 6128 2194 6140
rect 2403 6137 2415 6140
rect 2449 6168 2461 6171
rect 3329 6171 3387 6177
rect 3329 6168 3341 6171
rect 2449 6140 3341 6168
rect 2449 6137 2461 6140
rect 2403 6131 2461 6137
rect 3329 6137 3341 6140
rect 3375 6168 3387 6171
rect 4154 6168 4160 6180
rect 3375 6140 4160 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 5350 6128 5356 6180
rect 5408 6168 5414 6180
rect 5408 6140 5453 6168
rect 5408 6128 5414 6140
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 7745 6171 7803 6177
rect 7745 6168 7757 6171
rect 6328 6140 7757 6168
rect 6328 6128 6334 6140
rect 7745 6137 7757 6140
rect 7791 6168 7803 6171
rect 8018 6168 8024 6180
rect 7791 6140 8024 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8849 6171 8907 6177
rect 8352 6140 8397 6168
rect 8352 6128 8358 6140
rect 8849 6137 8861 6171
rect 8895 6168 8907 6171
rect 10042 6168 10048 6180
rect 8895 6140 10048 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 11348 6168 11376 6199
rect 11885 6171 11943 6177
rect 11885 6168 11897 6171
rect 11348 6140 11897 6168
rect 11885 6137 11897 6140
rect 11931 6168 11943 6171
rect 12342 6168 12348 6180
rect 11931 6140 12348 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6137 12679 6171
rect 13998 6168 14004 6180
rect 13959 6140 14004 6168
rect 12621 6131 12679 6137
rect 2961 6103 3019 6109
rect 2961 6069 2973 6103
rect 3007 6100 3019 6103
rect 3142 6100 3148 6112
rect 3007 6072 3148 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 3878 6060 3884 6112
rect 3936 6109 3942 6112
rect 3936 6103 3985 6109
rect 3936 6069 3939 6103
rect 3973 6069 3985 6103
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 3936 6063 3985 6069
rect 3936 6060 3942 6063
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5368 6100 5396 6128
rect 5123 6072 5396 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 6914 6060 6920 6112
rect 6972 6109 6978 6112
rect 6972 6103 7021 6109
rect 6972 6069 6975 6103
rect 7009 6069 7021 6103
rect 6972 6063 7021 6069
rect 6972 6060 6978 6063
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9732 6072 9781 6100
rect 9732 6060 9738 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 12158 6100 12164 6112
rect 12119 6072 12164 6100
rect 9769 6063 9827 6069
rect 12158 6060 12164 6072
rect 12216 6100 12222 6112
rect 12636 6100 12664 6131
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 16117 6171 16175 6177
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 16571 6171 16629 6177
rect 16571 6168 16583 6171
rect 16163 6140 16583 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 16571 6137 16583 6140
rect 16617 6168 16629 6171
rect 16942 6168 16948 6180
rect 16617 6140 16948 6168
rect 16617 6137 16629 6140
rect 16571 6131 16629 6137
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 17862 6168 17868 6180
rect 17775 6140 17868 6168
rect 17862 6128 17868 6140
rect 17920 6168 17926 6180
rect 18782 6168 18788 6180
rect 17920 6140 18644 6168
rect 18743 6140 18788 6168
rect 17920 6128 17926 6140
rect 12216 6072 12664 6100
rect 15381 6103 15439 6109
rect 12216 6060 12222 6072
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15746 6100 15752 6112
rect 15427 6072 15752 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 18616 6100 18644 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 18877 6171 18935 6177
rect 18877 6137 18889 6171
rect 18923 6137 18935 6171
rect 19426 6168 19432 6180
rect 19339 6140 19432 6168
rect 18877 6131 18935 6137
rect 18892 6100 18920 6131
rect 19426 6128 19432 6140
rect 19484 6168 19490 6180
rect 19484 6140 20392 6168
rect 19484 6128 19490 6140
rect 18616 6072 18920 6100
rect 20364 6100 20392 6140
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 20990 6168 20996 6180
rect 20496 6140 20541 6168
rect 20951 6140 20996 6168
rect 20496 6128 20502 6140
rect 20990 6128 20996 6140
rect 21048 6128 21054 6180
rect 21008 6100 21036 6128
rect 21652 6112 21680 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 22278 6236 22284 6248
rect 21968 6208 22284 6236
rect 21968 6196 21974 6208
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23400 6208 23673 6236
rect 21634 6100 21640 6112
rect 20364 6072 21036 6100
rect 21595 6072 21640 6100
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 23106 6060 23112 6112
rect 23164 6100 23170 6112
rect 23400 6109 23428 6208
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 23661 6199 23719 6205
rect 23934 6196 23940 6248
rect 23992 6236 23998 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23992 6208 24225 6236
rect 23992 6196 23998 6208
rect 24213 6205 24225 6208
rect 24259 6236 24271 6239
rect 25314 6236 25320 6248
rect 24259 6208 25320 6236
rect 24259 6205 24271 6208
rect 24213 6199 24271 6205
rect 25314 6196 25320 6208
rect 25372 6196 25378 6248
rect 29288 6245 29316 6276
rect 29273 6239 29331 6245
rect 29273 6205 29285 6239
rect 29319 6205 29331 6239
rect 29730 6236 29736 6248
rect 29691 6208 29736 6236
rect 29273 6199 29331 6205
rect 29730 6196 29736 6208
rect 29788 6196 29794 6248
rect 30944 6236 30972 6403
rect 32122 6400 32128 6412
rect 32180 6400 32186 6452
rect 32214 6400 32220 6452
rect 32272 6440 32278 6452
rect 34146 6440 34152 6452
rect 32272 6412 34152 6440
rect 32272 6400 32278 6412
rect 34146 6400 34152 6412
rect 34204 6440 34210 6452
rect 34241 6443 34299 6449
rect 34241 6440 34253 6443
rect 34204 6412 34253 6440
rect 34204 6400 34210 6412
rect 34241 6409 34253 6412
rect 34287 6440 34299 6443
rect 35894 6440 35900 6452
rect 34287 6412 35900 6440
rect 34287 6409 34299 6412
rect 34241 6403 34299 6409
rect 35894 6400 35900 6412
rect 35952 6400 35958 6452
rect 34977 6307 35035 6313
rect 34977 6273 34989 6307
rect 35023 6304 35035 6307
rect 35342 6304 35348 6316
rect 35023 6276 35348 6304
rect 35023 6273 35035 6276
rect 34977 6267 35035 6273
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 35618 6264 35624 6316
rect 35676 6304 35682 6316
rect 36817 6307 36875 6313
rect 36817 6304 36829 6307
rect 35676 6276 36829 6304
rect 35676 6264 35682 6276
rect 36817 6273 36829 6276
rect 36863 6273 36875 6307
rect 36817 6267 36875 6273
rect 31113 6239 31171 6245
rect 31113 6236 31125 6239
rect 30944 6208 31125 6236
rect 31113 6205 31125 6208
rect 31159 6205 31171 6239
rect 31570 6236 31576 6248
rect 31531 6208 31576 6236
rect 31113 6199 31171 6205
rect 31570 6196 31576 6208
rect 31628 6196 31634 6248
rect 33965 6239 34023 6245
rect 33965 6205 33977 6239
rect 34011 6236 34023 6239
rect 34422 6236 34428 6248
rect 34011 6208 34428 6236
rect 34011 6205 34023 6208
rect 33965 6199 34023 6205
rect 34422 6196 34428 6208
rect 34480 6196 34486 6248
rect 35802 6196 35808 6248
rect 35860 6236 35866 6248
rect 36265 6239 36323 6245
rect 36265 6236 36277 6239
rect 35860 6208 36277 6236
rect 35860 6196 35866 6208
rect 36265 6205 36277 6208
rect 36311 6205 36323 6239
rect 36265 6199 36323 6205
rect 24394 6168 24400 6180
rect 24355 6140 24400 6168
rect 24394 6128 24400 6140
rect 24452 6128 24458 6180
rect 24670 6128 24676 6180
rect 24728 6168 24734 6180
rect 24765 6171 24823 6177
rect 24765 6168 24777 6171
rect 24728 6140 24777 6168
rect 24728 6128 24734 6140
rect 24765 6137 24777 6140
rect 24811 6168 24823 6171
rect 24854 6168 24860 6180
rect 24811 6140 24860 6168
rect 24811 6137 24823 6140
rect 24765 6131 24823 6137
rect 24854 6128 24860 6140
rect 24912 6168 24918 6180
rect 25133 6171 25191 6177
rect 25133 6168 25145 6171
rect 24912 6140 25145 6168
rect 24912 6128 24918 6140
rect 25133 6137 25145 6140
rect 25179 6168 25191 6171
rect 25587 6171 25645 6177
rect 25587 6168 25599 6171
rect 25179 6140 25599 6168
rect 25179 6137 25191 6140
rect 25133 6131 25191 6137
rect 25587 6137 25599 6140
rect 25633 6168 25645 6171
rect 25958 6168 25964 6180
rect 25633 6140 25964 6168
rect 25633 6137 25645 6140
rect 25587 6131 25645 6137
rect 25958 6128 25964 6140
rect 26016 6128 26022 6180
rect 26513 6171 26571 6177
rect 26513 6137 26525 6171
rect 26559 6168 26571 6171
rect 27062 6168 27068 6180
rect 26559 6140 26924 6168
rect 27023 6140 27068 6168
rect 26559 6137 26571 6140
rect 26513 6131 26571 6137
rect 26896 6112 26924 6140
rect 27062 6128 27068 6140
rect 27120 6128 27126 6180
rect 27157 6171 27215 6177
rect 27157 6137 27169 6171
rect 27203 6137 27215 6171
rect 27157 6131 27215 6137
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 23164 6072 23397 6100
rect 23164 6060 23170 6072
rect 23385 6069 23397 6072
rect 23431 6069 23443 6103
rect 23385 6063 23443 6069
rect 26050 6060 26056 6112
rect 26108 6100 26114 6112
rect 26145 6103 26203 6109
rect 26145 6100 26157 6103
rect 26108 6072 26157 6100
rect 26108 6060 26114 6072
rect 26145 6069 26157 6072
rect 26191 6069 26203 6103
rect 26145 6063 26203 6069
rect 26878 6060 26884 6112
rect 26936 6100 26942 6112
rect 27172 6100 27200 6131
rect 27798 6128 27804 6180
rect 27856 6168 27862 6180
rect 28445 6171 28503 6177
rect 28445 6168 28457 6171
rect 27856 6140 28457 6168
rect 27856 6128 27862 6140
rect 28445 6137 28457 6140
rect 28491 6168 28503 6171
rect 31846 6168 31852 6180
rect 28491 6140 29408 6168
rect 31807 6140 31852 6168
rect 28491 6137 28503 6140
rect 28445 6131 28503 6137
rect 29380 6109 29408 6140
rect 31846 6128 31852 6140
rect 31904 6128 31910 6180
rect 33318 6168 33324 6180
rect 33279 6140 33324 6168
rect 33318 6128 33324 6140
rect 33376 6128 33382 6180
rect 33413 6171 33471 6177
rect 33413 6137 33425 6171
rect 33459 6137 33471 6171
rect 34609 6171 34667 6177
rect 34609 6168 34621 6171
rect 33413 6131 33471 6137
rect 34072 6140 34621 6168
rect 26936 6072 27200 6100
rect 29365 6103 29423 6109
rect 26936 6060 26942 6072
rect 29365 6069 29377 6103
rect 29411 6069 29423 6103
rect 29365 6063 29423 6069
rect 30377 6103 30435 6109
rect 30377 6069 30389 6103
rect 30423 6100 30435 6103
rect 30466 6100 30472 6112
rect 30423 6072 30472 6100
rect 30423 6069 30435 6072
rect 30377 6063 30435 6069
rect 30466 6060 30472 6072
rect 30524 6060 30530 6112
rect 30926 6060 30932 6112
rect 30984 6100 30990 6112
rect 32493 6103 32551 6109
rect 32493 6100 32505 6103
rect 30984 6072 32505 6100
rect 30984 6060 30990 6072
rect 32493 6069 32505 6072
rect 32539 6069 32551 6103
rect 33134 6100 33140 6112
rect 33095 6072 33140 6100
rect 32493 6063 32551 6069
rect 33134 6060 33140 6072
rect 33192 6100 33198 6112
rect 33428 6100 33456 6131
rect 34072 6100 34100 6140
rect 34609 6137 34621 6140
rect 34655 6137 34667 6171
rect 34609 6131 34667 6137
rect 35069 6171 35127 6177
rect 35069 6137 35081 6171
rect 35115 6137 35127 6171
rect 35069 6131 35127 6137
rect 35621 6171 35679 6177
rect 35621 6137 35633 6171
rect 35667 6168 35679 6171
rect 35986 6168 35992 6180
rect 35667 6140 35992 6168
rect 35667 6137 35679 6140
rect 35621 6131 35679 6137
rect 33192 6072 34100 6100
rect 34624 6100 34652 6131
rect 35084 6100 35112 6131
rect 35986 6128 35992 6140
rect 36044 6128 36050 6180
rect 34624 6072 35112 6100
rect 36280 6100 36308 6199
rect 36538 6168 36544 6180
rect 36499 6140 36544 6168
rect 36538 6128 36544 6140
rect 36596 6128 36602 6180
rect 36633 6171 36691 6177
rect 36633 6137 36645 6171
rect 36679 6137 36691 6171
rect 36633 6131 36691 6137
rect 36648 6100 36676 6131
rect 36280 6072 36676 6100
rect 33192 6060 33198 6072
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 4614 5896 4620 5908
rect 2915 5868 4620 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5896 5043 5899
rect 5350 5896 5356 5908
rect 5031 5868 5356 5896
rect 5031 5865 5043 5868
rect 4985 5859 5043 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 7466 5896 7472 5908
rect 5736 5868 7328 5896
rect 7427 5868 7472 5896
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5828 1823 5831
rect 2130 5828 2136 5840
rect 1811 5800 2136 5828
rect 1811 5797 1823 5800
rect 1765 5791 1823 5797
rect 2130 5788 2136 5800
rect 2188 5828 2194 5840
rect 2270 5831 2328 5837
rect 2270 5828 2282 5831
rect 2188 5800 2282 5828
rect 2188 5788 2194 5800
rect 2270 5797 2282 5800
rect 2316 5797 2328 5831
rect 2270 5791 2328 5797
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4427 5831 4485 5837
rect 4427 5828 4439 5831
rect 4212 5800 4439 5828
rect 4212 5788 4218 5800
rect 4427 5797 4439 5800
rect 4473 5828 4485 5831
rect 4473 5800 5120 5828
rect 4473 5797 4485 5800
rect 4427 5791 4485 5797
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 1949 5763 2007 5769
rect 1949 5760 1961 5763
rect 1912 5732 1961 5760
rect 1912 5720 1918 5732
rect 1949 5729 1961 5732
rect 1995 5729 2007 5763
rect 3234 5760 3240 5772
rect 3195 5732 3240 5760
rect 1949 5723 2007 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 4028 5732 4077 5760
rect 4028 5720 4034 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 5092 5760 5120 5800
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5629 5831 5687 5837
rect 5629 5828 5641 5831
rect 5316 5800 5641 5828
rect 5316 5788 5322 5800
rect 5629 5797 5641 5800
rect 5675 5797 5687 5831
rect 5629 5791 5687 5797
rect 5736 5760 5764 5868
rect 7300 5840 7328 5868
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8352 5868 8861 5896
rect 8352 5856 8358 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 12437 5899 12495 5905
rect 12437 5865 12449 5899
rect 12483 5896 12495 5899
rect 12618 5896 12624 5908
rect 12483 5868 12624 5896
rect 12483 5865 12495 5868
rect 12437 5859 12495 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 12710 5856 12716 5908
rect 12768 5896 12774 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12768 5868 12817 5896
rect 12768 5856 12774 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 14642 5896 14648 5908
rect 14603 5868 14648 5896
rect 12805 5859 12863 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15562 5896 15568 5908
rect 15523 5868 15568 5896
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 22370 5896 22376 5908
rect 22331 5868 22376 5896
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 23753 5899 23811 5905
rect 23753 5865 23765 5899
rect 23799 5896 23811 5899
rect 23934 5896 23940 5908
rect 23799 5868 23940 5896
rect 23799 5865 23811 5868
rect 23753 5859 23811 5865
rect 23934 5856 23940 5868
rect 23992 5856 23998 5908
rect 25222 5896 25228 5908
rect 25183 5868 25228 5896
rect 25222 5856 25228 5868
rect 25280 5856 25286 5908
rect 29546 5856 29552 5908
rect 29604 5896 29610 5908
rect 29641 5899 29699 5905
rect 29641 5896 29653 5899
rect 29604 5868 29653 5896
rect 29604 5856 29610 5868
rect 29641 5865 29653 5868
rect 29687 5865 29699 5899
rect 31202 5896 31208 5908
rect 31163 5868 31208 5896
rect 29641 5859 29699 5865
rect 31202 5856 31208 5868
rect 31260 5856 31266 5908
rect 33042 5896 33048 5908
rect 33003 5868 33048 5896
rect 33042 5856 33048 5868
rect 33100 5856 33106 5908
rect 33686 5896 33692 5908
rect 33647 5868 33692 5896
rect 33686 5856 33692 5868
rect 33744 5856 33750 5908
rect 34790 5896 34796 5908
rect 34751 5868 34796 5896
rect 34790 5856 34796 5868
rect 34848 5856 34854 5908
rect 35066 5896 35072 5908
rect 35027 5868 35072 5896
rect 35066 5856 35072 5868
rect 35124 5856 35130 5908
rect 36538 5856 36544 5908
rect 36596 5896 36602 5908
rect 36633 5899 36691 5905
rect 36633 5896 36645 5899
rect 36596 5868 36645 5896
rect 36596 5856 36602 5868
rect 36633 5865 36645 5868
rect 36679 5865 36691 5899
rect 36633 5859 36691 5865
rect 6270 5828 6276 5840
rect 6231 5800 6276 5828
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 8015 5831 8073 5837
rect 8015 5828 8027 5831
rect 7340 5800 8027 5828
rect 7340 5788 7346 5800
rect 8015 5797 8027 5800
rect 8061 5828 8073 5831
rect 8110 5828 8116 5840
rect 8061 5800 8116 5828
rect 8061 5797 8073 5800
rect 8015 5791 8073 5797
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 8588 5800 9873 5828
rect 5092 5732 5764 5760
rect 4065 5723 4123 5729
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7248 5732 7665 5760
rect 7248 5720 7254 5732
rect 7653 5729 7665 5732
rect 7699 5760 7711 5763
rect 8478 5760 8484 5772
rect 7699 5732 8484 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 8588 5769 8616 5800
rect 9861 5797 9873 5800
rect 9907 5828 9919 5831
rect 10410 5828 10416 5840
rect 9907 5800 10416 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 11879 5831 11937 5837
rect 11879 5797 11891 5831
rect 11925 5828 11937 5831
rect 11974 5828 11980 5840
rect 11925 5800 11980 5828
rect 11925 5797 11937 5800
rect 11879 5791 11937 5797
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 13449 5831 13507 5837
rect 13449 5797 13461 5831
rect 13495 5828 13507 5831
rect 13998 5828 14004 5840
rect 13495 5800 14004 5828
rect 13495 5797 13507 5800
rect 13449 5791 13507 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 16301 5831 16359 5837
rect 16301 5797 16313 5831
rect 16347 5828 16359 5831
rect 16390 5828 16396 5840
rect 16347 5800 16396 5828
rect 16347 5797 16359 5800
rect 16301 5791 16359 5797
rect 16390 5788 16396 5800
rect 16448 5828 16454 5840
rect 16755 5831 16813 5837
rect 16755 5828 16767 5831
rect 16448 5800 16767 5828
rect 16448 5788 16454 5800
rect 16755 5797 16767 5800
rect 16801 5828 16813 5831
rect 16942 5828 16948 5840
rect 16801 5800 16948 5828
rect 16801 5797 16813 5800
rect 16755 5791 16813 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 18785 5831 18843 5837
rect 18785 5828 18797 5831
rect 18432 5800 18797 5828
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 14826 5720 14832 5772
rect 14884 5760 14890 5772
rect 15194 5760 15200 5772
rect 14884 5732 15200 5760
rect 14884 5720 14890 5732
rect 15194 5720 15200 5732
rect 15252 5760 15258 5772
rect 18432 5769 18460 5800
rect 18785 5797 18797 5800
rect 18831 5828 18843 5831
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 18831 5800 20269 5828
rect 18831 5797 18843 5800
rect 18785 5791 18843 5797
rect 20257 5797 20269 5800
rect 20303 5828 20315 5831
rect 20438 5828 20444 5840
rect 20303 5800 20444 5828
rect 20303 5797 20315 5800
rect 20257 5791 20315 5797
rect 20438 5788 20444 5800
rect 20496 5788 20502 5840
rect 20806 5788 20812 5840
rect 20864 5828 20870 5840
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 20864 5800 21097 5828
rect 20864 5788 20870 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21085 5791 21143 5797
rect 21637 5831 21695 5837
rect 21637 5797 21649 5831
rect 21683 5828 21695 5831
rect 21726 5828 21732 5840
rect 21683 5800 21732 5828
rect 21683 5797 21695 5800
rect 21637 5791 21695 5797
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 22278 5788 22284 5840
rect 22336 5828 22342 5840
rect 23201 5831 23259 5837
rect 22336 5800 22968 5828
rect 22336 5788 22342 5800
rect 22940 5769 22968 5800
rect 23201 5797 23213 5831
rect 23247 5828 23259 5831
rect 23842 5828 23848 5840
rect 23247 5800 23848 5828
rect 23247 5797 23259 5800
rect 23201 5791 23259 5797
rect 23842 5788 23848 5800
rect 23900 5788 23906 5840
rect 24391 5831 24449 5837
rect 24391 5797 24403 5831
rect 24437 5828 24449 5831
rect 24854 5828 24860 5840
rect 24437 5800 24860 5828
rect 24437 5797 24449 5800
rect 24391 5791 24449 5797
rect 24854 5788 24860 5800
rect 24912 5788 24918 5840
rect 26326 5788 26332 5840
rect 26384 5828 26390 5840
rect 26697 5831 26755 5837
rect 26697 5828 26709 5831
rect 26384 5800 26709 5828
rect 26384 5788 26390 5800
rect 26697 5797 26709 5800
rect 26743 5797 26755 5831
rect 28258 5828 28264 5840
rect 28219 5800 28264 5828
rect 26697 5791 26755 5797
rect 28258 5788 28264 5800
rect 28316 5788 28322 5840
rect 30466 5788 30472 5840
rect 30524 5828 30530 5840
rect 30606 5831 30664 5837
rect 30606 5828 30618 5831
rect 30524 5800 30618 5828
rect 30524 5788 30530 5800
rect 30606 5797 30618 5800
rect 30652 5797 30664 5831
rect 30606 5791 30664 5797
rect 32214 5788 32220 5840
rect 32272 5828 32278 5840
rect 32446 5831 32504 5837
rect 32446 5828 32458 5831
rect 32272 5800 32458 5828
rect 32272 5788 32278 5800
rect 32446 5797 32458 5800
rect 32492 5797 32504 5831
rect 32446 5791 32504 5797
rect 34146 5788 34152 5840
rect 34204 5837 34210 5840
rect 34204 5831 34252 5837
rect 34204 5797 34206 5831
rect 34240 5797 34252 5831
rect 35434 5828 35440 5840
rect 35395 5800 35440 5828
rect 34204 5791 34252 5797
rect 34204 5788 34210 5791
rect 35434 5788 35440 5800
rect 35492 5788 35498 5840
rect 35802 5828 35808 5840
rect 35763 5800 35808 5828
rect 35802 5788 35808 5800
rect 35860 5788 35866 5840
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 15252 5732 15393 5760
rect 15252 5720 15258 5732
rect 15381 5729 15393 5732
rect 15427 5729 15439 5763
rect 15381 5723 15439 5729
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5760 17371 5763
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 17359 5732 18429 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5729 22799 5763
rect 22741 5723 22799 5729
rect 22925 5763 22983 5769
rect 22925 5729 22937 5763
rect 22971 5729 22983 5763
rect 22925 5723 22983 5729
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 4856 5664 5273 5692
rect 4856 5652 4862 5664
rect 5261 5661 5273 5664
rect 5307 5661 5319 5695
rect 6178 5692 6184 5704
rect 6139 5664 6184 5692
rect 5261 5655 5319 5661
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 6503 5664 9413 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 9401 5661 9413 5664
rect 9447 5692 9459 5695
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9447 5664 9781 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 9769 5655 9827 5661
rect 5626 5584 5632 5636
rect 5684 5624 5690 5636
rect 6472 5624 6500 5655
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 5684 5596 6500 5624
rect 5684 5584 5690 5596
rect 566 5516 572 5568
rect 624 5556 630 5568
rect 8386 5556 8392 5568
rect 624 5528 8392 5556
rect 624 5516 630 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 10502 5516 10508 5568
rect 10560 5556 10566 5568
rect 10965 5559 11023 5565
rect 10965 5556 10977 5559
rect 10560 5528 10977 5556
rect 10560 5516 10566 5528
rect 10965 5525 10977 5528
rect 11011 5525 11023 5559
rect 11422 5556 11428 5568
rect 11383 5528 11428 5556
rect 10965 5519 11023 5525
rect 11422 5516 11428 5528
rect 11480 5556 11486 5568
rect 11532 5556 11560 5655
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12124 5664 13369 5692
rect 12124 5652 12130 5664
rect 13357 5661 13369 5664
rect 13403 5692 13415 5695
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 13403 5664 15025 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 15344 5664 16405 5692
rect 15344 5652 15350 5664
rect 16393 5661 16405 5664
rect 16439 5692 16451 5695
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 16439 5664 17969 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 17957 5661 17969 5664
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5661 18751 5695
rect 18966 5692 18972 5704
rect 18927 5664 18972 5692
rect 18693 5655 18751 5661
rect 12526 5584 12532 5636
rect 12584 5624 12590 5636
rect 13446 5624 13452 5636
rect 12584 5596 13452 5624
rect 12584 5584 12590 5596
rect 13446 5584 13452 5596
rect 13504 5624 13510 5636
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 13504 5596 13921 5624
rect 13504 5584 13510 5596
rect 13909 5593 13921 5596
rect 13955 5593 13967 5627
rect 18708 5624 18736 5655
rect 18966 5652 18972 5664
rect 19024 5692 19030 5704
rect 20714 5692 20720 5704
rect 19024 5664 20720 5692
rect 19024 5652 19030 5664
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 20990 5692 20996 5704
rect 20903 5664 20996 5692
rect 20990 5652 20996 5664
rect 21048 5692 21054 5704
rect 21910 5692 21916 5704
rect 21048 5664 21916 5692
rect 21048 5652 21054 5664
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22756 5692 22784 5723
rect 33134 5720 33140 5772
rect 33192 5760 33198 5772
rect 33873 5763 33931 5769
rect 33873 5760 33885 5763
rect 33192 5732 33885 5760
rect 33192 5720 33198 5732
rect 33873 5729 33885 5732
rect 33919 5760 33931 5763
rect 34054 5760 34060 5772
rect 33919 5732 34060 5760
rect 33919 5729 33931 5732
rect 33873 5723 33931 5729
rect 34054 5720 34060 5732
rect 34112 5720 34118 5772
rect 23106 5692 23112 5704
rect 22756 5664 23112 5692
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 24026 5692 24032 5704
rect 23987 5664 24032 5692
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 26605 5695 26663 5701
rect 26605 5692 26617 5695
rect 26292 5664 26617 5692
rect 26292 5652 26298 5664
rect 26605 5661 26617 5664
rect 26651 5661 26663 5695
rect 27246 5692 27252 5704
rect 27207 5664 27252 5692
rect 26605 5655 26663 5661
rect 27246 5652 27252 5664
rect 27304 5652 27310 5704
rect 28166 5692 28172 5704
rect 28127 5664 28172 5692
rect 28166 5652 28172 5664
rect 28224 5692 28230 5704
rect 28350 5692 28356 5704
rect 28224 5664 28356 5692
rect 28224 5652 28230 5664
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 29270 5692 29276 5704
rect 29231 5664 29276 5692
rect 28445 5655 28503 5661
rect 19058 5624 19064 5636
rect 18708 5596 19064 5624
rect 13909 5587 13967 5593
rect 19058 5584 19064 5596
rect 19116 5584 19122 5636
rect 20732 5624 20760 5652
rect 22005 5627 22063 5633
rect 22005 5624 22017 5627
rect 20732 5596 22017 5624
rect 22005 5593 22017 5596
rect 22051 5593 22063 5627
rect 22005 5587 22063 5593
rect 24949 5627 25007 5633
rect 24949 5593 24961 5627
rect 24995 5624 25007 5627
rect 26326 5624 26332 5636
rect 24995 5596 26332 5624
rect 24995 5593 25007 5596
rect 24949 5587 25007 5593
rect 26326 5584 26332 5596
rect 26384 5584 26390 5636
rect 28460 5624 28488 5655
rect 29270 5652 29276 5664
rect 29328 5692 29334 5704
rect 29730 5692 29736 5704
rect 29328 5664 29736 5692
rect 29328 5652 29334 5664
rect 29730 5652 29736 5664
rect 29788 5652 29794 5704
rect 30282 5692 30288 5704
rect 30243 5664 30288 5692
rect 30282 5652 30288 5664
rect 30340 5652 30346 5704
rect 31938 5652 31944 5704
rect 31996 5692 32002 5704
rect 32125 5695 32183 5701
rect 32125 5692 32137 5695
rect 31996 5664 32137 5692
rect 31996 5652 32002 5664
rect 32125 5661 32137 5664
rect 32171 5692 32183 5695
rect 33042 5692 33048 5704
rect 32171 5664 33048 5692
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 33042 5652 33048 5664
rect 33100 5652 33106 5704
rect 35066 5652 35072 5704
rect 35124 5692 35130 5704
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 35124 5664 35725 5692
rect 35124 5652 35130 5664
rect 35713 5661 35725 5664
rect 35759 5661 35771 5695
rect 35986 5692 35992 5704
rect 35947 5664 35992 5692
rect 35713 5655 35771 5661
rect 35986 5652 35992 5664
rect 36044 5652 36050 5704
rect 28184 5596 28488 5624
rect 28184 5568 28212 5596
rect 11480 5528 11560 5556
rect 11480 5516 11486 5528
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 13872 5528 14289 5556
rect 13872 5516 13878 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 15838 5556 15844 5568
rect 15799 5528 15844 5556
rect 14277 5519 14335 5525
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 16850 5516 16856 5568
rect 16908 5556 16914 5568
rect 17589 5559 17647 5565
rect 17589 5556 17601 5559
rect 16908 5528 17601 5556
rect 16908 5516 16914 5528
rect 17589 5525 17601 5528
rect 17635 5525 17647 5559
rect 19702 5556 19708 5568
rect 19663 5528 19708 5556
rect 17589 5519 17647 5525
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 20622 5516 20628 5568
rect 20680 5556 20686 5568
rect 20717 5559 20775 5565
rect 20717 5556 20729 5559
rect 20680 5528 20729 5556
rect 20680 5516 20686 5528
rect 20717 5525 20729 5528
rect 20763 5525 20775 5559
rect 20717 5519 20775 5525
rect 28166 5516 28172 5568
rect 28224 5516 28230 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5352 2099 5355
rect 2682 5352 2688 5364
rect 2087 5324 2688 5352
rect 2087 5321 2099 5324
rect 2041 5315 2099 5321
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2056 5148 2084 5315
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5534 5352 5540 5364
rect 5495 5324 5540 5352
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6270 5352 6276 5364
rect 6227 5324 6276 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 7190 5352 7196 5364
rect 7151 5324 7196 5352
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8352 5324 8585 5352
rect 8352 5312 8358 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9582 5352 9588 5364
rect 8987 5324 9588 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 2406 5244 2412 5296
rect 2464 5284 2470 5296
rect 2593 5287 2651 5293
rect 2593 5284 2605 5287
rect 2464 5256 2605 5284
rect 2464 5244 2470 5256
rect 2593 5253 2605 5256
rect 2639 5284 2651 5287
rect 4172 5284 4200 5312
rect 2639 5256 4200 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 3050 5216 3056 5228
rect 2731 5188 3056 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 1443 5120 2084 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 3047 5083 3105 5089
rect 3047 5049 3059 5083
rect 3093 5080 3105 5083
rect 3160 5080 3188 5256
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 3936 5188 4537 5216
rect 3936 5176 3942 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4764 5188 4813 5216
rect 4764 5176 4770 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6236 5188 6469 5216
rect 6236 5176 6242 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 8956 5216 8984 5315
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10410 5352 10416 5364
rect 10371 5324 10416 5352
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 12986 5352 12992 5364
rect 12947 5324 12992 5352
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 15194 5352 15200 5364
rect 15155 5324 15200 5352
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 16390 5352 16396 5364
rect 16351 5324 16396 5352
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17034 5352 17040 5364
rect 16995 5324 17040 5352
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 22373 5355 22431 5361
rect 22373 5352 22385 5355
rect 22336 5324 22385 5352
rect 22336 5312 22342 5324
rect 22373 5321 22385 5324
rect 22419 5321 22431 5355
rect 24854 5352 24860 5364
rect 24815 5324 24860 5352
rect 22373 5315 22431 5321
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 26326 5352 26332 5364
rect 26287 5324 26332 5352
rect 26326 5312 26332 5324
rect 26384 5352 26390 5364
rect 28077 5355 28135 5361
rect 28077 5352 28089 5355
rect 26384 5324 28089 5352
rect 26384 5312 26390 5324
rect 28077 5321 28089 5324
rect 28123 5352 28135 5355
rect 28258 5352 28264 5364
rect 28123 5324 28264 5352
rect 28123 5321 28135 5324
rect 28077 5315 28135 5321
rect 28258 5312 28264 5324
rect 28316 5312 28322 5364
rect 28350 5312 28356 5364
rect 28408 5352 28414 5364
rect 28445 5355 28503 5361
rect 28445 5352 28457 5355
rect 28408 5324 28457 5352
rect 28408 5312 28414 5324
rect 28445 5321 28457 5324
rect 28491 5321 28503 5355
rect 28445 5315 28503 5321
rect 33134 5312 33140 5364
rect 33192 5352 33198 5364
rect 33505 5355 33563 5361
rect 33505 5352 33517 5355
rect 33192 5324 33517 5352
rect 33192 5312 33198 5324
rect 33505 5321 33517 5324
rect 33551 5321 33563 5355
rect 33505 5315 33563 5321
rect 34054 5312 34060 5364
rect 34112 5352 34118 5364
rect 34241 5355 34299 5361
rect 34241 5352 34253 5355
rect 34112 5324 34253 5352
rect 34112 5312 34118 5324
rect 34241 5321 34253 5324
rect 34287 5321 34299 5355
rect 34241 5315 34299 5321
rect 34606 5312 34612 5364
rect 34664 5352 34670 5364
rect 34974 5352 34980 5364
rect 34664 5324 34980 5352
rect 34664 5312 34670 5324
rect 34974 5312 34980 5324
rect 35032 5352 35038 5364
rect 35618 5352 35624 5364
rect 35032 5324 35624 5352
rect 35032 5312 35038 5324
rect 35618 5312 35624 5324
rect 35676 5312 35682 5364
rect 35894 5352 35900 5364
rect 35855 5324 35900 5352
rect 35894 5312 35900 5324
rect 35952 5312 35958 5364
rect 12621 5287 12679 5293
rect 12621 5253 12633 5287
rect 12667 5284 12679 5287
rect 12710 5284 12716 5296
rect 12667 5256 12716 5284
rect 12667 5253 12679 5256
rect 12621 5247 12679 5253
rect 12710 5244 12716 5256
rect 12768 5284 12774 5296
rect 13078 5284 13084 5296
rect 12768 5256 13084 5284
rect 12768 5244 12774 5256
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 13449 5287 13507 5293
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 16408 5284 16436 5312
rect 18230 5284 18236 5296
rect 13495 5256 16436 5284
rect 18191 5256 18236 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 7699 5188 8984 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 12032 5188 12265 5216
rect 12032 5176 12038 5188
rect 12253 5185 12265 5188
rect 12299 5216 12311 5219
rect 13464 5216 13492 5247
rect 12299 5188 13492 5216
rect 13541 5219 13599 5225
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 13722 5216 13728 5228
rect 13587 5188 13728 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 6822 5108 6828 5160
rect 6880 5148 6886 5160
rect 9582 5148 9588 5160
rect 6880 5120 9352 5148
rect 9543 5120 9588 5148
rect 6880 5108 6886 5120
rect 4617 5083 4675 5089
rect 4617 5080 4629 5083
rect 3093 5052 3188 5080
rect 3620 5052 4629 5080
rect 3093 5049 3105 5052
rect 3047 5043 3105 5049
rect 3620 5024 3648 5052
rect 4617 5049 4629 5052
rect 4663 5049 4675 5083
rect 4617 5043 4675 5049
rect 7561 5083 7619 5089
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 8015 5083 8073 5089
rect 8015 5080 8027 5083
rect 7607 5052 8027 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 8015 5049 8027 5052
rect 8061 5080 8073 5083
rect 8110 5080 8116 5092
rect 8061 5052 8116 5080
rect 8061 5049 8073 5052
rect 8015 5043 8073 5049
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 9324 5089 9352 5120
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9950 5148 9956 5160
rect 9911 5120 9956 5148
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 11146 5148 11152 5160
rect 10919 5120 11152 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12526 5148 12532 5160
rect 12483 5120 12532 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12526 5108 12532 5120
rect 12584 5148 12590 5160
rect 12986 5148 12992 5160
rect 12584 5120 12992 5148
rect 12584 5108 12590 5120
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 9309 5083 9367 5089
rect 9309 5049 9321 5083
rect 9355 5080 9367 5083
rect 9968 5080 9996 5108
rect 9355 5052 9996 5080
rect 10965 5083 11023 5089
rect 9355 5049 9367 5052
rect 9309 5043 9367 5049
rect 10965 5049 10977 5083
rect 11011 5049 11023 5083
rect 11514 5080 11520 5092
rect 11475 5052 11520 5080
rect 10965 5043 11023 5049
rect 3602 5012 3608 5024
rect 3563 4984 3608 5012
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 9674 5012 9680 5024
rect 9635 4984 9680 5012
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10980 5012 11008 5043
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 13918 5089 13946 5256
rect 18230 5244 18236 5256
rect 18288 5244 18294 5296
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 22152 5256 22197 5284
rect 22152 5244 22158 5256
rect 26050 5244 26056 5296
rect 26108 5284 26114 5296
rect 26605 5287 26663 5293
rect 26605 5284 26617 5287
rect 26108 5256 26617 5284
rect 26108 5244 26114 5256
rect 26605 5253 26617 5256
rect 26651 5284 26663 5287
rect 26697 5287 26755 5293
rect 26697 5284 26709 5287
rect 26651 5256 26709 5284
rect 26651 5253 26663 5256
rect 26605 5247 26663 5253
rect 26697 5253 26709 5256
rect 26743 5253 26755 5287
rect 32125 5287 32183 5293
rect 32125 5284 32137 5287
rect 26697 5247 26755 5253
rect 31772 5256 32137 5284
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15378 5216 15384 5228
rect 14875 5188 15384 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 20714 5176 20720 5228
rect 20772 5216 20778 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20772 5188 21097 5216
rect 20772 5176 20778 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21726 5216 21732 5228
rect 21687 5188 21732 5216
rect 21085 5179 21143 5185
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 25961 5219 26019 5225
rect 25961 5185 25973 5219
rect 26007 5216 26019 5219
rect 26970 5216 26976 5228
rect 26007 5188 26976 5216
rect 26007 5185 26019 5188
rect 25961 5179 26019 5185
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 27246 5216 27252 5228
rect 27207 5188 27252 5216
rect 27246 5176 27252 5188
rect 27304 5176 27310 5228
rect 28166 5176 28172 5228
rect 28224 5216 28230 5228
rect 31772 5225 31800 5256
rect 32125 5253 32137 5256
rect 32171 5284 32183 5287
rect 32214 5284 32220 5296
rect 32171 5256 32220 5284
rect 32171 5253 32183 5256
rect 32125 5247 32183 5253
rect 32214 5244 32220 5256
rect 32272 5244 32278 5296
rect 33229 5287 33287 5293
rect 33229 5253 33241 5287
rect 33275 5284 33287 5287
rect 34698 5284 34704 5296
rect 33275 5256 34704 5284
rect 33275 5253 33287 5256
rect 33229 5247 33287 5253
rect 34698 5244 34704 5256
rect 34756 5284 34762 5296
rect 36265 5287 36323 5293
rect 36265 5284 36277 5287
rect 34756 5256 36277 5284
rect 34756 5244 34762 5256
rect 36265 5253 36277 5256
rect 36311 5284 36323 5287
rect 36630 5284 36636 5296
rect 36311 5256 36636 5284
rect 36311 5253 36323 5256
rect 36265 5247 36323 5253
rect 36630 5244 36636 5256
rect 36688 5244 36694 5296
rect 29641 5219 29699 5225
rect 29641 5216 29653 5219
rect 28224 5188 29653 5216
rect 28224 5176 28230 5188
rect 29641 5185 29653 5188
rect 29687 5185 29699 5219
rect 31757 5219 31815 5225
rect 31757 5216 31769 5219
rect 29641 5179 29699 5185
rect 30484 5188 31769 5216
rect 30484 5160 30512 5188
rect 31757 5185 31769 5188
rect 31803 5185 31815 5219
rect 31757 5179 31815 5185
rect 31846 5176 31852 5228
rect 31904 5216 31910 5228
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31904 5188 32321 5216
rect 31904 5176 31910 5188
rect 32309 5185 32321 5188
rect 32355 5216 32367 5219
rect 32950 5216 32956 5228
rect 32355 5188 32956 5216
rect 32355 5185 32367 5188
rect 32309 5179 32367 5185
rect 32950 5176 32956 5188
rect 33008 5176 33014 5228
rect 34974 5216 34980 5228
rect 34935 5188 34980 5216
rect 34974 5176 34980 5188
rect 35032 5176 35038 5228
rect 35250 5216 35256 5228
rect 35211 5188 35256 5216
rect 35250 5176 35256 5188
rect 35308 5176 35314 5228
rect 35986 5176 35992 5228
rect 36044 5216 36050 5228
rect 36817 5219 36875 5225
rect 36817 5216 36829 5219
rect 36044 5188 36829 5216
rect 36044 5176 36050 5188
rect 36817 5185 36829 5188
rect 36863 5185 36875 5219
rect 36817 5179 36875 5185
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 18046 5108 18052 5120
rect 18104 5148 18110 5160
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 18104 5120 18521 5148
rect 18104 5108 18110 5120
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 19150 5148 19156 5160
rect 19111 5120 19156 5148
rect 18509 5111 18567 5117
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 19702 5148 19708 5160
rect 19291 5120 19708 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 24302 5148 24308 5160
rect 23707 5120 24308 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24302 5108 24308 5120
rect 24360 5108 24366 5160
rect 30377 5151 30435 5157
rect 30377 5117 30389 5151
rect 30423 5148 30435 5151
rect 30466 5148 30472 5160
rect 30423 5120 30472 5148
rect 30423 5117 30435 5120
rect 30377 5111 30435 5117
rect 30466 5108 30472 5120
rect 30524 5108 30530 5160
rect 30834 5148 30840 5160
rect 30795 5120 30840 5148
rect 30834 5108 30840 5120
rect 30892 5148 30898 5160
rect 31297 5151 31355 5157
rect 31297 5148 31309 5151
rect 30892 5120 31309 5148
rect 30892 5108 30898 5120
rect 31297 5117 31309 5120
rect 31343 5117 31355 5151
rect 31297 5111 31355 5117
rect 13903 5083 13961 5089
rect 13903 5049 13915 5083
rect 13949 5049 13961 5083
rect 15378 5080 15384 5092
rect 15339 5052 15384 5080
rect 13903 5043 13961 5049
rect 15378 5040 15384 5052
rect 15436 5040 15442 5092
rect 15473 5083 15531 5089
rect 15473 5049 15485 5083
rect 15519 5080 15531 5083
rect 15838 5080 15844 5092
rect 15519 5052 15844 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 11882 5012 11888 5024
rect 10980 4984 11888 5012
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 14461 5015 14519 5021
rect 14461 4981 14473 5015
rect 14507 5012 14519 5015
rect 15488 5012 15516 5043
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 19168 5080 19196 5108
rect 19566 5083 19624 5089
rect 19566 5080 19578 5083
rect 19168 5052 19578 5080
rect 19566 5049 19578 5052
rect 19612 5049 19624 5083
rect 21177 5083 21235 5089
rect 19566 5043 19624 5049
rect 20456 5052 21036 5080
rect 14507 4984 15516 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 17000 4984 17325 5012
rect 17000 4972 17006 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17313 4975 17371 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 20456 5021 20484 5052
rect 20165 5015 20223 5021
rect 20165 4981 20177 5015
rect 20211 5012 20223 5015
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 20211 4984 20453 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 20806 5012 20812 5024
rect 20588 4984 20812 5012
rect 20588 4972 20594 4984
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 21008 5012 21036 5052
rect 21177 5049 21189 5083
rect 21223 5049 21235 5083
rect 21177 5043 21235 5049
rect 23477 5083 23535 5089
rect 23477 5049 23489 5083
rect 23523 5080 23535 5083
rect 24023 5083 24081 5089
rect 24023 5080 24035 5083
rect 23523 5052 24035 5080
rect 23523 5049 23535 5052
rect 23477 5043 23535 5049
rect 24023 5049 24035 5052
rect 24069 5080 24081 5083
rect 24854 5080 24860 5092
rect 24069 5052 24860 5080
rect 24069 5049 24081 5052
rect 24023 5043 24081 5049
rect 21192 5012 21220 5043
rect 24854 5040 24860 5052
rect 24912 5040 24918 5092
rect 25406 5080 25412 5092
rect 25367 5052 25412 5080
rect 25406 5040 25412 5052
rect 25464 5040 25470 5092
rect 26605 5083 26663 5089
rect 26605 5049 26617 5083
rect 26651 5080 26663 5083
rect 27065 5083 27123 5089
rect 27065 5080 27077 5083
rect 26651 5052 27077 5080
rect 26651 5049 26663 5052
rect 26605 5043 26663 5049
rect 27065 5049 27077 5052
rect 27111 5080 27123 5083
rect 28997 5083 29055 5089
rect 28997 5080 29009 5083
rect 27111 5052 29009 5080
rect 27111 5049 27123 5052
rect 27065 5043 27123 5049
rect 28997 5049 29009 5052
rect 29043 5049 29055 5083
rect 29362 5080 29368 5092
rect 29323 5052 29368 5080
rect 28997 5043 29055 5049
rect 22554 5012 22560 5024
rect 21008 4984 21220 5012
rect 22515 4984 22560 5012
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 23106 5012 23112 5024
rect 23067 4984 23112 5012
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 24578 5012 24584 5024
rect 24539 4984 24584 5012
rect 24578 4972 24584 4984
rect 24636 4972 24642 5024
rect 29012 5012 29040 5043
rect 29362 5040 29368 5052
rect 29420 5040 29426 5092
rect 29457 5083 29515 5089
rect 29457 5049 29469 5083
rect 29503 5049 29515 5083
rect 29457 5043 29515 5049
rect 29472 5012 29500 5043
rect 32214 5040 32220 5092
rect 32272 5080 32278 5092
rect 32630 5083 32688 5089
rect 32630 5080 32642 5083
rect 32272 5052 32642 5080
rect 32272 5040 32278 5052
rect 32630 5049 32642 5052
rect 32676 5080 32688 5083
rect 33686 5080 33692 5092
rect 32676 5052 33692 5080
rect 32676 5049 32688 5052
rect 32630 5043 32688 5049
rect 33686 5040 33692 5052
rect 33744 5080 33750 5092
rect 33873 5083 33931 5089
rect 33873 5080 33885 5083
rect 33744 5052 33885 5080
rect 33744 5040 33750 5052
rect 33873 5049 33885 5052
rect 33919 5049 33931 5083
rect 33873 5043 33931 5049
rect 35066 5040 35072 5092
rect 35124 5080 35130 5092
rect 35124 5052 35169 5080
rect 35124 5040 35130 5052
rect 36354 5040 36360 5092
rect 36412 5080 36418 5092
rect 36541 5083 36599 5089
rect 36541 5080 36553 5083
rect 36412 5052 36553 5080
rect 36412 5040 36418 5052
rect 36541 5049 36553 5052
rect 36587 5049 36599 5083
rect 36541 5043 36599 5049
rect 36630 5040 36636 5092
rect 36688 5080 36694 5092
rect 36688 5052 36733 5080
rect 36688 5040 36694 5052
rect 29012 4984 29500 5012
rect 30374 4972 30380 5024
rect 30432 5012 30438 5024
rect 30653 5015 30711 5021
rect 30653 5012 30665 5015
rect 30432 4984 30665 5012
rect 30432 4972 30438 4984
rect 30653 4981 30665 4984
rect 30699 4981 30711 5015
rect 30653 4975 30711 4981
rect 30926 4972 30932 5024
rect 30984 5012 30990 5024
rect 31021 5015 31079 5021
rect 31021 5012 31033 5015
rect 30984 4984 31033 5012
rect 30984 4972 30990 4984
rect 31021 4981 31033 4984
rect 31067 4981 31079 5015
rect 31021 4975 31079 4981
rect 34701 5015 34759 5021
rect 34701 4981 34713 5015
rect 34747 5012 34759 5015
rect 35084 5012 35112 5040
rect 34747 4984 35112 5012
rect 34747 4981 34759 4984
rect 34701 4975 34759 4981
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1854 4808 1860 4820
rect 1719 4780 1860 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6086 4808 6092 4820
rect 5859 4780 6092 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 12158 4808 12164 4820
rect 12119 4780 12164 4808
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12529 4811 12587 4817
rect 12529 4777 12541 4811
rect 12575 4808 12587 4811
rect 12618 4808 12624 4820
rect 12575 4780 12624 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 12618 4768 12624 4780
rect 12676 4808 12682 4820
rect 13998 4808 14004 4820
rect 12676 4780 13216 4808
rect 13959 4780 14004 4808
rect 12676 4768 12682 4780
rect 2127 4743 2185 4749
rect 2127 4709 2139 4743
rect 2173 4740 2185 4743
rect 2406 4740 2412 4752
rect 2173 4712 2412 4740
rect 2173 4709 2185 4712
rect 2127 4703 2185 4709
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 3602 4700 3608 4752
rect 3660 4740 3666 4752
rect 3970 4740 3976 4752
rect 3660 4712 3976 4740
rect 3660 4700 3666 4712
rect 3970 4700 3976 4712
rect 4028 4740 4034 4752
rect 4249 4743 4307 4749
rect 4249 4740 4261 4743
rect 4028 4712 4261 4740
rect 4028 4700 4034 4712
rect 4249 4709 4261 4712
rect 4295 4740 4307 4743
rect 5077 4743 5135 4749
rect 5077 4740 5089 4743
rect 4295 4712 5089 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 5077 4709 5089 4712
rect 5123 4709 5135 4743
rect 5077 4703 5135 4709
rect 8110 4700 8116 4752
rect 8168 4749 8174 4752
rect 8168 4743 8216 4749
rect 8168 4709 8170 4743
rect 8204 4709 8216 4743
rect 9214 4740 9220 4752
rect 8168 4703 8216 4709
rect 8772 4712 9220 4740
rect 8168 4700 8174 4703
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6638 4672 6644 4684
rect 6595 4644 6644 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 6822 4672 6828 4684
rect 6783 4644 6828 4672
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7834 4672 7840 4684
rect 7795 4644 7840 4672
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8772 4681 8800 4712
rect 9214 4700 9220 4712
rect 9272 4740 9278 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9272 4712 9873 4740
rect 9272 4700 9278 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 9861 4703 9919 4709
rect 10413 4743 10471 4749
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 10502 4740 10508 4752
rect 10459 4712 10508 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 11603 4743 11661 4749
rect 11603 4709 11615 4743
rect 11649 4740 11661 4743
rect 11974 4740 11980 4752
rect 11649 4712 11980 4740
rect 11649 4709 11661 4712
rect 11603 4703 11661 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 12802 4740 12808 4752
rect 12763 4712 12808 4740
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 13078 4740 13084 4752
rect 13039 4712 13084 4740
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 13188 4749 13216 4780
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 20530 4808 20536 4820
rect 19659 4780 20536 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 21910 4808 21916 4820
rect 21871 4780 21916 4808
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 23566 4768 23572 4820
rect 23624 4768 23630 4820
rect 24302 4808 24308 4820
rect 24263 4780 24308 4808
rect 24302 4768 24308 4780
rect 24360 4808 24366 4820
rect 24949 4811 25007 4817
rect 24949 4808 24961 4811
rect 24360 4780 24961 4808
rect 24360 4768 24366 4780
rect 24949 4777 24961 4780
rect 24995 4777 25007 4811
rect 26326 4808 26332 4820
rect 26287 4780 26332 4808
rect 24949 4771 25007 4777
rect 26326 4768 26332 4780
rect 26384 4768 26390 4820
rect 29362 4808 29368 4820
rect 29323 4780 29368 4808
rect 29362 4768 29368 4780
rect 29420 4768 29426 4820
rect 32950 4808 32956 4820
rect 32911 4780 32956 4808
rect 32950 4768 32956 4780
rect 33008 4768 33014 4820
rect 34974 4808 34980 4820
rect 34935 4780 34980 4808
rect 34974 4768 34980 4780
rect 35032 4768 35038 4820
rect 35066 4768 35072 4820
rect 35124 4808 35130 4820
rect 36081 4811 36139 4817
rect 36081 4808 36093 4811
rect 35124 4780 36093 4808
rect 35124 4768 35130 4780
rect 36081 4777 36093 4780
rect 36127 4777 36139 4811
rect 36081 4771 36139 4777
rect 36354 4768 36360 4820
rect 36412 4808 36418 4820
rect 36449 4811 36507 4817
rect 36449 4808 36461 4811
rect 36412 4780 36461 4808
rect 36412 4768 36418 4780
rect 36449 4777 36461 4780
rect 36495 4777 36507 4811
rect 36449 4771 36507 4777
rect 13173 4743 13231 4749
rect 13173 4709 13185 4743
rect 13219 4709 13231 4743
rect 13173 4703 13231 4709
rect 13538 4700 13544 4752
rect 13596 4740 13602 4752
rect 14182 4740 14188 4752
rect 13596 4712 14188 4740
rect 13596 4700 13602 4712
rect 14182 4700 14188 4712
rect 14240 4740 14246 4752
rect 14369 4743 14427 4749
rect 14369 4740 14381 4743
rect 14240 4712 14381 4740
rect 14240 4700 14246 4712
rect 14369 4709 14381 4712
rect 14415 4709 14427 4743
rect 14369 4703 14427 4709
rect 19055 4743 19113 4749
rect 19055 4709 19067 4743
rect 19101 4740 19113 4743
rect 19150 4740 19156 4752
rect 19101 4712 19156 4740
rect 19101 4709 19113 4712
rect 19055 4703 19113 4709
rect 19150 4700 19156 4712
rect 19208 4700 19214 4752
rect 19886 4740 19892 4752
rect 19847 4712 19892 4740
rect 19886 4700 19892 4712
rect 19944 4700 19950 4752
rect 20717 4743 20775 4749
rect 20717 4709 20729 4743
rect 20763 4740 20775 4743
rect 20806 4740 20812 4752
rect 20763 4712 20812 4740
rect 20763 4709 20775 4712
rect 20717 4703 20775 4709
rect 20806 4700 20812 4712
rect 20864 4740 20870 4752
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 20864 4712 21097 4740
rect 20864 4700 20870 4712
rect 21085 4709 21097 4712
rect 21131 4709 21143 4743
rect 21085 4703 21143 4709
rect 21637 4743 21695 4749
rect 21637 4709 21649 4743
rect 21683 4740 21695 4743
rect 21726 4740 21732 4752
rect 21683 4712 21732 4740
rect 21683 4709 21695 4712
rect 21637 4703 21695 4709
rect 21726 4700 21732 4712
rect 21784 4700 21790 4752
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4641 8815 4675
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 8757 4635 8815 4641
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15838 4672 15844 4684
rect 15799 4644 15844 4672
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 16316 4644 16865 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 2590 4604 2596 4616
rect 1811 4576 2596 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 4154 4604 4160 4616
rect 3559 4576 4160 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4798 4604 4804 4616
rect 4759 4576 4804 4604
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 7055 4576 7297 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7285 4573 7297 4576
rect 7331 4604 7343 4607
rect 7466 4604 7472 4616
rect 7331 4576 7472 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 9766 4604 9772 4616
rect 9727 4576 9772 4604
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 11238 4604 11244 4616
rect 11199 4576 11244 4604
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 13446 4604 13452 4616
rect 13407 4576 13452 4604
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4604 15715 4607
rect 16316 4604 16344 4644
rect 16853 4641 16865 4644
rect 16899 4672 16911 4675
rect 17770 4672 17776 4684
rect 16899 4644 17776 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 17770 4632 17776 4644
rect 17828 4632 17834 4684
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 23584 4681 23612 4768
rect 24026 4740 24032 4752
rect 23987 4712 24032 4740
rect 24026 4700 24032 4712
rect 24084 4740 24090 4752
rect 24673 4743 24731 4749
rect 24673 4740 24685 4743
rect 24084 4712 24685 4740
rect 24084 4700 24090 4712
rect 24673 4709 24685 4712
rect 24719 4709 24731 4743
rect 24673 4703 24731 4709
rect 26234 4700 26240 4752
rect 26292 4740 26298 4752
rect 26697 4743 26755 4749
rect 26697 4740 26709 4743
rect 26292 4712 26709 4740
rect 26292 4700 26298 4712
rect 26697 4709 26709 4712
rect 26743 4709 26755 4743
rect 28258 4740 28264 4752
rect 28219 4712 28264 4740
rect 26697 4703 26755 4709
rect 28258 4700 28264 4712
rect 28316 4700 28322 4752
rect 31202 4740 31208 4752
rect 31163 4712 31208 4740
rect 31202 4700 31208 4712
rect 31260 4700 31266 4752
rect 33686 4700 33692 4752
rect 33744 4749 33750 4752
rect 33744 4743 33792 4749
rect 33744 4709 33746 4743
rect 33780 4740 33792 4743
rect 35482 4743 35540 4749
rect 35482 4740 35494 4743
rect 33780 4712 35494 4740
rect 33780 4709 33792 4712
rect 33744 4703 33792 4709
rect 35482 4709 35494 4712
rect 35528 4740 35540 4743
rect 35894 4740 35900 4752
rect 35528 4712 35900 4740
rect 35528 4709 35540 4712
rect 35482 4703 35540 4709
rect 33744 4700 33750 4703
rect 35894 4700 35900 4712
rect 35952 4700 35958 4752
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 18380 4644 18705 4672
rect 18380 4632 18386 4644
rect 18693 4641 18705 4644
rect 18739 4672 18751 4675
rect 20257 4675 20315 4681
rect 20257 4672 20269 4675
rect 18739 4644 20269 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 20257 4641 20269 4644
rect 20303 4641 20315 4675
rect 20257 4635 20315 4641
rect 23569 4675 23627 4681
rect 23569 4641 23581 4675
rect 23615 4641 23627 4675
rect 23750 4672 23756 4684
rect 23711 4644 23756 4672
rect 23569 4635 23627 4641
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 24946 4672 24952 4684
rect 24907 4644 24952 4672
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 25317 4675 25375 4681
rect 25317 4641 25329 4675
rect 25363 4641 25375 4675
rect 25317 4635 25375 4641
rect 15703 4576 16344 4604
rect 16393 4607 16451 4613
rect 15703 4573 15715 4576
rect 15657 4567 15715 4573
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16666 4604 16672 4616
rect 16439 4576 16672 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16666 4564 16672 4576
rect 16724 4604 16730 4616
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 16724 4576 17233 4604
rect 16724 4564 16730 4576
rect 17221 4573 17233 4576
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4604 21051 4607
rect 21266 4604 21272 4616
rect 21039 4576 21272 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 21266 4564 21272 4576
rect 21324 4604 21330 4616
rect 22554 4604 22560 4616
rect 21324 4576 22560 4604
rect 21324 4564 21330 4576
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 23768 4604 23796 4632
rect 25130 4604 25136 4616
rect 23768 4576 25136 4604
rect 25130 4564 25136 4576
rect 25188 4604 25194 4616
rect 25332 4604 25360 4635
rect 30374 4632 30380 4684
rect 30432 4672 30438 4684
rect 30469 4675 30527 4681
rect 30469 4672 30481 4675
rect 30432 4644 30481 4672
rect 30432 4632 30438 4644
rect 30469 4641 30481 4644
rect 30515 4641 30527 4675
rect 30926 4672 30932 4684
rect 30887 4644 30932 4672
rect 30469 4635 30527 4641
rect 30926 4632 30932 4644
rect 30984 4632 30990 4684
rect 25188 4576 25360 4604
rect 25188 4564 25194 4576
rect 26142 4564 26148 4616
rect 26200 4604 26206 4616
rect 26605 4607 26663 4613
rect 26605 4604 26617 4607
rect 26200 4576 26617 4604
rect 26200 4564 26206 4576
rect 26605 4573 26617 4576
rect 26651 4604 26663 4607
rect 27246 4604 27252 4616
rect 26651 4576 27252 4604
rect 26651 4573 26663 4576
rect 26605 4567 26663 4573
rect 27246 4564 27252 4576
rect 27304 4564 27310 4616
rect 28166 4604 28172 4616
rect 28127 4576 28172 4604
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28810 4604 28816 4616
rect 28771 4576 28816 4604
rect 28810 4564 28816 4576
rect 28868 4564 28874 4616
rect 32122 4604 32128 4616
rect 32083 4576 32128 4604
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 33413 4607 33471 4613
rect 33413 4573 33425 4607
rect 33459 4604 33471 4607
rect 33962 4604 33968 4616
rect 33459 4576 33968 4604
rect 33459 4573 33471 4576
rect 33413 4567 33471 4573
rect 33962 4564 33968 4576
rect 34020 4564 34026 4616
rect 35158 4604 35164 4616
rect 35119 4576 35164 4604
rect 35158 4564 35164 4576
rect 35216 4564 35222 4616
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 8846 4536 8852 4548
rect 8352 4508 8852 4536
rect 8352 4496 8358 4508
rect 8846 4496 8852 4508
rect 8904 4536 8910 4548
rect 9401 4539 9459 4545
rect 9401 4536 9413 4539
rect 8904 4508 9413 4536
rect 8904 4496 8910 4508
rect 9401 4505 9413 4508
rect 9447 4536 9459 4539
rect 9582 4536 9588 4548
rect 9447 4508 9588 4536
rect 9447 4505 9459 4508
rect 9401 4499 9459 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 18046 4536 18052 4548
rect 16960 4508 18052 4536
rect 16960 4480 16988 4508
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 27154 4536 27160 4548
rect 27067 4508 27160 4536
rect 27154 4496 27160 4508
rect 27212 4536 27218 4548
rect 28828 4536 28856 4564
rect 32582 4536 32588 4548
rect 27212 4508 28856 4536
rect 32543 4508 32588 4536
rect 27212 4496 27218 4508
rect 32582 4496 32588 4508
rect 32640 4496 32646 4548
rect 2682 4468 2688 4480
rect 2643 4440 2688 4468
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 8110 4468 8116 4480
rect 7791 4440 8116 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8260 4440 9045 4468
rect 8260 4428 8266 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 10778 4468 10784 4480
rect 10739 4440 10784 4468
rect 9033 4431 9091 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 15102 4468 15108 4480
rect 15063 4440 15108 4468
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16669 4471 16727 4477
rect 16669 4468 16681 4471
rect 16356 4440 16681 4468
rect 16356 4428 16362 4440
rect 16669 4437 16681 4440
rect 16715 4468 16727 4471
rect 16942 4468 16948 4480
rect 16715 4440 16948 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16942 4428 16948 4440
rect 17000 4477 17006 4480
rect 17000 4471 17049 4477
rect 17000 4437 17003 4471
rect 17037 4437 17049 4471
rect 17126 4468 17132 4480
rect 17087 4440 17132 4468
rect 17000 4431 17049 4437
rect 17000 4428 17006 4431
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 17310 4468 17316 4480
rect 17271 4440 17316 4468
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 18230 4428 18236 4480
rect 18288 4468 18294 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 18288 4440 18429 4468
rect 18288 4428 18294 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 18417 4431 18475 4437
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 28350 4468 28356 4480
rect 22704 4440 28356 4468
rect 22704 4428 22710 4440
rect 28350 4428 28356 4440
rect 28408 4468 28414 4480
rect 28718 4468 28724 4480
rect 28408 4440 28724 4468
rect 28408 4428 28414 4440
rect 28718 4428 28724 4440
rect 28776 4428 28782 4480
rect 31478 4468 31484 4480
rect 31439 4440 31484 4468
rect 31478 4428 31484 4440
rect 31536 4428 31542 4480
rect 34333 4471 34391 4477
rect 34333 4437 34345 4471
rect 34379 4468 34391 4471
rect 34606 4468 34612 4480
rect 34379 4440 34612 4468
rect 34379 4437 34391 4440
rect 34333 4431 34391 4437
rect 34606 4428 34612 4440
rect 34664 4428 34670 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 2406 4264 2412 4276
rect 2367 4236 2412 4264
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 3970 4264 3976 4276
rect 3931 4236 3976 4264
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 6365 4267 6423 4273
rect 6365 4233 6377 4267
rect 6411 4264 6423 4267
rect 6822 4264 6828 4276
rect 6411 4236 6828 4264
rect 6411 4233 6423 4236
rect 6365 4227 6423 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 11974 4264 11980 4276
rect 11931 4236 11980 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12805 4267 12863 4273
rect 12805 4233 12817 4267
rect 12851 4264 12863 4267
rect 13906 4264 13912 4276
rect 12851 4236 13912 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 18187 4267 18245 4273
rect 18187 4264 18199 4267
rect 18104 4236 18199 4264
rect 18104 4224 18110 4236
rect 18187 4233 18199 4236
rect 18233 4233 18245 4267
rect 18187 4227 18245 4233
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 21266 4264 21272 4276
rect 21227 4236 21272 4264
rect 20901 4227 20959 4233
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 21637 4267 21695 4273
rect 21637 4264 21649 4267
rect 21416 4236 21649 4264
rect 21416 4224 21422 4236
rect 21637 4233 21649 4236
rect 21683 4264 21695 4267
rect 22278 4264 22284 4276
rect 21683 4236 22284 4264
rect 21683 4233 21695 4236
rect 21637 4227 21695 4233
rect 22278 4224 22284 4236
rect 22336 4224 22342 4276
rect 23385 4267 23443 4273
rect 23385 4233 23397 4267
rect 23431 4264 23443 4267
rect 23474 4264 23480 4276
rect 23431 4236 23480 4264
rect 23431 4233 23443 4236
rect 23385 4227 23443 4233
rect 23474 4224 23480 4236
rect 23532 4224 23538 4276
rect 27617 4267 27675 4273
rect 27617 4233 27629 4267
rect 27663 4264 27675 4267
rect 28169 4267 28227 4273
rect 28169 4264 28181 4267
rect 27663 4236 28181 4264
rect 27663 4233 27675 4236
rect 27617 4227 27675 4233
rect 28169 4233 28181 4236
rect 28215 4264 28227 4267
rect 28258 4264 28264 4276
rect 28215 4236 28264 4264
rect 28215 4233 28227 4236
rect 28169 4227 28227 4233
rect 28258 4224 28264 4236
rect 28316 4224 28322 4276
rect 30374 4224 30380 4276
rect 30432 4264 30438 4276
rect 30469 4267 30527 4273
rect 30469 4264 30481 4267
rect 30432 4236 30481 4264
rect 30432 4224 30438 4236
rect 30469 4233 30481 4236
rect 30515 4264 30527 4267
rect 32214 4264 32220 4276
rect 30515 4236 32220 4264
rect 30515 4233 30527 4236
rect 30469 4227 30527 4233
rect 32214 4224 32220 4236
rect 32272 4224 32278 4276
rect 33686 4264 33692 4276
rect 33647 4236 33692 4264
rect 33686 4224 33692 4236
rect 33744 4224 33750 4276
rect 35894 4264 35900 4276
rect 35855 4236 35900 4264
rect 35894 4224 35900 4236
rect 35952 4224 35958 4276
rect 35986 4224 35992 4276
rect 36044 4264 36050 4276
rect 36265 4267 36323 4273
rect 36265 4264 36277 4267
rect 36044 4236 36277 4264
rect 36044 4224 36050 4236
rect 36265 4233 36277 4236
rect 36311 4233 36323 4267
rect 36265 4227 36323 4233
rect 3234 4196 3240 4208
rect 2700 4168 3240 4196
rect 2700 4137 2728 4168
rect 3234 4156 3240 4168
rect 3292 4156 3298 4208
rect 4798 4196 4804 4208
rect 4172 4168 4804 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3016 4100 3341 4128
rect 3016 4088 3022 4100
rect 3329 4097 3341 4100
rect 3375 4128 3387 4131
rect 4172 4128 4200 4168
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 6638 4196 6644 4208
rect 5675 4168 6644 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 16574 4196 16580 4208
rect 16535 4168 16580 4196
rect 16574 4156 16580 4168
rect 16632 4196 16638 4208
rect 17126 4196 17132 4208
rect 16632 4168 17132 4196
rect 16632 4156 16638 4168
rect 17126 4156 17132 4168
rect 17184 4196 17190 4208
rect 17313 4199 17371 4205
rect 17313 4196 17325 4199
rect 17184 4168 17325 4196
rect 17184 4156 17190 4168
rect 17313 4165 17325 4168
rect 17359 4196 17371 4199
rect 17586 4196 17592 4208
rect 17359 4168 17592 4196
rect 17359 4165 17371 4168
rect 17313 4159 17371 4165
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 23750 4196 23756 4208
rect 23492 4168 23756 4196
rect 3375 4100 4200 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4304 4100 4537 4128
rect 4304 4088 4310 4100
rect 4525 4097 4537 4100
rect 4571 4128 4583 4131
rect 4706 4128 4712 4140
rect 4571 4100 4712 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7524 4100 7849 4128
rect 7524 4088 7530 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 11330 4128 11336 4140
rect 11291 4100 11336 4128
rect 7837 4091 7895 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11422 4088 11428 4140
rect 11480 4128 11486 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11480 4100 11529 4128
rect 11480 4088 11486 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 14734 4128 14740 4140
rect 14695 4100 14740 4128
rect 11517 4091 11575 4097
rect 14734 4088 14740 4100
rect 14792 4128 14798 4140
rect 15286 4128 15292 4140
rect 14792 4100 15292 4128
rect 14792 4088 14798 4100
rect 1648 4063 1706 4069
rect 1648 4029 1660 4063
rect 1694 4060 1706 4063
rect 5721 4063 5779 4069
rect 1694 4032 2176 4060
rect 1694 4029 1706 4032
rect 1648 4023 1706 4029
rect 2148 4001 2176 4032
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6086 4060 6092 4072
rect 5767 4032 6092 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 10689 4063 10747 4069
rect 6871 4032 7420 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 2498 3992 2504 4004
rect 2179 3964 2504 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 2777 3995 2835 4001
rect 2777 3961 2789 3995
rect 2823 3961 2835 3995
rect 4246 3992 4252 4004
rect 4207 3964 4252 3992
rect 2777 3955 2835 3961
rect 1719 3927 1777 3933
rect 1719 3893 1731 3927
rect 1765 3924 1777 3927
rect 1946 3924 1952 3936
rect 1765 3896 1952 3924
rect 1765 3893 1777 3896
rect 1719 3887 1777 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2792 3924 2820 3955
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 4341 3995 4399 4001
rect 4341 3961 4353 3995
rect 4387 3961 4399 3995
rect 4341 3955 4399 3961
rect 2866 3924 2872 3936
rect 2779 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3924 2930 3936
rect 3697 3927 3755 3933
rect 3697 3924 3709 3927
rect 2924 3896 3709 3924
rect 2924 3884 2930 3896
rect 3697 3893 3709 3896
rect 3743 3924 3755 3927
rect 4356 3924 4384 3955
rect 5810 3952 5816 4004
rect 5868 3992 5874 4004
rect 7282 3992 7288 4004
rect 5868 3964 7288 3992
rect 5868 3952 5874 3964
rect 5258 3924 5264 3936
rect 3743 3896 4384 3924
rect 5219 3896 5264 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3924 5966 3936
rect 6454 3924 6460 3936
rect 5960 3896 6460 3924
rect 5960 3884 5966 3896
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 7024 3933 7052 3964
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 7392 3936 7420 4032
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 10689 4023 10747 4029
rect 11164 4032 11253 4060
rect 7742 3992 7748 4004
rect 7703 3964 7748 3992
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 8199 3995 8257 4001
rect 8199 3961 8211 3995
rect 8245 3961 8257 3995
rect 9582 3992 9588 4004
rect 9543 3964 9588 3992
rect 8199 3955 8257 3961
rect 7009 3927 7067 3933
rect 7009 3893 7021 3927
rect 7055 3893 7067 3927
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 7009 3887 7067 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7760 3924 7788 3952
rect 8110 3924 8116 3936
rect 7760 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3924 8174 3936
rect 8220 3924 8248 3955
rect 9582 3952 9588 3964
rect 9640 3952 9646 4004
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10704 3992 10732 4023
rect 10778 3992 10784 4004
rect 9999 3964 10784 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10778 3952 10784 3964
rect 10836 3992 10842 4004
rect 11054 3992 11060 4004
rect 10836 3964 11060 3992
rect 10836 3952 10842 3964
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 8754 3924 8760 3936
rect 8168 3896 8248 3924
rect 8715 3896 8760 3924
rect 8168 3884 8174 3896
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3924 10290 3936
rect 11164 3924 11192 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4060 13231 4063
rect 13538 4060 13544 4072
rect 13219 4032 13544 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 13814 4060 13820 4072
rect 13775 4032 13820 4060
rect 13814 4020 13820 4032
rect 13872 4060 13878 4072
rect 14936 4069 14964 4100
rect 15286 4088 15292 4100
rect 15344 4128 15350 4140
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 15344 4100 15761 4128
rect 15344 4088 15350 4100
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16448 4131 16506 4137
rect 16448 4128 16460 4131
rect 16356 4100 16460 4128
rect 16356 4088 16362 4100
rect 16448 4097 16460 4100
rect 16494 4097 16506 4131
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 16448 4091 16506 4097
rect 16666 4088 16672 4100
rect 16724 4128 16730 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 16724 4100 17785 4128
rect 16724 4088 16730 4100
rect 17773 4097 17785 4100
rect 17819 4128 17831 4131
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 17819 4100 18429 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18417 4097 18429 4100
rect 18463 4097 18475 4131
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 18417 4091 18475 4097
rect 18524 4100 19441 4128
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13872 4032 14289 4060
rect 13872 4020 13878 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4029 14979 4063
rect 15102 4060 15108 4072
rect 15063 4032 15108 4060
rect 14921 4023 14979 4029
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 18230 4020 18236 4072
rect 18288 4069 18294 4072
rect 18288 4063 18337 4069
rect 18288 4029 18291 4063
rect 18325 4060 18337 4063
rect 18524 4060 18552 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 19886 4088 19892 4140
rect 19944 4128 19950 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19944 4100 19993 4128
rect 19944 4088 19950 4100
rect 19981 4097 19993 4100
rect 20027 4128 20039 4131
rect 20622 4128 20628 4140
rect 20027 4100 20628 4128
rect 20027 4097 20039 4100
rect 19981 4091 20039 4097
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4128 23075 4131
rect 23382 4128 23388 4140
rect 23063 4100 23388 4128
rect 23063 4097 23075 4100
rect 23017 4091 23075 4097
rect 23382 4088 23388 4100
rect 23440 4128 23446 4140
rect 23492 4128 23520 4168
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 24946 4196 24952 4208
rect 24872 4168 24952 4196
rect 23440 4100 23520 4128
rect 24489 4131 24547 4137
rect 23440 4088 23446 4100
rect 24489 4097 24501 4131
rect 24535 4128 24547 4131
rect 24872 4128 24900 4168
rect 24946 4156 24952 4168
rect 25004 4156 25010 4208
rect 35084 4168 35388 4196
rect 30926 4128 30932 4140
rect 24535 4100 24900 4128
rect 30887 4100 30932 4128
rect 24535 4097 24547 4100
rect 24489 4091 24547 4097
rect 30926 4088 30932 4100
rect 30984 4128 30990 4140
rect 32401 4131 32459 4137
rect 32401 4128 32413 4131
rect 30984 4100 32413 4128
rect 30984 4088 30990 4100
rect 32401 4097 32413 4100
rect 32447 4128 32459 4131
rect 34606 4128 34612 4140
rect 32447 4100 33088 4128
rect 34567 4100 34612 4128
rect 32447 4097 32459 4100
rect 32401 4091 32459 4097
rect 18782 4060 18788 4072
rect 18325 4032 18552 4060
rect 18743 4032 18788 4060
rect 18325 4029 18337 4032
rect 18288 4023 18337 4029
rect 18288 4020 18294 4023
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 21818 4060 21824 4072
rect 21779 4032 21824 4060
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 22186 4060 22192 4072
rect 22147 4032 22192 4060
rect 22186 4020 22192 4032
rect 22244 4020 22250 4072
rect 24949 4063 25007 4069
rect 24949 4029 24961 4063
rect 24995 4060 25007 4063
rect 25498 4060 25504 4072
rect 24995 4032 25504 4060
rect 24995 4029 25007 4032
rect 24949 4023 25007 4029
rect 25498 4020 25504 4032
rect 25556 4020 25562 4072
rect 25869 4063 25927 4069
rect 25869 4029 25881 4063
rect 25915 4060 25927 4063
rect 26234 4060 26240 4072
rect 25915 4032 26240 4060
rect 25915 4029 25927 4032
rect 25869 4023 25927 4029
rect 26234 4020 26240 4032
rect 26292 4020 26298 4072
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26697 4063 26755 4069
rect 26697 4060 26709 4063
rect 26384 4032 26709 4060
rect 26384 4020 26390 4032
rect 26697 4029 26709 4032
rect 26743 4029 26755 4063
rect 29546 4060 29552 4072
rect 29507 4032 29552 4060
rect 26697 4023 26755 4029
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 29914 4060 29920 4072
rect 29875 4032 29920 4060
rect 29914 4020 29920 4032
rect 29972 4020 29978 4072
rect 32582 4060 32588 4072
rect 32543 4032 32588 4060
rect 32582 4020 32588 4032
rect 32640 4020 32646 4072
rect 33060 4069 33088 4100
rect 34606 4088 34612 4100
rect 34664 4088 34670 4140
rect 34977 4131 35035 4137
rect 34977 4097 34989 4131
rect 35023 4128 35035 4131
rect 35084 4128 35112 4168
rect 35250 4128 35256 4140
rect 35023 4100 35112 4128
rect 35211 4100 35256 4128
rect 35023 4097 35035 4100
rect 34977 4091 35035 4097
rect 35250 4088 35256 4100
rect 35308 4088 35314 4140
rect 35360 4128 35388 4168
rect 36004 4128 36032 4224
rect 35360 4100 36032 4128
rect 33045 4063 33103 4069
rect 33045 4029 33057 4063
rect 33091 4029 33103 4063
rect 36446 4060 36452 4072
rect 36407 4032 36452 4060
rect 33045 4023 33103 4029
rect 36446 4020 36452 4032
rect 36504 4060 36510 4072
rect 36998 4060 37004 4072
rect 36504 4032 37004 4060
rect 36504 4020 36510 4032
rect 36998 4020 37004 4032
rect 37056 4020 37062 4072
rect 37550 4020 37556 4072
rect 37608 4069 37614 4072
rect 37608 4063 37646 4069
rect 37634 4060 37646 4063
rect 38013 4063 38071 4069
rect 38013 4060 38025 4063
rect 37634 4032 38025 4060
rect 37634 4029 37646 4032
rect 37608 4023 37646 4029
rect 38013 4029 38025 4032
rect 38059 4029 38071 4063
rect 38013 4023 38071 4029
rect 37608 4020 37614 4023
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12802 3992 12808 4004
rect 12299 3964 12808 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 15194 3952 15200 4004
rect 15252 3992 15258 4004
rect 15473 3995 15531 4001
rect 15473 3992 15485 3995
rect 15252 3964 15485 3992
rect 15252 3952 15258 3964
rect 15473 3961 15485 3964
rect 15519 3992 15531 3995
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 15519 3964 16313 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 16301 3961 16313 3964
rect 16347 3992 16359 3995
rect 16482 3992 16488 4004
rect 16347 3964 16488 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 17034 3992 17040 4004
rect 16995 3964 17040 3992
rect 17034 3952 17040 3964
rect 17092 3952 17098 4004
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 18049 3995 18107 4001
rect 18049 3992 18061 3995
rect 17828 3964 18061 3992
rect 17828 3952 17834 3964
rect 18049 3961 18061 3964
rect 18095 3961 18107 3995
rect 19150 3992 19156 4004
rect 19063 3964 19156 3992
rect 18049 3955 18107 3961
rect 19150 3952 19156 3964
rect 19208 3992 19214 4004
rect 20302 3995 20360 4001
rect 20302 3992 20314 3995
rect 19208 3964 20314 3992
rect 19208 3952 19214 3964
rect 19812 3936 19840 3964
rect 20302 3961 20314 3964
rect 20348 3961 20360 3995
rect 20302 3955 20360 3961
rect 24857 3995 24915 4001
rect 24857 3961 24869 3995
rect 24903 3992 24915 3995
rect 25038 3992 25044 4004
rect 24903 3964 25044 3992
rect 24903 3961 24915 3964
rect 24857 3955 24915 3961
rect 25038 3952 25044 3964
rect 25096 3992 25102 4004
rect 25311 3995 25369 4001
rect 25311 3992 25323 3995
rect 25096 3964 25323 3992
rect 25096 3952 25102 3964
rect 25311 3961 25323 3964
rect 25357 3992 25369 3995
rect 26605 3995 26663 4001
rect 26605 3992 26617 3995
rect 25357 3964 26617 3992
rect 25357 3961 25369 3964
rect 25311 3955 25369 3961
rect 26605 3961 26617 3964
rect 26651 3992 26663 3995
rect 27059 3995 27117 4001
rect 27059 3992 27071 3995
rect 26651 3964 27071 3992
rect 26651 3961 26663 3964
rect 26605 3955 26663 3961
rect 27059 3961 27071 3964
rect 27105 3992 27117 3995
rect 28718 3992 28724 4004
rect 27105 3964 28724 3992
rect 27105 3961 27117 3964
rect 27059 3955 27117 3961
rect 28718 3952 28724 3964
rect 28776 3952 28782 4004
rect 29089 3995 29147 4001
rect 29089 3961 29101 3995
rect 29135 3992 29147 3995
rect 29932 3992 29960 4020
rect 30098 3992 30104 4004
rect 29135 3964 29960 3992
rect 30059 3964 30104 3992
rect 29135 3961 29147 3964
rect 29089 3955 29147 3961
rect 30098 3952 30104 3964
rect 30156 3952 30162 4004
rect 31110 3992 31116 4004
rect 31071 3964 31116 3992
rect 31110 3952 31116 3964
rect 31168 3952 31174 4004
rect 31205 3995 31263 4001
rect 31205 3961 31217 3995
rect 31251 3992 31263 3995
rect 31478 3992 31484 4004
rect 31251 3964 31484 3992
rect 31251 3961 31263 3964
rect 31205 3955 31263 3961
rect 31478 3952 31484 3964
rect 31536 3952 31542 4004
rect 31570 3952 31576 4004
rect 31628 3992 31634 4004
rect 31757 3995 31815 4001
rect 31757 3992 31769 3995
rect 31628 3964 31769 3992
rect 31628 3952 31634 3964
rect 31757 3961 31769 3964
rect 31803 3961 31815 3995
rect 33318 3992 33324 4004
rect 33279 3964 33324 3992
rect 31757 3955 31815 3961
rect 33318 3952 33324 3964
rect 33376 3952 33382 4004
rect 35069 3995 35127 4001
rect 35069 3961 35081 3995
rect 35115 3961 35127 3995
rect 35069 3955 35127 3961
rect 10284 3896 11192 3924
rect 13541 3927 13599 3933
rect 10284 3884 10290 3896
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 13722 3924 13728 3936
rect 13587 3896 13728 3924
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14918 3884 14924 3936
rect 14976 3924 14982 3936
rect 16117 3927 16175 3933
rect 16117 3924 16129 3927
rect 14976 3896 16129 3924
rect 14976 3884 14982 3896
rect 16117 3893 16129 3896
rect 16163 3924 16175 3927
rect 16574 3924 16580 3936
rect 16163 3896 16580 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 19794 3924 19800 3936
rect 19755 3896 19800 3924
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 22005 3927 22063 3933
rect 22005 3893 22017 3927
rect 22051 3924 22063 3927
rect 22186 3924 22192 3936
rect 22051 3896 22192 3924
rect 22051 3893 22063 3896
rect 22005 3887 22063 3893
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 23661 3927 23719 3933
rect 23661 3893 23673 3927
rect 23707 3924 23719 3927
rect 24210 3924 24216 3936
rect 23707 3896 24216 3924
rect 23707 3893 23719 3896
rect 23661 3887 23719 3893
rect 24210 3884 24216 3896
rect 24268 3884 24274 3936
rect 26237 3927 26295 3933
rect 26237 3893 26249 3927
rect 26283 3924 26295 3927
rect 26326 3924 26332 3936
rect 26283 3896 26332 3924
rect 26283 3893 26295 3896
rect 26237 3887 26295 3893
rect 26326 3884 26332 3896
rect 26384 3884 26390 3936
rect 27338 3884 27344 3936
rect 27396 3924 27402 3936
rect 28166 3924 28172 3936
rect 27396 3896 28172 3924
rect 27396 3884 27402 3896
rect 28166 3884 28172 3896
rect 28224 3924 28230 3936
rect 28445 3927 28503 3933
rect 28445 3924 28457 3927
rect 28224 3896 28457 3924
rect 28224 3884 28230 3896
rect 28445 3893 28457 3896
rect 28491 3893 28503 3927
rect 33962 3924 33968 3936
rect 33923 3896 33968 3924
rect 28445 3887 28503 3893
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 34606 3884 34612 3936
rect 34664 3924 34670 3936
rect 35084 3924 35112 3955
rect 34664 3896 35112 3924
rect 36633 3927 36691 3933
rect 34664 3884 34670 3896
rect 36633 3893 36645 3927
rect 36679 3924 36691 3927
rect 36814 3924 36820 3936
rect 36679 3896 36820 3924
rect 36679 3893 36691 3896
rect 36633 3887 36691 3893
rect 36814 3884 36820 3896
rect 36872 3884 36878 3936
rect 37274 3884 37280 3936
rect 37332 3924 37338 3936
rect 37691 3927 37749 3933
rect 37691 3924 37703 3927
rect 37332 3896 37703 3924
rect 37332 3884 37338 3896
rect 37691 3893 37703 3896
rect 37737 3893 37749 3927
rect 37691 3887 37749 3893
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3237 3723 3295 3729
rect 3237 3720 3249 3723
rect 2832 3692 3249 3720
rect 2832 3680 2838 3692
rect 3237 3689 3249 3692
rect 3283 3720 3295 3723
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 3283 3692 4169 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 5166 3720 5172 3732
rect 5127 3692 5172 3720
rect 4157 3683 4215 3689
rect 5166 3680 5172 3692
rect 5224 3720 5230 3732
rect 5350 3720 5356 3732
rect 5224 3692 5356 3720
rect 5224 3680 5230 3692
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6822 3720 6828 3732
rect 6783 3692 6828 3720
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7561 3723 7619 3729
rect 7561 3689 7573 3723
rect 7607 3720 7619 3723
rect 8018 3720 8024 3732
rect 7607 3692 8024 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10134 3720 10140 3732
rect 9907 3692 10140 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 11057 3723 11115 3729
rect 11057 3689 11069 3723
rect 11103 3720 11115 3723
rect 11238 3720 11244 3732
rect 11103 3692 11244 3720
rect 11103 3689 11115 3692
rect 11057 3683 11115 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 12492 3692 13461 3720
rect 12492 3680 12498 3692
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13906 3720 13912 3732
rect 13867 3692 13912 3720
rect 13449 3683 13507 3689
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 15013 3723 15071 3729
rect 15013 3689 15025 3723
rect 15059 3720 15071 3723
rect 15102 3720 15108 3732
rect 15059 3692 15108 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15102 3680 15108 3692
rect 15160 3720 15166 3732
rect 15562 3720 15568 3732
rect 15160 3692 15568 3720
rect 15160 3680 15166 3692
rect 15562 3680 15568 3692
rect 15620 3720 15626 3732
rect 15838 3720 15844 3732
rect 15620 3692 15844 3720
rect 15620 3680 15626 3692
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 17862 3720 17868 3732
rect 17823 3692 17868 3720
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 20165 3723 20223 3729
rect 20165 3720 20177 3723
rect 18340 3692 20177 3720
rect 1762 3612 1768 3664
rect 1820 3652 1826 3664
rect 1943 3655 2001 3661
rect 1943 3652 1955 3655
rect 1820 3624 1955 3652
rect 1820 3612 1826 3624
rect 1943 3621 1955 3624
rect 1989 3652 2001 3655
rect 2406 3652 2412 3664
rect 1989 3624 2412 3652
rect 1989 3621 2001 3624
rect 1943 3615 2001 3621
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 2866 3652 2872 3664
rect 2827 3624 2872 3652
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4246 3652 4252 3664
rect 3927 3624 4252 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4632 3624 6224 3652
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3752 3556 4077 3584
rect 3752 3544 3758 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1670 3516 1676 3528
rect 1627 3488 1676 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 4080 3516 4108 3547
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4632 3593 4660 3624
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4212 3556 4629 3584
rect 4212 3544 4218 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 5810 3584 5816 3596
rect 5771 3556 5816 3584
rect 4617 3547 4675 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6196 3593 6224 3624
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 6270 3584 6276 3596
rect 6227 3556 6276 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6270 3544 6276 3556
rect 6328 3584 6334 3596
rect 6840 3584 6868 3680
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8205 3655 8263 3661
rect 8205 3652 8217 3655
rect 8168 3624 8217 3652
rect 8168 3612 8174 3624
rect 8205 3621 8217 3624
rect 8251 3652 8263 3655
rect 8754 3652 8760 3664
rect 8251 3624 8760 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 10505 3655 10563 3661
rect 10505 3621 10517 3655
rect 10551 3652 10563 3655
rect 10870 3652 10876 3664
rect 10551 3624 10876 3652
rect 10551 3621 10563 3624
rect 10505 3615 10563 3621
rect 10870 3612 10876 3624
rect 10928 3652 10934 3664
rect 12802 3652 12808 3664
rect 10928 3624 11376 3652
rect 12715 3624 12808 3652
rect 10928 3612 10934 3624
rect 11348 3596 11376 3624
rect 12802 3612 12808 3624
rect 12860 3652 12866 3664
rect 13630 3652 13636 3664
rect 12860 3624 13636 3652
rect 12860 3612 12866 3624
rect 13630 3612 13636 3624
rect 13688 3612 13694 3664
rect 16390 3652 16396 3664
rect 16351 3624 16396 3652
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17494 3652 17500 3664
rect 17267 3624 17500 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17494 3612 17500 3624
rect 17552 3652 17558 3664
rect 17770 3652 17776 3664
rect 17552 3624 17776 3652
rect 17552 3612 17558 3624
rect 17770 3612 17776 3624
rect 17828 3652 17834 3664
rect 18233 3655 18291 3661
rect 18233 3652 18245 3655
rect 17828 3624 18245 3652
rect 17828 3612 17834 3624
rect 18233 3621 18245 3624
rect 18279 3621 18291 3655
rect 18233 3615 18291 3621
rect 9674 3584 9680 3596
rect 6328 3556 6868 3584
rect 9635 3556 9680 3584
rect 6328 3544 6334 3556
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 11054 3584 11060 3596
rect 11015 3556 11060 3584
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 11330 3584 11336 3596
rect 11291 3556 11336 3584
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 11606 3584 11612 3596
rect 11567 3556 11612 3584
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 12986 3593 12992 3596
rect 12952 3587 12992 3593
rect 12952 3553 12964 3587
rect 12952 3547 12992 3553
rect 12986 3544 12992 3547
rect 13044 3544 13050 3596
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 16482 3584 16488 3596
rect 15703 3556 16488 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17368 3587 17426 3593
rect 17368 3584 17380 3587
rect 17000 3556 17380 3584
rect 17000 3544 17006 3556
rect 17368 3553 17380 3556
rect 17414 3584 17426 3587
rect 17954 3584 17960 3596
rect 17414 3556 17960 3584
rect 17414 3553 17426 3556
rect 17368 3547 17426 3553
rect 17954 3544 17960 3556
rect 18012 3584 18018 3596
rect 18340 3584 18368 3692
rect 20165 3689 20177 3692
rect 20211 3720 20223 3723
rect 20533 3723 20591 3729
rect 20533 3720 20545 3723
rect 20211 3692 20545 3720
rect 20211 3689 20223 3692
rect 20165 3683 20223 3689
rect 20533 3689 20545 3692
rect 20579 3689 20591 3723
rect 22186 3720 22192 3732
rect 22147 3692 22192 3720
rect 20533 3683 20591 3689
rect 22186 3680 22192 3692
rect 22244 3720 22250 3732
rect 23293 3723 23351 3729
rect 22244 3692 22416 3720
rect 22244 3680 22250 3692
rect 19886 3652 19892 3664
rect 19847 3624 19892 3652
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 20901 3655 20959 3661
rect 20901 3621 20913 3655
rect 20947 3652 20959 3655
rect 21266 3652 21272 3664
rect 20947 3624 21272 3652
rect 20947 3621 20959 3624
rect 20901 3615 20959 3621
rect 21266 3612 21272 3624
rect 21324 3612 21330 3664
rect 19058 3584 19064 3596
rect 18012 3556 18368 3584
rect 18971 3556 19064 3584
rect 18012 3544 18018 3556
rect 19058 3544 19064 3556
rect 19116 3584 19122 3596
rect 19429 3587 19487 3593
rect 19429 3584 19441 3587
rect 19116 3556 19441 3584
rect 19116 3544 19122 3556
rect 19429 3553 19441 3556
rect 19475 3553 19487 3587
rect 19610 3584 19616 3596
rect 19571 3556 19616 3584
rect 19429 3547 19487 3553
rect 5902 3516 5908 3528
rect 4080 3488 5908 3516
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8202 3516 8208 3528
rect 8159 3488 8208 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8754 3516 8760 3528
rect 8715 3488 8760 3516
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 13262 3516 13268 3528
rect 13219 3488 13268 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 13262 3476 13268 3488
rect 13320 3516 13326 3528
rect 14090 3516 14096 3528
rect 13320 3488 14096 3516
rect 13320 3476 13326 3488
rect 14090 3476 14096 3488
rect 14148 3516 14154 3528
rect 14185 3519 14243 3525
rect 14185 3516 14197 3519
rect 14148 3488 14197 3516
rect 14148 3476 14154 3488
rect 14185 3485 14197 3488
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15068 3488 16037 3516
rect 15068 3476 15074 3488
rect 16025 3485 16037 3488
rect 16071 3516 16083 3519
rect 16666 3516 16672 3528
rect 16071 3488 16672 3516
rect 16071 3485 16083 3488
rect 16025 3479 16083 3485
rect 16666 3476 16672 3488
rect 16724 3516 16730 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16724 3488 16865 3516
rect 16724 3476 16730 3488
rect 16853 3485 16865 3488
rect 16899 3516 16911 3519
rect 17126 3516 17132 3528
rect 16899 3488 17132 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 17126 3476 17132 3488
rect 17184 3516 17190 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17184 3488 17601 3516
rect 17184 3476 17190 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 19444 3516 19472 3547
rect 19610 3544 19616 3556
rect 19668 3544 19674 3596
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 20806 3584 20812 3596
rect 20128 3556 20812 3584
rect 20128 3544 20134 3556
rect 20806 3544 20812 3556
rect 20864 3584 20870 3596
rect 22388 3593 22416 3692
rect 23293 3689 23305 3723
rect 23339 3720 23351 3723
rect 23474 3720 23480 3732
rect 23339 3692 23480 3720
rect 23339 3689 23351 3692
rect 23293 3683 23351 3689
rect 23474 3680 23480 3692
rect 23532 3720 23538 3732
rect 25130 3720 25136 3732
rect 23532 3692 24348 3720
rect 25091 3692 25136 3720
rect 23532 3680 23538 3692
rect 22735 3655 22793 3661
rect 22735 3621 22747 3655
rect 22781 3652 22793 3655
rect 23106 3652 23112 3664
rect 22781 3624 23112 3652
rect 22781 3621 22793 3624
rect 22735 3615 22793 3621
rect 23106 3612 23112 3624
rect 23164 3612 23170 3664
rect 24210 3652 24216 3664
rect 24171 3624 24216 3652
rect 24210 3612 24216 3624
rect 24268 3612 24274 3664
rect 24320 3661 24348 3692
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 26234 3720 26240 3732
rect 26195 3692 26240 3720
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 28074 3720 28080 3732
rect 28035 3692 28080 3720
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 30098 3720 30104 3732
rect 30059 3692 30104 3720
rect 30098 3680 30104 3692
rect 30156 3720 30162 3732
rect 31113 3723 31171 3729
rect 30156 3692 30236 3720
rect 30156 3680 30162 3692
rect 24305 3655 24363 3661
rect 24305 3621 24317 3655
rect 24351 3621 24363 3655
rect 24305 3615 24363 3621
rect 25961 3655 26019 3661
rect 25961 3621 25973 3655
rect 26007 3652 26019 3655
rect 26142 3652 26148 3664
rect 26007 3624 26148 3652
rect 26007 3621 26019 3624
rect 25961 3615 26019 3621
rect 26142 3612 26148 3624
rect 26200 3612 26206 3664
rect 26789 3655 26847 3661
rect 26789 3621 26801 3655
rect 26835 3652 26847 3655
rect 26878 3652 26884 3664
rect 26835 3624 26884 3652
rect 26835 3621 26847 3624
rect 26789 3615 26847 3621
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 27338 3652 27344 3664
rect 27299 3624 27344 3652
rect 27338 3612 27344 3624
rect 27396 3612 27402 3664
rect 28531 3655 28589 3661
rect 28531 3621 28543 3655
rect 28577 3652 28589 3655
rect 28718 3652 28724 3664
rect 28577 3624 28724 3652
rect 28577 3621 28589 3624
rect 28531 3615 28589 3621
rect 28718 3612 28724 3624
rect 28776 3612 28782 3664
rect 30208 3593 30236 3692
rect 31113 3689 31125 3723
rect 31159 3720 31171 3723
rect 31478 3720 31484 3732
rect 31159 3692 31484 3720
rect 31159 3689 31171 3692
rect 31113 3683 31171 3689
rect 31478 3680 31484 3692
rect 31536 3680 31542 3732
rect 34609 3723 34667 3729
rect 34609 3689 34621 3723
rect 34655 3720 34667 3723
rect 34655 3692 35664 3720
rect 34655 3689 34667 3692
rect 34609 3683 34667 3689
rect 30466 3612 30472 3664
rect 30524 3661 30530 3664
rect 30524 3655 30572 3661
rect 30524 3621 30526 3655
rect 30560 3621 30572 3655
rect 30524 3615 30572 3621
rect 30524 3612 30530 3615
rect 33778 3612 33784 3664
rect 33836 3652 33842 3664
rect 35636 3661 35664 3692
rect 34010 3655 34068 3661
rect 34010 3652 34022 3655
rect 33836 3624 34022 3652
rect 33836 3612 33842 3624
rect 34010 3621 34022 3624
rect 34056 3621 34068 3655
rect 34010 3615 34068 3621
rect 35621 3655 35679 3661
rect 35621 3621 35633 3655
rect 35667 3652 35679 3655
rect 36262 3652 36268 3664
rect 35667 3624 36268 3652
rect 35667 3621 35679 3624
rect 35621 3615 35679 3621
rect 36262 3612 36268 3624
rect 36320 3612 36326 3664
rect 21085 3587 21143 3593
rect 21085 3584 21097 3587
rect 20864 3556 21097 3584
rect 20864 3544 20870 3556
rect 21085 3553 21097 3556
rect 21131 3553 21143 3587
rect 21085 3547 21143 3553
rect 22373 3587 22431 3593
rect 22373 3553 22385 3587
rect 22419 3553 22431 3587
rect 22373 3547 22431 3553
rect 30193 3587 30251 3593
rect 30193 3553 30205 3587
rect 30239 3553 30251 3587
rect 30193 3547 30251 3553
rect 31110 3544 31116 3596
rect 31168 3584 31174 3596
rect 31389 3587 31447 3593
rect 31389 3584 31401 3587
rect 31168 3556 31401 3584
rect 31168 3544 31174 3556
rect 31389 3553 31401 3556
rect 31435 3584 31447 3587
rect 31570 3584 31576 3596
rect 31435 3556 31576 3584
rect 31435 3553 31447 3556
rect 31389 3547 31447 3553
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 32214 3584 32220 3596
rect 32175 3556 32220 3584
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 32585 3587 32643 3593
rect 32585 3553 32597 3587
rect 32631 3553 32643 3587
rect 32585 3547 32643 3553
rect 20622 3516 20628 3528
rect 19444 3488 20628 3516
rect 17589 3479 17647 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 24026 3516 24032 3528
rect 21499 3488 24032 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 24486 3516 24492 3528
rect 24447 3488 24492 3516
rect 24486 3476 24492 3488
rect 24544 3516 24550 3528
rect 24854 3516 24860 3528
rect 24544 3488 24860 3516
rect 24544 3476 24550 3488
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 26326 3476 26332 3528
rect 26384 3516 26390 3528
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 26384 3488 26709 3516
rect 26384 3476 26390 3488
rect 26697 3485 26709 3488
rect 26743 3516 26755 3519
rect 26786 3516 26792 3528
rect 26743 3488 26792 3516
rect 26743 3485 26755 3488
rect 26697 3479 26755 3485
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 28166 3516 28172 3528
rect 28127 3488 28172 3516
rect 28166 3476 28172 3488
rect 28224 3476 28230 3528
rect 31478 3476 31484 3528
rect 31536 3516 31542 3528
rect 31662 3516 31668 3528
rect 31536 3488 31668 3516
rect 31536 3476 31542 3488
rect 31662 3476 31668 3488
rect 31720 3516 31726 3528
rect 32600 3516 32628 3547
rect 33318 3544 33324 3596
rect 33376 3584 33382 3596
rect 33689 3587 33747 3593
rect 33689 3584 33701 3587
rect 33376 3556 33701 3584
rect 33376 3544 33382 3556
rect 33689 3553 33701 3556
rect 33735 3553 33747 3587
rect 33689 3547 33747 3553
rect 31720 3488 32628 3516
rect 32861 3519 32919 3525
rect 31720 3476 31726 3488
rect 32861 3485 32873 3519
rect 32907 3516 32919 3519
rect 35158 3516 35164 3528
rect 32907 3488 35164 3516
rect 32907 3485 32919 3488
rect 32861 3479 32919 3485
rect 35158 3476 35164 3488
rect 35216 3476 35222 3528
rect 35529 3519 35587 3525
rect 35529 3485 35541 3519
rect 35575 3516 35587 3519
rect 35894 3516 35900 3528
rect 35575 3488 35900 3516
rect 35575 3485 35587 3488
rect 35529 3479 35587 3485
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 36044 3488 36089 3516
rect 36044 3476 36050 3488
rect 7742 3408 7748 3460
rect 7800 3408 7806 3460
rect 13081 3451 13139 3457
rect 13081 3417 13093 3451
rect 13127 3448 13139 3451
rect 13906 3448 13912 3460
rect 13127 3420 13912 3448
rect 13127 3417 13139 3420
rect 13081 3411 13139 3417
rect 13906 3408 13912 3420
rect 13964 3448 13970 3460
rect 15933 3451 15991 3457
rect 15933 3448 15945 3451
rect 13964 3420 15945 3448
rect 13964 3408 13970 3420
rect 15933 3417 15945 3420
rect 15979 3448 15991 3451
rect 17497 3451 17555 3457
rect 17497 3448 17509 3451
rect 15979 3420 17509 3448
rect 15979 3417 15991 3420
rect 15933 3411 15991 3417
rect 17497 3417 17509 3420
rect 17543 3448 17555 3451
rect 18230 3448 18236 3460
rect 17543 3420 18236 3448
rect 17543 3417 17555 3420
rect 17497 3411 17555 3417
rect 18230 3408 18236 3420
rect 18288 3408 18294 3460
rect 2498 3380 2504 3392
rect 2459 3352 2504 3380
rect 2498 3340 2504 3352
rect 2556 3340 2562 3392
rect 7760 3380 7788 3408
rect 7929 3383 7987 3389
rect 7929 3380 7941 3383
rect 7760 3352 7941 3380
rect 7929 3349 7941 3352
rect 7975 3380 7987 3383
rect 8754 3380 8760 3392
rect 7975 3352 8760 3380
rect 7975 3349 7987 3352
rect 7929 3343 7987 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 12526 3380 12532 3392
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14553 3383 14611 3389
rect 14553 3380 14565 3383
rect 14056 3352 14565 3380
rect 14056 3340 14062 3352
rect 14553 3349 14565 3352
rect 14599 3349 14611 3383
rect 14553 3343 14611 3349
rect 15746 3340 15752 3392
rect 15804 3389 15810 3392
rect 15804 3383 15853 3389
rect 15804 3349 15807 3383
rect 15841 3349 15853 3383
rect 18598 3380 18604 3392
rect 18559 3352 18604 3380
rect 15804 3343 15853 3349
rect 15804 3340 15810 3343
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 21818 3380 21824 3392
rect 21779 3352 21824 3380
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 25498 3380 25504 3392
rect 25459 3352 25504 3380
rect 25498 3340 25504 3352
rect 25556 3340 25562 3392
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 29089 3383 29147 3389
rect 29089 3380 29101 3383
rect 28960 3352 29101 3380
rect 28960 3340 28966 3352
rect 29089 3349 29101 3352
rect 29135 3380 29147 3383
rect 29362 3380 29368 3392
rect 29135 3352 29368 3380
rect 29135 3349 29147 3352
rect 29089 3343 29147 3349
rect 29362 3340 29368 3352
rect 29420 3340 29426 3392
rect 29457 3383 29515 3389
rect 29457 3349 29469 3383
rect 29503 3380 29515 3383
rect 29546 3380 29552 3392
rect 29503 3352 29552 3380
rect 29503 3349 29515 3352
rect 29457 3343 29515 3349
rect 29546 3340 29552 3352
rect 29604 3340 29610 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 1762 3176 1768 3188
rect 1719 3148 1768 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 3694 3176 3700 3188
rect 3655 3148 3700 3176
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 4154 3176 4160 3188
rect 4111 3148 4160 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5442 3176 5448 3188
rect 5123 3148 5448 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 2777 3111 2835 3117
rect 2777 3077 2789 3111
rect 2823 3108 2835 3111
rect 2958 3108 2964 3120
rect 2823 3080 2964 3108
rect 2823 3077 2835 3080
rect 2777 3071 2835 3077
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1544 3012 2237 3040
rect 1544 3000 1550 3012
rect 2225 3009 2237 3012
rect 2271 3040 2283 3043
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2271 3012 3157 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 5092 2984 5120 3139
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 8110 3176 8116 3188
rect 8071 3148 8116 3176
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9548 3148 9873 3176
rect 9548 3136 9554 3148
rect 9861 3145 9873 3148
rect 9907 3176 9919 3179
rect 9950 3176 9956 3188
rect 9907 3148 9956 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10505 3179 10563 3185
rect 10505 3176 10517 3179
rect 10284 3148 10517 3176
rect 10284 3136 10290 3148
rect 10505 3145 10517 3148
rect 10551 3145 10563 3179
rect 12158 3176 12164 3188
rect 12119 3148 12164 3176
rect 10505 3139 10563 3145
rect 5258 3108 5264 3120
rect 5219 3080 5264 3108
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 6288 3040 6316 3136
rect 10520 3040 10548 3139
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 13320 3148 13461 3176
rect 13320 3136 13326 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 15102 3176 15108 3188
rect 13449 3139 13507 3145
rect 14108 3148 15108 3176
rect 12526 3108 12532 3120
rect 12439 3080 12532 3108
rect 12526 3068 12532 3080
rect 12584 3108 12590 3120
rect 14108 3117 14136 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 16298 3176 16304 3188
rect 15804 3148 16304 3176
rect 15804 3136 15810 3148
rect 16298 3136 16304 3148
rect 16356 3176 16362 3188
rect 16577 3179 16635 3185
rect 16577 3176 16589 3179
rect 16356 3148 16589 3176
rect 16356 3136 16362 3148
rect 16577 3145 16589 3148
rect 16623 3145 16635 3179
rect 16577 3139 16635 3145
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17221 3179 17279 3185
rect 17221 3176 17233 3179
rect 17184 3148 17233 3176
rect 17184 3136 17190 3148
rect 17221 3145 17233 3148
rect 17267 3145 17279 3179
rect 17221 3139 17279 3145
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17644 3148 17785 3176
rect 17644 3136 17650 3148
rect 17773 3145 17785 3148
rect 17819 3176 17831 3179
rect 17819 3148 18184 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 18156 3117 18184 3148
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 20901 3179 20959 3185
rect 20901 3176 20913 3179
rect 20864 3148 20913 3176
rect 20864 3136 20870 3148
rect 20901 3145 20913 3148
rect 20947 3145 20959 3179
rect 21266 3176 21272 3188
rect 21227 3148 21272 3176
rect 20901 3139 20959 3145
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21692 3148 21833 3176
rect 21692 3136 21698 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 23474 3176 23480 3188
rect 23435 3148 23480 3176
rect 21821 3139 21879 3145
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 24210 3176 24216 3188
rect 24171 3148 24216 3176
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 26053 3179 26111 3185
rect 26053 3145 26065 3179
rect 26099 3176 26111 3179
rect 26878 3176 26884 3188
rect 26099 3148 26884 3176
rect 26099 3145 26111 3148
rect 26053 3139 26111 3145
rect 26878 3136 26884 3148
rect 26936 3136 26942 3188
rect 28077 3179 28135 3185
rect 28077 3145 28089 3179
rect 28123 3176 28135 3179
rect 28166 3176 28172 3188
rect 28123 3148 28172 3176
rect 28123 3145 28135 3148
rect 28077 3139 28135 3145
rect 28166 3136 28172 3148
rect 28224 3136 28230 3188
rect 28718 3176 28724 3188
rect 28631 3148 28724 3176
rect 28718 3136 28724 3148
rect 28776 3176 28782 3188
rect 30285 3179 30343 3185
rect 30285 3176 30297 3179
rect 28776 3148 30297 3176
rect 28776 3136 28782 3148
rect 30285 3145 30297 3148
rect 30331 3176 30343 3179
rect 30466 3176 30472 3188
rect 30331 3148 30472 3176
rect 30331 3145 30343 3148
rect 30285 3139 30343 3145
rect 30466 3136 30472 3148
rect 30524 3136 30530 3188
rect 31941 3179 31999 3185
rect 31941 3145 31953 3179
rect 31987 3176 31999 3179
rect 32214 3176 32220 3188
rect 31987 3148 32220 3176
rect 31987 3145 31999 3148
rect 31941 3139 31999 3145
rect 32214 3136 32220 3148
rect 32272 3136 32278 3188
rect 33318 3136 33324 3188
rect 33376 3176 33382 3188
rect 34057 3179 34115 3185
rect 34057 3176 34069 3179
rect 33376 3148 34069 3176
rect 33376 3136 33382 3148
rect 34057 3145 34069 3148
rect 34103 3145 34115 3179
rect 34698 3176 34704 3188
rect 34659 3148 34704 3176
rect 34057 3139 34115 3145
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 35894 3176 35900 3188
rect 35855 3148 35900 3176
rect 35894 3136 35900 3148
rect 35952 3136 35958 3188
rect 36262 3176 36268 3188
rect 36223 3148 36268 3176
rect 36262 3136 36268 3148
rect 36320 3136 36326 3188
rect 37366 3136 37372 3188
rect 37424 3176 37430 3188
rect 37599 3179 37657 3185
rect 37599 3176 37611 3179
rect 37424 3148 37611 3176
rect 37424 3136 37430 3148
rect 37599 3145 37611 3148
rect 37645 3145 37657 3179
rect 37599 3139 37657 3145
rect 13909 3111 13967 3117
rect 13909 3108 13921 3111
rect 12584 3080 13921 3108
rect 12584 3068 12590 3080
rect 13909 3077 13921 3080
rect 13955 3108 13967 3111
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 13955 3080 14105 3108
rect 13955 3077 13967 3080
rect 13909 3071 13967 3077
rect 14093 3077 14105 3080
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 18141 3111 18199 3117
rect 18141 3077 18153 3111
rect 18187 3077 18199 3111
rect 18141 3071 18199 3077
rect 13078 3040 13084 3052
rect 6288 3012 7328 3040
rect 10520 3012 10824 3040
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4617 2975 4675 2981
rect 4617 2972 4629 2975
rect 4203 2944 4629 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4617 2941 4629 2944
rect 4663 2972 4675 2975
rect 4706 2972 4712 2984
rect 4663 2944 4712 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 5074 2972 5080 2984
rect 4987 2944 5080 2972
rect 5074 2932 5080 2944
rect 5132 2972 5138 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 5132 2944 5181 2972
rect 5132 2932 5138 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5442 2972 5448 2984
rect 5403 2944 5448 2972
rect 5169 2935 5227 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5810 2932 5816 2984
rect 5868 2972 5874 2984
rect 5994 2972 6000 2984
rect 5868 2944 6000 2972
rect 5868 2932 5874 2944
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6564 2944 6837 2972
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2904 2375 2907
rect 2498 2904 2504 2916
rect 2363 2876 2504 2904
rect 2363 2873 2375 2876
rect 2317 2867 2375 2873
rect 2038 2836 2044 2848
rect 1951 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2836 2102 2848
rect 2332 2836 2360 2867
rect 2498 2864 2504 2876
rect 2556 2864 2562 2916
rect 5902 2904 5908 2916
rect 5863 2876 5908 2904
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6564 2845 6592 2944
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 7098 2972 7104 2984
rect 6871 2944 7104 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7300 2981 7328 3012
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7926 2972 7932 2984
rect 7331 2944 7932 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8846 2972 8852 2984
rect 8527 2944 8852 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8846 2932 8852 2944
rect 8904 2972 8910 2984
rect 10796 2981 10824 3012
rect 12452 3012 12848 3040
rect 13039 3012 13084 3040
rect 12452 2981 12480 3012
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8904 2944 8953 2972
rect 8904 2932 8910 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 10689 2975 10747 2981
rect 10689 2972 10701 2975
rect 10275 2944 10701 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 10689 2941 10701 2944
rect 10735 2941 10747 2975
rect 10689 2935 10747 2941
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2941 10839 2975
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 10781 2935 10839 2941
rect 11808 2944 12449 2972
rect 8754 2904 8760 2916
rect 8667 2876 8760 2904
rect 8754 2864 8760 2876
rect 8812 2904 8818 2916
rect 9262 2907 9320 2913
rect 9262 2904 9274 2907
rect 8812 2876 9274 2904
rect 8812 2864 8818 2876
rect 9262 2873 9274 2876
rect 9308 2873 9320 2907
rect 10704 2904 10732 2935
rect 11606 2904 11612 2916
rect 10704 2876 11612 2904
rect 9262 2867 9320 2873
rect 11606 2864 11612 2876
rect 11664 2904 11670 2916
rect 11808 2913 11836 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12820 2972 12848 3012
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 16022 3040 16028 3052
rect 14016 3012 15608 3040
rect 15983 3012 16028 3040
rect 14016 2984 14044 3012
rect 13998 2972 14004 2984
rect 12820 2944 14004 2972
rect 12713 2935 12771 2941
rect 11793 2907 11851 2913
rect 11793 2904 11805 2907
rect 11664 2876 11805 2904
rect 11664 2864 11670 2876
rect 11793 2873 11805 2876
rect 11839 2873 11851 2907
rect 11793 2867 11851 2873
rect 12158 2864 12164 2916
rect 12216 2904 12222 2916
rect 12728 2904 12756 2935
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 15580 2981 15608 3012
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 18414 3000 18420 3052
rect 18472 3040 18478 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18472 3012 18521 3040
rect 18472 3000 18478 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 21652 3040 21680 3136
rect 27154 3108 27160 3120
rect 27115 3080 27160 3108
rect 27154 3068 27160 3080
rect 27212 3068 27218 3120
rect 33686 3108 33692 3120
rect 33647 3080 33692 3108
rect 33686 3068 33692 3080
rect 33744 3068 33750 3120
rect 22738 3040 22744 3052
rect 18509 3003 18567 3009
rect 19904 3012 21680 3040
rect 22699 3012 22744 3040
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 15565 2975 15623 2981
rect 15565 2941 15577 2975
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 15841 2975 15899 2981
rect 15712 2944 15757 2972
rect 15712 2932 15718 2944
rect 15841 2941 15853 2975
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 15381 2907 15439 2913
rect 15381 2904 15393 2907
rect 12216 2876 15393 2904
rect 12216 2864 12222 2876
rect 15381 2873 15393 2876
rect 15427 2904 15439 2907
rect 15856 2904 15884 2935
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 18012 2944 18061 2972
rect 18012 2932 18018 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 18049 2935 18107 2941
rect 18322 2932 18328 2944
rect 18380 2972 18386 2984
rect 18598 2972 18604 2984
rect 18380 2944 18604 2972
rect 18380 2932 18386 2944
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 19904 2981 19932 3012
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 19852 2944 19901 2972
rect 19852 2932 19858 2944
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2941 20131 2975
rect 21652 2972 21680 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3040 23811 3043
rect 26329 3043 26387 3049
rect 26329 3040 26341 3043
rect 23799 3012 26341 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 26329 3009 26341 3012
rect 26375 3040 26387 3043
rect 26605 3043 26663 3049
rect 26605 3040 26617 3043
rect 26375 3012 26617 3040
rect 26375 3009 26387 3012
rect 26329 3003 26387 3009
rect 26605 3009 26617 3012
rect 26651 3009 26663 3043
rect 26605 3003 26663 3009
rect 28307 3043 28365 3049
rect 28307 3009 28319 3043
rect 28353 3040 28365 3043
rect 29362 3040 29368 3052
rect 28353 3012 29368 3040
rect 28353 3009 28365 3012
rect 28307 3003 28365 3009
rect 29362 3000 29368 3012
rect 29420 3000 29426 3052
rect 29638 3040 29644 3052
rect 29599 3012 29644 3040
rect 29638 3000 29644 3012
rect 29696 3040 29702 3052
rect 30098 3040 30104 3052
rect 29696 3012 30104 3040
rect 29696 3000 29702 3012
rect 30098 3000 30104 3012
rect 30156 3000 30162 3052
rect 31573 3043 31631 3049
rect 31573 3009 31585 3043
rect 31619 3040 31631 3043
rect 31938 3040 31944 3052
rect 31619 3012 31944 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 31938 3000 31944 3012
rect 31996 3000 32002 3052
rect 33137 3043 33195 3049
rect 33137 3009 33149 3043
rect 33183 3040 33195 3043
rect 33962 3040 33968 3052
rect 33183 3012 33968 3040
rect 33183 3009 33195 3012
rect 33137 3003 33195 3009
rect 33962 3000 33968 3012
rect 34020 3000 34026 3052
rect 34974 3040 34980 3052
rect 34935 3012 34980 3040
rect 34974 3000 34980 3012
rect 35032 3000 35038 3052
rect 35066 3000 35072 3052
rect 35124 3040 35130 3052
rect 35253 3043 35311 3049
rect 35253 3040 35265 3043
rect 35124 3012 35265 3040
rect 35124 3000 35130 3012
rect 35253 3009 35265 3012
rect 35299 3009 35311 3043
rect 35912 3040 35940 3136
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 35912 3012 36461 3040
rect 35253 3003 35311 3009
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 22005 2975 22063 2981
rect 22005 2972 22017 2975
rect 21652 2944 22017 2972
rect 20073 2935 20131 2941
rect 22005 2941 22017 2944
rect 22051 2941 22063 2975
rect 22005 2935 22063 2941
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2972 22615 2975
rect 23382 2972 23388 2984
rect 22603 2944 23388 2972
rect 22603 2941 22615 2944
rect 22557 2935 22615 2941
rect 15427 2876 15884 2904
rect 15427 2873 15439 2876
rect 15381 2867 15439 2873
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 19153 2907 19211 2913
rect 19153 2904 19165 2907
rect 17828 2876 19165 2904
rect 17828 2864 17834 2876
rect 19153 2873 19165 2876
rect 19199 2904 19211 2907
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 19199 2876 19533 2904
rect 19199 2873 19211 2876
rect 19153 2867 19211 2873
rect 19521 2873 19533 2876
rect 19567 2904 19579 2907
rect 19610 2904 19616 2916
rect 19567 2876 19616 2904
rect 19567 2873 19579 2876
rect 19521 2867 19579 2873
rect 19610 2864 19616 2876
rect 19668 2904 19674 2916
rect 20088 2904 20116 2935
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 24762 2972 24768 2984
rect 24723 2944 24768 2972
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 28074 2932 28080 2984
rect 28132 2972 28138 2984
rect 28204 2975 28262 2981
rect 28204 2972 28216 2975
rect 28132 2944 28216 2972
rect 28132 2932 28138 2944
rect 28204 2941 28216 2944
rect 28250 2941 28262 2975
rect 30742 2972 30748 2984
rect 30655 2944 30748 2972
rect 28204 2935 28262 2941
rect 30742 2932 30748 2944
rect 30800 2972 30806 2984
rect 30837 2975 30895 2981
rect 30837 2972 30849 2975
rect 30800 2944 30849 2972
rect 30800 2932 30806 2944
rect 30837 2941 30849 2944
rect 30883 2941 30895 2975
rect 30837 2935 30895 2941
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 31389 2975 31447 2981
rect 31389 2972 31401 2975
rect 31352 2944 31401 2972
rect 31352 2932 31358 2944
rect 31389 2941 31401 2944
rect 31435 2972 31447 2975
rect 31478 2972 31484 2984
rect 31435 2944 31484 2972
rect 31435 2941 31447 2944
rect 31389 2935 31447 2941
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 32306 2972 32312 2984
rect 32219 2944 32312 2972
rect 32306 2932 32312 2944
rect 32364 2972 32370 2984
rect 32401 2975 32459 2981
rect 32401 2972 32413 2975
rect 32364 2944 32413 2972
rect 32364 2932 32370 2944
rect 32401 2941 32413 2944
rect 32447 2941 32459 2975
rect 32858 2972 32864 2984
rect 32819 2944 32864 2972
rect 32401 2935 32459 2941
rect 32858 2932 32864 2944
rect 32916 2932 32922 2984
rect 36998 2932 37004 2984
rect 37056 2972 37062 2984
rect 37496 2975 37554 2981
rect 37496 2972 37508 2975
rect 37056 2944 37508 2972
rect 37056 2932 37062 2944
rect 37496 2941 37508 2944
rect 37542 2972 37554 2975
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37542 2944 37933 2972
rect 37542 2941 37554 2944
rect 37496 2935 37554 2941
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 23106 2904 23112 2916
rect 19668 2876 20116 2904
rect 23019 2876 23112 2904
rect 19668 2864 19674 2876
rect 23106 2864 23112 2876
rect 23164 2904 23170 2916
rect 24673 2907 24731 2913
rect 24673 2904 24685 2907
rect 23164 2876 24685 2904
rect 23164 2864 23170 2876
rect 24673 2873 24685 2876
rect 24719 2904 24731 2907
rect 25038 2904 25044 2916
rect 24719 2876 25044 2904
rect 24719 2873 24731 2876
rect 24673 2867 24731 2873
rect 25038 2864 25044 2876
rect 25096 2913 25102 2916
rect 25096 2907 25144 2913
rect 25096 2873 25098 2907
rect 25132 2873 25144 2907
rect 26697 2907 26755 2913
rect 25096 2867 25144 2873
rect 25700 2876 26556 2904
rect 25096 2864 25102 2867
rect 2096 2808 2360 2836
rect 4341 2839 4399 2845
rect 2096 2796 2102 2808
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 4387 2808 6561 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 6914 2836 6920 2848
rect 6875 2808 6920 2836
rect 6549 2799 6607 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 13964 2808 14473 2836
rect 13964 2796 13970 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 15010 2836 15016 2848
rect 14971 2808 15016 2836
rect 14461 2799 14519 2805
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 19702 2836 19708 2848
rect 19663 2808 19708 2836
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 25700 2845 25728 2876
rect 25685 2839 25743 2845
rect 25685 2805 25697 2839
rect 25731 2805 25743 2839
rect 26528 2836 26556 2876
rect 26697 2873 26709 2907
rect 26743 2873 26755 2907
rect 26697 2867 26755 2873
rect 29089 2907 29147 2913
rect 29089 2873 29101 2907
rect 29135 2904 29147 2907
rect 29365 2907 29423 2913
rect 29365 2904 29377 2907
rect 29135 2876 29377 2904
rect 29135 2873 29147 2876
rect 29089 2867 29147 2873
rect 29365 2873 29377 2876
rect 29411 2873 29423 2907
rect 29365 2867 29423 2873
rect 26712 2836 26740 2867
rect 27525 2839 27583 2845
rect 27525 2836 27537 2839
rect 26528 2808 27537 2836
rect 25685 2799 25743 2805
rect 27525 2805 27537 2808
rect 27571 2805 27583 2839
rect 29380 2836 29408 2867
rect 29454 2864 29460 2916
rect 29512 2904 29518 2916
rect 29512 2876 29557 2904
rect 29512 2864 29518 2876
rect 34698 2864 34704 2916
rect 34756 2904 34762 2916
rect 35069 2907 35127 2913
rect 35069 2904 35081 2907
rect 34756 2876 35081 2904
rect 34756 2864 34762 2876
rect 35069 2873 35081 2876
rect 35115 2873 35127 2907
rect 35069 2867 35127 2873
rect 29730 2836 29736 2848
rect 29380 2808 29736 2836
rect 27525 2799 27583 2805
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 1670 2632 1676 2644
rect 1631 2604 1676 2632
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 2038 2632 2044 2644
rect 1999 2604 2044 2632
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 4764 2604 5365 2632
rect 4764 2592 4770 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 6052 2604 6285 2632
rect 6052 2592 6058 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 6273 2595 6331 2601
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 8018 2632 8024 2644
rect 7147 2604 8024 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8628 2604 9137 2632
rect 8628 2592 8634 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 9125 2595 9183 2601
rect 2056 2564 2084 2592
rect 2317 2567 2375 2573
rect 2317 2564 2329 2567
rect 2056 2536 2329 2564
rect 2317 2533 2329 2536
rect 2363 2533 2375 2567
rect 2317 2527 2375 2533
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 4062 2564 4068 2576
rect 2915 2536 4068 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 4433 2567 4491 2573
rect 4433 2533 4445 2567
rect 4479 2564 4491 2567
rect 7926 2564 7932 2576
rect 4479 2536 5212 2564
rect 7887 2536 7932 2564
rect 4479 2533 4491 2536
rect 4433 2527 4491 2533
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4724 2468 4905 2496
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 2004 2400 2237 2428
rect 2004 2388 2010 2400
rect 2225 2397 2237 2400
rect 2271 2428 2283 2431
rect 3145 2431 3203 2437
rect 3145 2428 3157 2431
rect 2271 2400 3157 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 3145 2397 3157 2400
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 4724 2301 4752 2468
rect 4893 2465 4905 2468
rect 4939 2496 4951 2499
rect 5074 2496 5080 2508
rect 4939 2468 5080 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5184 2505 5212 2536
rect 7926 2524 7932 2536
rect 7984 2564 7990 2576
rect 8846 2564 8852 2576
rect 7984 2536 8616 2564
rect 8807 2536 8852 2564
rect 7984 2524 7990 2536
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5350 2496 5356 2508
rect 5215 2468 5356 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5350 2456 5356 2468
rect 5408 2496 5414 2508
rect 5810 2496 5816 2508
rect 5408 2468 5816 2496
rect 5408 2456 5414 2468
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 6086 2496 6092 2508
rect 6043 2468 6092 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 6012 2428 6040 2459
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6914 2496 6920 2508
rect 6779 2468 6920 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 8588 2505 8616 2536
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7699 2468 8401 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8389 2465 8401 2468
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 5031 2400 6040 2428
rect 8404 2428 8432 2459
rect 8662 2428 8668 2440
rect 8404 2400 8668 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9140 2428 9168 2595
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 12710 2592 12716 2644
rect 12768 2592 12774 2644
rect 13262 2632 13268 2644
rect 13223 2604 13268 2632
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 16945 2635 17003 2641
rect 16632 2604 16677 2632
rect 16632 2592 16638 2604
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17310 2632 17316 2644
rect 16991 2604 17316 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 9950 2564 9956 2576
rect 9911 2536 9956 2564
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 10502 2564 10508 2576
rect 10463 2536 10508 2564
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11149 2567 11207 2573
rect 11149 2564 11161 2567
rect 11112 2536 11161 2564
rect 11112 2524 11118 2536
rect 11149 2533 11161 2536
rect 11195 2564 11207 2567
rect 12621 2567 12679 2573
rect 12621 2564 12633 2567
rect 11195 2536 12633 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 12621 2533 12633 2536
rect 12667 2564 12679 2567
rect 12728 2564 12756 2592
rect 12894 2564 12900 2576
rect 12667 2536 12900 2564
rect 12667 2533 12679 2536
rect 12621 2527 12679 2533
rect 12894 2524 12900 2536
rect 12952 2524 12958 2576
rect 10520 2496 10548 2524
rect 11368 2499 11426 2505
rect 11368 2496 11380 2499
rect 10520 2468 11380 2496
rect 11368 2465 11380 2468
rect 11414 2465 11426 2499
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 11368 2459 11426 2465
rect 12912 2468 13645 2496
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9140 2400 9873 2428
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11471 2431 11529 2437
rect 11471 2397 11483 2431
rect 11517 2428 11529 2431
rect 11882 2428 11888 2440
rect 11517 2400 11888 2428
rect 11517 2397 11529 2400
rect 11471 2391 11529 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12768 2431 12826 2437
rect 12768 2428 12780 2431
rect 12676 2400 12780 2428
rect 12676 2388 12682 2400
rect 12768 2397 12780 2400
rect 12814 2428 12826 2431
rect 12912 2428 12940 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 14148 2468 14197 2496
rect 14148 2456 14154 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 15212 2496 15240 2592
rect 17052 2505 17080 2604
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17494 2632 17500 2644
rect 17455 2604 17500 2632
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 17586 2592 17592 2644
rect 17644 2632 17650 2644
rect 18046 2632 18052 2644
rect 17644 2604 18052 2632
rect 17644 2592 17650 2604
rect 18046 2592 18052 2604
rect 18104 2632 18110 2644
rect 19705 2635 19763 2641
rect 18104 2604 18460 2632
rect 18104 2592 18110 2604
rect 18322 2564 18328 2576
rect 18283 2536 18328 2564
rect 18322 2524 18328 2536
rect 18380 2524 18386 2576
rect 18432 2505 18460 2604
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 19794 2632 19800 2644
rect 19751 2604 19800 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 20898 2632 20904 2644
rect 20859 2604 20904 2632
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 21358 2632 21364 2644
rect 21319 2604 21364 2632
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 23382 2632 23388 2644
rect 23343 2604 23388 2632
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 23566 2592 23572 2644
rect 23624 2632 23630 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 23624 2604 23765 2632
rect 23624 2592 23630 2604
rect 23753 2601 23765 2604
rect 23799 2601 23811 2635
rect 23753 2595 23811 2601
rect 24854 2592 24860 2644
rect 24912 2632 24918 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 24912 2604 25421 2632
rect 24912 2592 24918 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 26326 2632 26332 2644
rect 26287 2604 26332 2632
rect 25409 2595 25467 2601
rect 20622 2564 20628 2576
rect 20583 2536 20628 2564
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15212 2468 15577 2496
rect 14185 2459 14243 2465
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 19978 2496 19984 2508
rect 19935 2468 19984 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20916 2496 20944 2592
rect 23109 2567 23167 2573
rect 23109 2533 23121 2567
rect 23155 2564 23167 2567
rect 24762 2564 24768 2576
rect 23155 2536 24768 2564
rect 23155 2533 23167 2536
rect 23109 2527 23167 2533
rect 24762 2524 24768 2536
rect 24820 2564 24826 2576
rect 25041 2567 25099 2573
rect 25041 2564 25053 2567
rect 24820 2536 25053 2564
rect 24820 2524 24826 2536
rect 25041 2533 25053 2536
rect 25087 2533 25099 2567
rect 25041 2527 25099 2533
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20916 2468 21189 2496
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 22646 2496 22652 2508
rect 22607 2468 22652 2496
rect 21177 2459 21235 2465
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 22925 2499 22983 2505
rect 22925 2465 22937 2499
rect 22971 2465 22983 2499
rect 22925 2459 22983 2465
rect 12814 2400 12940 2428
rect 12989 2431 13047 2437
rect 12814 2397 12826 2400
rect 12768 2391 12826 2397
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 12989 2391 13047 2397
rect 15120 2400 15485 2428
rect 12069 2363 12127 2369
rect 12069 2329 12081 2363
rect 12115 2360 12127 2363
rect 13004 2360 13032 2391
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 12115 2332 14381 2360
rect 12115 2329 12127 2332
rect 12069 2323 12127 2329
rect 14369 2329 14381 2332
rect 14415 2360 14427 2363
rect 15010 2360 15016 2372
rect 14415 2332 15016 2360
rect 14415 2329 14427 2332
rect 14369 2323 14427 2329
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 3476 2264 4721 2292
rect 3476 2252 3482 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 12437 2295 12495 2301
rect 12437 2261 12449 2295
rect 12483 2292 12495 2295
rect 12802 2292 12808 2304
rect 12483 2264 12808 2292
rect 12483 2261 12495 2264
rect 12437 2255 12495 2261
rect 12802 2252 12808 2264
rect 12860 2292 12866 2304
rect 12897 2295 12955 2301
rect 12897 2292 12909 2295
rect 12860 2264 12909 2292
rect 12860 2252 12866 2264
rect 12897 2261 12909 2264
rect 12943 2261 12955 2295
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 12897 2255 12955 2261
rect 14826 2252 14832 2264
rect 14884 2292 14890 2304
rect 15120 2292 15148 2400
rect 15473 2397 15485 2400
rect 15519 2428 15531 2431
rect 15654 2428 15660 2440
rect 15519 2400 15660 2428
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 21729 2431 21787 2437
rect 21729 2397 21741 2431
rect 21775 2428 21787 2431
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21775 2400 22109 2428
rect 21775 2397 21787 2400
rect 21729 2391 21787 2397
rect 22097 2397 22109 2400
rect 22143 2428 22155 2431
rect 22940 2428 22968 2459
rect 23566 2456 23572 2508
rect 23624 2496 23630 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23624 2468 24041 2496
rect 23624 2456 23630 2468
rect 24029 2465 24041 2468
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 24489 2499 24547 2505
rect 24489 2465 24501 2499
rect 24535 2465 24547 2499
rect 25424 2496 25452 2595
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 27246 2632 27252 2644
rect 27207 2604 27252 2632
rect 27246 2592 27252 2604
rect 27304 2592 27310 2644
rect 28813 2635 28871 2641
rect 28813 2601 28825 2635
rect 28859 2632 28871 2635
rect 28902 2632 28908 2644
rect 28859 2604 28908 2632
rect 28859 2601 28871 2604
rect 28813 2595 28871 2601
rect 28902 2592 28908 2604
rect 28960 2592 28966 2644
rect 29454 2632 29460 2644
rect 29415 2604 29460 2632
rect 29454 2592 29460 2604
rect 29512 2592 29518 2644
rect 29914 2592 29920 2644
rect 29972 2632 29978 2644
rect 30929 2635 30987 2641
rect 30929 2632 30941 2635
rect 29972 2604 30941 2632
rect 29972 2592 29978 2604
rect 27264 2564 27292 2592
rect 28166 2564 28172 2576
rect 27264 2536 27936 2564
rect 28127 2536 28172 2564
rect 25628 2499 25686 2505
rect 25628 2496 25640 2499
rect 25424 2468 25640 2496
rect 24489 2459 24547 2465
rect 25628 2465 25640 2468
rect 25674 2465 25686 2499
rect 26694 2496 26700 2508
rect 26607 2468 26700 2496
rect 25628 2459 25686 2465
rect 23382 2428 23388 2440
rect 22143 2400 23388 2428
rect 22143 2397 22155 2400
rect 22097 2391 22155 2397
rect 23382 2388 23388 2400
rect 23440 2428 23446 2440
rect 24504 2428 24532 2459
rect 26694 2456 26700 2468
rect 26752 2496 26758 2508
rect 27706 2496 27712 2508
rect 26752 2468 27712 2496
rect 26752 2456 26758 2468
rect 27706 2456 27712 2468
rect 27764 2456 27770 2508
rect 27908 2505 27936 2536
rect 28166 2524 28172 2536
rect 28224 2524 28230 2576
rect 27893 2499 27951 2505
rect 27893 2465 27905 2499
rect 27939 2465 27951 2499
rect 29472 2496 29500 2592
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29472 2468 29745 2496
rect 27893 2459 27951 2465
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 29733 2459 29791 2465
rect 30024 2496 30052 2604
rect 30929 2601 30941 2604
rect 30975 2632 30987 2635
rect 31294 2632 31300 2644
rect 30975 2604 31300 2632
rect 30975 2601 30987 2604
rect 30929 2595 30987 2601
rect 31294 2592 31300 2604
rect 31352 2592 31358 2644
rect 31754 2592 31760 2644
rect 31812 2632 31818 2644
rect 32585 2635 32643 2641
rect 32585 2632 32597 2635
rect 31812 2604 32597 2632
rect 31812 2592 31818 2604
rect 32585 2601 32597 2604
rect 32631 2601 32643 2635
rect 32585 2595 32643 2601
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 33045 2635 33103 2641
rect 33045 2632 33057 2635
rect 32916 2604 33057 2632
rect 32916 2592 32922 2604
rect 33045 2601 33057 2604
rect 33091 2601 33103 2635
rect 34054 2632 34060 2644
rect 34015 2604 34060 2632
rect 33045 2595 33103 2601
rect 34054 2592 34060 2604
rect 34112 2592 34118 2644
rect 34974 2632 34980 2644
rect 34935 2604 34980 2632
rect 34974 2592 34980 2604
rect 35032 2592 35038 2644
rect 35986 2632 35992 2644
rect 35947 2604 35992 2632
rect 35986 2592 35992 2604
rect 36044 2592 36050 2644
rect 30098 2524 30104 2576
rect 30156 2564 30162 2576
rect 31312 2564 31340 2592
rect 32217 2567 32275 2573
rect 32217 2564 32229 2567
rect 30156 2536 30696 2564
rect 31312 2536 32229 2564
rect 30156 2524 30162 2536
rect 30193 2499 30251 2505
rect 30193 2496 30205 2499
rect 30024 2468 30205 2496
rect 24670 2428 24676 2440
rect 23440 2400 24532 2428
rect 24631 2400 24676 2428
rect 23440 2388 23446 2400
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 29181 2431 29239 2437
rect 29181 2397 29193 2431
rect 29227 2428 29239 2431
rect 30024 2428 30052 2468
rect 30193 2465 30205 2468
rect 30239 2465 30251 2499
rect 30668 2496 30696 2536
rect 32217 2533 32229 2536
rect 32263 2564 32275 2567
rect 32876 2564 32904 2592
rect 32263 2536 32904 2564
rect 32263 2533 32275 2536
rect 32217 2527 32275 2533
rect 31332 2499 31390 2505
rect 31332 2496 31344 2499
rect 30668 2468 31344 2496
rect 30193 2459 30251 2465
rect 31332 2465 31344 2468
rect 31378 2496 31390 2499
rect 31757 2499 31815 2505
rect 31757 2496 31769 2499
rect 31378 2468 31769 2496
rect 31378 2465 31390 2468
rect 31332 2459 31390 2465
rect 31757 2465 31769 2468
rect 31803 2465 31815 2499
rect 31757 2459 31815 2465
rect 33664 2499 33722 2505
rect 33664 2465 33676 2499
rect 33710 2496 33722 2499
rect 34072 2496 34100 2592
rect 33710 2468 34100 2496
rect 35504 2499 35562 2505
rect 33710 2465 33722 2468
rect 33664 2459 33722 2465
rect 35504 2465 35516 2499
rect 35550 2496 35562 2499
rect 36004 2496 36032 2592
rect 35550 2468 36032 2496
rect 35550 2465 35562 2468
rect 35504 2459 35562 2465
rect 36354 2456 36360 2508
rect 36412 2496 36418 2508
rect 36484 2499 36542 2505
rect 36484 2496 36496 2499
rect 36412 2468 36496 2496
rect 36412 2456 36418 2468
rect 36484 2465 36496 2468
rect 36530 2496 36542 2499
rect 36909 2499 36967 2505
rect 36909 2496 36921 2499
rect 36530 2468 36921 2496
rect 36530 2465 36542 2468
rect 36484 2459 36542 2465
rect 36909 2465 36921 2468
rect 36955 2465 36967 2499
rect 36909 2459 36967 2465
rect 30282 2428 30288 2440
rect 29227 2400 30052 2428
rect 30243 2400 30288 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36587 2431 36645 2437
rect 36587 2428 36599 2431
rect 35952 2400 36599 2428
rect 35952 2388 35958 2400
rect 36587 2397 36599 2400
rect 36633 2397 36645 2431
rect 36587 2391 36645 2397
rect 17221 2363 17279 2369
rect 17221 2329 17233 2363
rect 17267 2360 17279 2363
rect 17770 2360 17776 2372
rect 17267 2332 17776 2360
rect 17267 2329 17279 2332
rect 17221 2323 17279 2329
rect 17770 2320 17776 2332
rect 17828 2320 17834 2372
rect 35575 2363 35633 2369
rect 35575 2329 35587 2363
rect 35621 2360 35633 2363
rect 36354 2360 36360 2372
rect 35621 2332 36360 2360
rect 35621 2329 35633 2332
rect 35575 2323 35633 2329
rect 36354 2320 36360 2332
rect 36412 2320 36418 2372
rect 20070 2292 20076 2304
rect 14884 2264 15148 2292
rect 20031 2264 20076 2292
rect 14884 2252 14890 2264
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 25731 2295 25789 2301
rect 25731 2261 25743 2295
rect 25777 2292 25789 2295
rect 25958 2292 25964 2304
rect 25777 2264 25964 2292
rect 25777 2261 25789 2264
rect 25731 2255 25789 2261
rect 25958 2252 25964 2264
rect 26016 2252 26022 2304
rect 31435 2295 31493 2301
rect 31435 2261 31447 2295
rect 31481 2292 31493 2295
rect 31662 2292 31668 2304
rect 31481 2264 31668 2292
rect 31481 2261 31493 2264
rect 31435 2255 31493 2261
rect 31662 2252 31668 2264
rect 31720 2252 31726 2304
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 33735 2295 33793 2301
rect 33735 2292 33747 2295
rect 33192 2264 33747 2292
rect 33192 2252 33198 2264
rect 33735 2261 33747 2264
rect 33781 2261 33793 2295
rect 33735 2255 33793 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 22094 552 22100 604
rect 22152 592 22158 604
rect 22278 592 22284 604
rect 22152 564 22284 592
rect 22152 552 22158 564
rect 22278 552 22284 564
rect 22336 552 22342 604
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 35624 12971 35676 12980
rect 35624 12937 35633 12971
rect 35633 12937 35667 12971
rect 35667 12937 35676 12971
rect 35624 12928 35676 12937
rect 5448 12724 5500 12776
rect 35440 12767 35492 12776
rect 11336 12656 11388 12708
rect 1952 12588 2004 12640
rect 3700 12588 3752 12640
rect 5264 12588 5316 12640
rect 5448 12631 5500 12640
rect 5448 12597 5457 12631
rect 5457 12597 5491 12631
rect 5491 12597 5500 12631
rect 5448 12588 5500 12597
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 35440 12733 35449 12767
rect 35449 12733 35483 12767
rect 35483 12733 35492 12767
rect 35440 12724 35492 12733
rect 18420 12588 18472 12640
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 1492 12384 1544 12436
rect 1676 12248 1728 12300
rect 2872 12248 2924 12300
rect 3976 12248 4028 12300
rect 4252 12248 4304 12300
rect 5908 12291 5960 12300
rect 5908 12257 5952 12291
rect 5952 12257 5960 12291
rect 5908 12248 5960 12257
rect 10048 12248 10100 12300
rect 11336 12291 11388 12300
rect 11336 12257 11354 12291
rect 11354 12257 11388 12291
rect 11336 12248 11388 12257
rect 12164 12248 12216 12300
rect 13452 12248 13504 12300
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 2688 12044 2740 12053
rect 4160 12044 4212 12096
rect 6736 12044 6788 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 11796 12044 11848 12096
rect 14004 12044 14056 12096
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 14832 11704 14884 11756
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 2412 11679 2464 11688
rect 2412 11645 2421 11679
rect 2421 11645 2455 11679
rect 2455 11645 2464 11679
rect 2412 11636 2464 11645
rect 2596 11611 2648 11620
rect 2596 11577 2605 11611
rect 2605 11577 2639 11611
rect 2639 11577 2648 11611
rect 2596 11568 2648 11577
rect 4896 11679 4948 11688
rect 4896 11645 4940 11679
rect 4940 11645 4948 11679
rect 4896 11636 4948 11645
rect 7012 11636 7064 11688
rect 8116 11636 8168 11688
rect 10508 11636 10560 11688
rect 11244 11679 11296 11688
rect 11244 11645 11288 11679
rect 11288 11645 11296 11679
rect 11244 11636 11296 11645
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 4252 11568 4304 11620
rect 5448 11568 5500 11620
rect 10048 11568 10100 11620
rect 18328 11636 18380 11688
rect 19432 11636 19484 11688
rect 15016 11611 15068 11620
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 4988 11500 5040 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6920 11500 6972 11552
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 11428 11500 11480 11552
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 12716 11500 12768 11552
rect 13452 11500 13504 11552
rect 14004 11500 14056 11552
rect 15016 11577 15025 11611
rect 15025 11577 15059 11611
rect 15059 11577 15068 11611
rect 15016 11568 15068 11577
rect 18788 11500 18840 11552
rect 20076 11500 20128 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 17040 11296 17092 11348
rect 35624 11339 35676 11348
rect 35624 11305 35633 11339
rect 35633 11305 35667 11339
rect 35667 11305 35676 11339
rect 35624 11296 35676 11305
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 4252 11160 4304 11212
rect 5172 11203 5224 11212
rect 5172 11169 5190 11203
rect 5190 11169 5224 11203
rect 5172 11160 5224 11169
rect 6184 11203 6236 11212
rect 6184 11169 6202 11203
rect 6202 11169 6236 11203
rect 6184 11160 6236 11169
rect 7104 11203 7156 11212
rect 7104 11169 7148 11203
rect 7148 11169 7156 11203
rect 7104 11160 7156 11169
rect 8208 11203 8260 11212
rect 8208 11169 8226 11203
rect 8226 11169 8260 11203
rect 8208 11160 8260 11169
rect 9772 11160 9824 11212
rect 2228 11092 2280 11144
rect 9588 11092 9640 11144
rect 11704 11160 11756 11212
rect 1860 10956 1912 11008
rect 3516 10956 3568 11008
rect 4712 11024 4764 11076
rect 5448 11024 5500 11076
rect 6368 11024 6420 11076
rect 9864 11067 9916 11076
rect 9864 11033 9873 11067
rect 9873 11033 9907 11067
rect 9907 11033 9916 11067
rect 9864 11024 9916 11033
rect 10968 11024 11020 11076
rect 7472 10956 7524 11008
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 11244 10956 11296 11008
rect 13360 10956 13412 11008
rect 14004 11160 14056 11212
rect 16672 11160 16724 11212
rect 18512 11203 18564 11212
rect 18512 11169 18530 11203
rect 18530 11169 18564 11203
rect 18512 11160 18564 11169
rect 19524 11203 19576 11212
rect 19524 11169 19542 11203
rect 19542 11169 19576 11203
rect 19524 11160 19576 11169
rect 22100 11203 22152 11212
rect 22100 11169 22118 11203
rect 22118 11169 22152 11203
rect 22100 11160 22152 11169
rect 26608 11203 26660 11212
rect 26608 11169 26652 11203
rect 26652 11169 26660 11203
rect 26608 11160 26660 11169
rect 34152 11160 34204 11212
rect 35256 11160 35308 11212
rect 14924 11092 14976 11144
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 18604 11024 18656 11076
rect 19616 11024 19668 11076
rect 24308 11024 24360 11076
rect 27528 11024 27580 11076
rect 34060 10956 34112 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 1400 10752 1452 10804
rect 4068 10752 4120 10804
rect 6644 10752 6696 10804
rect 7104 10752 7156 10804
rect 8024 10752 8076 10804
rect 8300 10752 8352 10804
rect 9588 10752 9640 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 18512 10795 18564 10804
rect 18512 10761 18521 10795
rect 18521 10761 18555 10795
rect 18555 10761 18564 10795
rect 18512 10752 18564 10761
rect 26240 10795 26292 10804
rect 26240 10761 26249 10795
rect 26249 10761 26283 10795
rect 26283 10761 26292 10795
rect 26240 10752 26292 10761
rect 35624 10795 35676 10804
rect 35624 10761 35633 10795
rect 35633 10761 35667 10795
rect 35667 10761 35676 10795
rect 35624 10752 35676 10761
rect 2044 10684 2096 10736
rect 4068 10616 4120 10668
rect 4252 10616 4304 10668
rect 11520 10616 11572 10668
rect 14004 10616 14056 10668
rect 2504 10548 2556 10600
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 5172 10548 5224 10600
rect 5816 10591 5868 10600
rect 5816 10557 5834 10591
rect 5834 10557 5868 10591
rect 5816 10548 5868 10557
rect 10324 10591 10376 10600
rect 10324 10557 10368 10591
rect 10368 10557 10376 10591
rect 10324 10548 10376 10557
rect 11888 10548 11940 10600
rect 12992 10548 13044 10600
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 15292 10548 15344 10600
rect 16304 10591 16356 10600
rect 3976 10480 4028 10532
rect 8576 10480 8628 10532
rect 12072 10480 12124 10532
rect 15108 10480 15160 10532
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 18052 10591 18104 10600
rect 18052 10557 18096 10591
rect 18096 10557 18104 10591
rect 18052 10548 18104 10557
rect 18972 10548 19024 10600
rect 19984 10548 20036 10600
rect 20720 10548 20772 10600
rect 16488 10480 16540 10532
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 7288 10412 7340 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 9404 10412 9456 10464
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 10692 10412 10744 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 16212 10412 16264 10464
rect 16672 10412 16724 10464
rect 17868 10412 17920 10464
rect 19064 10412 19116 10464
rect 20720 10412 20772 10464
rect 22376 10548 22428 10600
rect 25688 10591 25740 10600
rect 25688 10557 25732 10591
rect 25732 10557 25740 10591
rect 25688 10548 25740 10557
rect 26148 10548 26200 10600
rect 26700 10591 26752 10600
rect 26700 10557 26744 10591
rect 26744 10557 26752 10591
rect 27160 10591 27212 10600
rect 26700 10548 26752 10557
rect 27160 10557 27169 10591
rect 27169 10557 27203 10591
rect 27203 10557 27212 10591
rect 27160 10548 27212 10557
rect 28172 10591 28224 10600
rect 28172 10557 28181 10591
rect 28181 10557 28215 10591
rect 28215 10557 28224 10591
rect 28172 10548 28224 10557
rect 21732 10480 21784 10532
rect 22100 10480 22152 10532
rect 27988 10480 28040 10532
rect 33416 10548 33468 10600
rect 35256 10591 35308 10600
rect 35256 10557 35265 10591
rect 35265 10557 35299 10591
rect 35299 10557 35308 10591
rect 35256 10548 35308 10557
rect 35440 10591 35492 10600
rect 35440 10557 35449 10591
rect 35449 10557 35483 10591
rect 35483 10557 35492 10591
rect 35440 10548 35492 10557
rect 21824 10412 21876 10464
rect 22008 10412 22060 10464
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 27252 10412 27304 10464
rect 33600 10412 33652 10464
rect 33784 10455 33836 10464
rect 33784 10421 33793 10455
rect 33793 10421 33827 10455
rect 33827 10421 33836 10455
rect 33784 10412 33836 10421
rect 34152 10412 34204 10464
rect 34796 10412 34848 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 3516 10251 3568 10260
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 6828 10208 6880 10260
rect 10784 10251 10836 10260
rect 10784 10217 10793 10251
rect 10793 10217 10827 10251
rect 10827 10217 10836 10251
rect 10784 10208 10836 10217
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 14004 10208 14056 10260
rect 27252 10208 27304 10260
rect 35716 10208 35768 10260
rect 2780 10140 2832 10192
rect 27436 10183 27488 10192
rect 27436 10149 27445 10183
rect 27445 10149 27479 10183
rect 27479 10149 27488 10183
rect 27436 10140 27488 10149
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 2320 10072 2372 10124
rect 3056 10115 3108 10124
rect 3056 10081 3074 10115
rect 3074 10081 3108 10115
rect 3056 10072 3108 10081
rect 4252 10115 4304 10124
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 5724 10115 5776 10124
rect 5724 10081 5742 10115
rect 5742 10081 5776 10115
rect 5724 10072 5776 10081
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 6920 10072 6972 10124
rect 9036 10072 9088 10124
rect 9772 10072 9824 10124
rect 11520 10072 11572 10124
rect 13728 10072 13780 10124
rect 15384 10072 15436 10124
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 19340 10115 19392 10124
rect 19340 10081 19384 10115
rect 19384 10081 19392 10115
rect 19340 10072 19392 10081
rect 4620 10047 4672 10056
rect 1860 9936 1912 9988
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 12440 10004 12492 10056
rect 12624 10004 12676 10056
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 20812 10004 20864 10056
rect 12808 9936 12860 9988
rect 20628 9936 20680 9988
rect 22928 10115 22980 10124
rect 21548 10004 21600 10056
rect 22928 10081 22937 10115
rect 22937 10081 22971 10115
rect 22971 10081 22980 10115
rect 22928 10072 22980 10081
rect 24124 10072 24176 10124
rect 25504 10115 25556 10124
rect 25504 10081 25522 10115
rect 25522 10081 25556 10115
rect 25504 10072 25556 10081
rect 28908 10115 28960 10124
rect 28908 10081 28926 10115
rect 28926 10081 28960 10115
rect 28908 10072 28960 10081
rect 33416 10115 33468 10124
rect 33416 10081 33460 10115
rect 33460 10081 33468 10115
rect 33416 10072 33468 10081
rect 34704 10072 34756 10124
rect 35808 10072 35860 10124
rect 36268 10072 36320 10124
rect 37188 10072 37240 10124
rect 22468 10004 22520 10056
rect 27528 10004 27580 10056
rect 29184 10004 29236 10056
rect 21640 9936 21692 9988
rect 2504 9868 2556 9920
rect 3240 9868 3292 9920
rect 5540 9868 5592 9920
rect 9588 9868 9640 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 13176 9868 13228 9920
rect 14096 9868 14148 9920
rect 19708 9868 19760 9920
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 21272 9868 21324 9920
rect 21456 9868 21508 9920
rect 23756 9868 23808 9920
rect 24492 9868 24544 9920
rect 24584 9911 24636 9920
rect 24584 9877 24593 9911
rect 24593 9877 24627 9911
rect 24627 9877 24636 9911
rect 24584 9868 24636 9877
rect 25964 9868 26016 9920
rect 28448 9868 28500 9920
rect 34152 9868 34204 9920
rect 35256 9868 35308 9920
rect 35348 9868 35400 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 3056 9664 3108 9716
rect 3332 9664 3384 9716
rect 2780 9596 2832 9648
rect 4528 9664 4580 9716
rect 6644 9664 6696 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 9772 9664 9824 9716
rect 11520 9707 11572 9716
rect 11520 9673 11529 9707
rect 11529 9673 11563 9707
rect 11563 9673 11572 9707
rect 11520 9664 11572 9673
rect 12808 9664 12860 9716
rect 13084 9664 13136 9716
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 6920 9596 6972 9648
rect 11796 9639 11848 9648
rect 3516 9528 3568 9580
rect 5816 9528 5868 9580
rect 7564 9528 7616 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 2412 9460 2464 9512
rect 5172 9460 5224 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 13728 9596 13780 9648
rect 15292 9596 15344 9648
rect 16304 9596 16356 9648
rect 17960 9664 18012 9716
rect 19340 9707 19392 9716
rect 19340 9673 19349 9707
rect 19349 9673 19383 9707
rect 19383 9673 19392 9707
rect 19340 9664 19392 9673
rect 20812 9664 20864 9716
rect 25504 9707 25556 9716
rect 25504 9673 25513 9707
rect 25513 9673 25547 9707
rect 25547 9673 25556 9707
rect 25504 9664 25556 9673
rect 33416 9707 33468 9716
rect 33416 9673 33425 9707
rect 33425 9673 33459 9707
rect 33459 9673 33468 9707
rect 33416 9664 33468 9673
rect 12808 9528 12860 9580
rect 13176 9528 13228 9580
rect 13912 9528 13964 9580
rect 15660 9528 15712 9580
rect 8668 9460 8720 9512
rect 10508 9503 10560 9512
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 10876 9460 10928 9512
rect 11520 9460 11572 9512
rect 14648 9460 14700 9512
rect 2044 9392 2096 9444
rect 3516 9392 3568 9444
rect 3700 9435 3752 9444
rect 3700 9401 3709 9435
rect 3709 9401 3743 9435
rect 3743 9401 3752 9435
rect 3700 9392 3752 9401
rect 6276 9392 6328 9444
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7012 9392 7064 9401
rect 12532 9392 12584 9444
rect 13544 9392 13596 9444
rect 16120 9435 16172 9444
rect 16120 9401 16129 9435
rect 16129 9401 16163 9435
rect 16163 9401 16172 9435
rect 16672 9435 16724 9444
rect 16120 9392 16172 9401
rect 16672 9401 16681 9435
rect 16681 9401 16715 9435
rect 16715 9401 16724 9435
rect 16672 9392 16724 9401
rect 7104 9324 7156 9376
rect 8300 9324 8352 9376
rect 9036 9324 9088 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11796 9324 11848 9376
rect 12808 9324 12860 9376
rect 13268 9324 13320 9376
rect 13820 9324 13872 9376
rect 17040 9324 17092 9376
rect 26608 9596 26660 9648
rect 28632 9596 28684 9648
rect 32312 9639 32364 9648
rect 32312 9605 32321 9639
rect 32321 9605 32355 9639
rect 32355 9605 32364 9639
rect 32312 9596 32364 9605
rect 35532 9639 35584 9648
rect 35532 9605 35541 9639
rect 35541 9605 35575 9639
rect 35575 9605 35584 9639
rect 35532 9596 35584 9605
rect 36636 9639 36688 9648
rect 36636 9605 36645 9639
rect 36645 9605 36679 9639
rect 36679 9605 36688 9639
rect 36636 9596 36688 9605
rect 20536 9528 20588 9580
rect 21916 9528 21968 9580
rect 24768 9571 24820 9580
rect 24768 9537 24777 9571
rect 24777 9537 24811 9571
rect 24811 9537 24820 9571
rect 24768 9528 24820 9537
rect 27252 9528 27304 9580
rect 17960 9460 18012 9512
rect 18512 9503 18564 9512
rect 18512 9469 18521 9503
rect 18521 9469 18555 9503
rect 18555 9469 18564 9503
rect 18512 9460 18564 9469
rect 19524 9460 19576 9512
rect 19892 9460 19944 9512
rect 22468 9503 22520 9512
rect 22468 9469 22477 9503
rect 22477 9469 22511 9503
rect 22511 9469 22520 9503
rect 22468 9460 22520 9469
rect 17684 9324 17736 9376
rect 18236 9392 18288 9444
rect 21456 9435 21508 9444
rect 21456 9401 21465 9435
rect 21465 9401 21499 9435
rect 21499 9401 21508 9435
rect 21456 9392 21508 9401
rect 21548 9435 21600 9444
rect 21548 9401 21557 9435
rect 21557 9401 21591 9435
rect 21591 9401 21600 9435
rect 21548 9392 21600 9401
rect 22100 9392 22152 9444
rect 22928 9435 22980 9444
rect 22928 9401 22937 9435
rect 22937 9401 22971 9435
rect 22971 9401 22980 9435
rect 22928 9392 22980 9401
rect 24032 9435 24084 9444
rect 24032 9401 24041 9435
rect 24041 9401 24075 9435
rect 24075 9401 24084 9435
rect 24492 9460 24544 9512
rect 26240 9460 26292 9512
rect 24032 9392 24084 9401
rect 24860 9392 24912 9444
rect 27436 9392 27488 9444
rect 28080 9435 28132 9444
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 26700 9324 26752 9376
rect 26884 9367 26936 9376
rect 26884 9333 26893 9367
rect 26893 9333 26927 9367
rect 26927 9333 26936 9367
rect 26884 9324 26936 9333
rect 28080 9401 28089 9435
rect 28089 9401 28123 9435
rect 28123 9401 28132 9435
rect 28080 9392 28132 9401
rect 30196 9460 30248 9512
rect 32588 9571 32640 9580
rect 32588 9537 32597 9571
rect 32597 9537 32631 9571
rect 32631 9537 32640 9571
rect 32588 9528 32640 9537
rect 35164 9571 35216 9580
rect 35164 9537 35173 9571
rect 35173 9537 35207 9571
rect 35207 9537 35216 9571
rect 35164 9528 35216 9537
rect 33692 9460 33744 9512
rect 36452 9503 36504 9512
rect 36452 9469 36461 9503
rect 36461 9469 36495 9503
rect 36495 9469 36504 9503
rect 36452 9460 36504 9469
rect 36084 9392 36136 9444
rect 28724 9324 28776 9376
rect 28908 9324 28960 9376
rect 29092 9324 29144 9376
rect 29828 9367 29880 9376
rect 29828 9333 29837 9367
rect 29837 9333 29871 9367
rect 29871 9333 29880 9367
rect 29828 9324 29880 9333
rect 30472 9367 30524 9376
rect 30472 9333 30481 9367
rect 30481 9333 30515 9367
rect 30515 9333 30524 9367
rect 30472 9324 30524 9333
rect 32680 9324 32732 9376
rect 33324 9324 33376 9376
rect 33508 9324 33560 9376
rect 34704 9367 34756 9376
rect 34704 9333 34713 9367
rect 34713 9333 34747 9367
rect 34747 9333 34756 9367
rect 34704 9324 34756 9333
rect 35164 9324 35216 9376
rect 35900 9367 35952 9376
rect 35900 9333 35909 9367
rect 35909 9333 35943 9367
rect 35943 9333 35952 9367
rect 35900 9324 35952 9333
rect 37280 9324 37332 9376
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 2504 9120 2556 9172
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 10600 9120 10652 9172
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 12624 9120 12676 9172
rect 13176 9120 13228 9172
rect 16120 9120 16172 9172
rect 17960 9120 18012 9172
rect 18696 9163 18748 9172
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 18696 9120 18748 9129
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 20628 9120 20680 9172
rect 21824 9120 21876 9172
rect 22192 9120 22244 9172
rect 23480 9120 23532 9172
rect 26700 9120 26752 9172
rect 28908 9120 28960 9172
rect 33600 9163 33652 9172
rect 33600 9129 33609 9163
rect 33609 9129 33643 9163
rect 33643 9129 33652 9163
rect 33600 9120 33652 9129
rect 2872 9052 2924 9104
rect 3700 9052 3752 9104
rect 4252 9095 4304 9104
rect 4252 9061 4261 9095
rect 4261 9061 4295 9095
rect 4295 9061 4304 9095
rect 4252 9052 4304 9061
rect 7380 9095 7432 9104
rect 7380 9061 7389 9095
rect 7389 9061 7423 9095
rect 7423 9061 7432 9095
rect 7380 9052 7432 9061
rect 11888 9052 11940 9104
rect 13452 9052 13504 9104
rect 15384 9052 15436 9104
rect 17224 9095 17276 9104
rect 17224 9061 17233 9095
rect 17233 9061 17267 9095
rect 17267 9061 17276 9095
rect 17224 9052 17276 9061
rect 18512 9095 18564 9104
rect 18512 9061 18521 9095
rect 18521 9061 18555 9095
rect 18555 9061 18564 9095
rect 21272 9095 21324 9104
rect 18512 9052 18564 9061
rect 1676 8984 1728 9036
rect 5632 9027 5684 9036
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 6276 8984 6328 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10140 8984 10192 9036
rect 10876 8984 10928 9036
rect 15200 8984 15252 9036
rect 18236 8984 18288 9036
rect 21272 9061 21281 9095
rect 21281 9061 21315 9095
rect 21315 9061 21324 9095
rect 21272 9052 21324 9061
rect 21364 9095 21416 9104
rect 21364 9061 21373 9095
rect 21373 9061 21407 9095
rect 21407 9061 21416 9095
rect 21364 9052 21416 9061
rect 24584 9052 24636 9104
rect 26976 9052 27028 9104
rect 27712 9052 27764 9104
rect 27988 9052 28040 9104
rect 29000 9095 29052 9104
rect 2688 8916 2740 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 5080 8916 5132 8968
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 19800 8984 19852 9036
rect 20812 8984 20864 9036
rect 22836 9027 22888 9036
rect 22836 8993 22854 9027
rect 22854 8993 22888 9027
rect 22836 8984 22888 8993
rect 23940 8984 23992 9036
rect 24860 9027 24912 9036
rect 4528 8848 4580 8900
rect 5448 8848 5500 8900
rect 6000 8848 6052 8900
rect 8392 8848 8444 8900
rect 8760 8848 8812 8900
rect 12256 8891 12308 8900
rect 12256 8857 12265 8891
rect 12265 8857 12299 8891
rect 12299 8857 12308 8891
rect 12256 8848 12308 8857
rect 16672 8848 16724 8900
rect 19248 8916 19300 8968
rect 19340 8916 19392 8968
rect 21824 8891 21876 8900
rect 21824 8857 21833 8891
rect 21833 8857 21867 8891
rect 21867 8857 21876 8891
rect 21824 8848 21876 8857
rect 24860 8993 24869 9027
rect 24869 8993 24903 9027
rect 24903 8993 24912 9027
rect 24860 8984 24912 8993
rect 24952 8984 25004 9036
rect 25412 8916 25464 8968
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 27620 8916 27672 8968
rect 28080 8916 28132 8968
rect 28540 8916 28592 8968
rect 29000 9061 29009 9095
rect 29009 9061 29043 9095
rect 29043 9061 29052 9095
rect 29000 9052 29052 9061
rect 34060 9095 34112 9104
rect 34060 9061 34069 9095
rect 34069 9061 34103 9095
rect 34103 9061 34112 9095
rect 34060 9052 34112 9061
rect 35624 9095 35676 9104
rect 35624 9061 35633 9095
rect 35633 9061 35667 9095
rect 35667 9061 35676 9095
rect 35624 9052 35676 9061
rect 30380 9027 30432 9036
rect 30380 8993 30424 9027
rect 30424 8993 30432 9027
rect 32312 9027 32364 9036
rect 30380 8984 30432 8993
rect 32312 8993 32321 9027
rect 32321 8993 32355 9027
rect 32355 8993 32364 9027
rect 32312 8984 32364 8993
rect 32772 8984 32824 9036
rect 29184 8959 29236 8968
rect 29184 8925 29193 8959
rect 29193 8925 29227 8959
rect 29227 8925 29236 8959
rect 29184 8916 29236 8925
rect 32956 8916 33008 8968
rect 33324 8916 33376 8968
rect 34152 8916 34204 8968
rect 29828 8848 29880 8900
rect 33876 8848 33928 8900
rect 34336 8916 34388 8968
rect 36268 8916 36320 8968
rect 36728 8848 36780 8900
rect 1492 8780 1544 8832
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 3516 8823 3568 8832
rect 3516 8789 3525 8823
rect 3525 8789 3559 8823
rect 3559 8789 3568 8823
rect 3516 8780 3568 8789
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 8852 8823 8904 8832
rect 8852 8789 8861 8823
rect 8861 8789 8895 8823
rect 8895 8789 8904 8823
rect 8852 8780 8904 8789
rect 19524 8780 19576 8832
rect 19800 8780 19852 8832
rect 21456 8780 21508 8832
rect 24124 8780 24176 8832
rect 27528 8780 27580 8832
rect 27620 8780 27672 8832
rect 28080 8780 28132 8832
rect 30564 8780 30616 8832
rect 31392 8780 31444 8832
rect 33324 8823 33376 8832
rect 33324 8789 33333 8823
rect 33333 8789 33367 8823
rect 33367 8789 33376 8823
rect 33324 8780 33376 8789
rect 34980 8823 35032 8832
rect 34980 8789 34989 8823
rect 34989 8789 35023 8823
rect 35023 8789 35032 8823
rect 34980 8780 35032 8789
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 3148 8576 3200 8628
rect 4252 8576 4304 8628
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 5632 8576 5684 8628
rect 7380 8576 7432 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 12624 8576 12676 8628
rect 12900 8576 12952 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 17132 8576 17184 8628
rect 18512 8576 18564 8628
rect 19248 8619 19300 8628
rect 19248 8585 19257 8619
rect 19257 8585 19291 8619
rect 19291 8585 19300 8619
rect 19248 8576 19300 8585
rect 21272 8576 21324 8628
rect 22836 8619 22888 8628
rect 22836 8585 22845 8619
rect 22845 8585 22879 8619
rect 22879 8585 22888 8619
rect 22836 8576 22888 8585
rect 23940 8619 23992 8628
rect 23940 8585 23949 8619
rect 23949 8585 23983 8619
rect 23983 8585 23992 8619
rect 23940 8576 23992 8585
rect 27804 8576 27856 8628
rect 29000 8576 29052 8628
rect 34060 8576 34112 8628
rect 35624 8576 35676 8628
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 36636 8619 36688 8628
rect 36636 8585 36645 8619
rect 36645 8585 36679 8619
rect 36679 8585 36688 8619
rect 36636 8576 36688 8585
rect 2412 8551 2464 8560
rect 2412 8517 2421 8551
rect 2421 8517 2455 8551
rect 2455 8517 2464 8551
rect 2412 8508 2464 8517
rect 3884 8508 3936 8560
rect 5816 8551 5868 8560
rect 1952 8440 2004 8492
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 5080 8440 5132 8492
rect 5816 8517 5825 8551
rect 5825 8517 5859 8551
rect 5859 8517 5868 8551
rect 5816 8508 5868 8517
rect 7288 8508 7340 8560
rect 6000 8440 6052 8492
rect 10048 8508 10100 8560
rect 12256 8508 12308 8560
rect 2872 8347 2924 8356
rect 2872 8313 2881 8347
rect 2881 8313 2915 8347
rect 2915 8313 2924 8347
rect 2872 8304 2924 8313
rect 3148 8347 3200 8356
rect 3148 8313 3157 8347
rect 3157 8313 3191 8347
rect 3191 8313 3200 8347
rect 3148 8304 3200 8313
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 8668 8372 8720 8424
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 11336 8440 11388 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13268 8508 13320 8560
rect 15384 8508 15436 8560
rect 16948 8508 17000 8560
rect 17960 8508 18012 8560
rect 18972 8508 19024 8560
rect 23572 8508 23624 8560
rect 29184 8508 29236 8560
rect 33876 8551 33928 8560
rect 13728 8440 13780 8492
rect 14648 8440 14700 8492
rect 14740 8372 14792 8424
rect 10968 8347 11020 8356
rect 10968 8313 10977 8347
rect 10977 8313 11011 8347
rect 11011 8313 11020 8347
rect 10968 8304 11020 8313
rect 11888 8347 11940 8356
rect 11888 8313 11897 8347
rect 11897 8313 11931 8347
rect 11931 8313 11940 8347
rect 11888 8304 11940 8313
rect 2780 8236 2832 8288
rect 3792 8236 3844 8288
rect 7288 8236 7340 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 14648 8304 14700 8356
rect 14924 8440 14976 8492
rect 19708 8440 19760 8492
rect 20076 8440 20128 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 29460 8440 29512 8492
rect 33876 8517 33885 8551
rect 33885 8517 33919 8551
rect 33919 8517 33928 8551
rect 35532 8551 35584 8560
rect 33876 8508 33928 8517
rect 35532 8517 35541 8551
rect 35541 8517 35575 8551
rect 35575 8517 35584 8551
rect 35532 8508 35584 8517
rect 33600 8440 33652 8492
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 16856 8372 16908 8424
rect 14924 8304 14976 8356
rect 15384 8304 15436 8356
rect 12900 8236 12952 8288
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 16488 8236 16540 8288
rect 17224 8304 17276 8356
rect 18512 8304 18564 8356
rect 19340 8304 19392 8356
rect 21272 8372 21324 8424
rect 24400 8415 24452 8424
rect 24400 8381 24409 8415
rect 24409 8381 24443 8415
rect 24443 8381 24452 8415
rect 24400 8372 24452 8381
rect 20720 8304 20772 8356
rect 21548 8347 21600 8356
rect 21548 8313 21557 8347
rect 21557 8313 21591 8347
rect 21591 8313 21600 8347
rect 21548 8304 21600 8313
rect 24952 8372 25004 8424
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 31392 8372 31444 8424
rect 25412 8347 25464 8356
rect 25412 8313 25421 8347
rect 25421 8313 25455 8347
rect 25455 8313 25464 8347
rect 25412 8304 25464 8313
rect 27804 8347 27856 8356
rect 27804 8313 27813 8347
rect 27813 8313 27847 8347
rect 27847 8313 27856 8347
rect 27804 8304 27856 8313
rect 27988 8304 28040 8356
rect 28540 8304 28592 8356
rect 26792 8236 26844 8288
rect 26976 8236 27028 8288
rect 30380 8347 30432 8356
rect 30380 8313 30389 8347
rect 30389 8313 30423 8347
rect 30423 8313 30432 8347
rect 30380 8304 30432 8313
rect 32312 8304 32364 8356
rect 32772 8347 32824 8356
rect 32772 8313 32781 8347
rect 32781 8313 32815 8347
rect 32815 8313 32824 8347
rect 32772 8304 32824 8313
rect 36268 8372 36320 8424
rect 33324 8304 33376 8356
rect 34612 8304 34664 8356
rect 32220 8236 32272 8288
rect 33968 8236 34020 8288
rect 38016 8415 38068 8424
rect 38016 8381 38025 8415
rect 38025 8381 38059 8415
rect 38059 8381 38068 8415
rect 38016 8372 38068 8381
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 2688 8032 2740 8084
rect 3148 8032 3200 8084
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 2504 8007 2556 8016
rect 2504 7973 2507 8007
rect 2507 7973 2541 8007
rect 2541 7973 2556 8007
rect 2504 7964 2556 7973
rect 4160 8007 4212 8016
rect 4160 7973 4169 8007
rect 4169 7973 4203 8007
rect 4203 7973 4212 8007
rect 4160 7964 4212 7973
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 5080 7964 5132 8016
rect 2228 7896 2280 7948
rect 5448 7896 5500 7948
rect 6460 7896 6512 7948
rect 6828 8032 6880 8084
rect 6920 8032 6972 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 8944 8032 8996 8084
rect 10600 8032 10652 8084
rect 10968 8032 11020 8084
rect 12348 8032 12400 8084
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 15384 8032 15436 8084
rect 7288 7964 7340 8016
rect 8392 7896 8444 7948
rect 9956 7939 10008 7948
rect 9956 7905 10000 7939
rect 10000 7905 10008 7939
rect 11980 7964 12032 8016
rect 12900 8007 12952 8016
rect 12900 7973 12909 8007
rect 12909 7973 12943 8007
rect 12943 7973 12952 8007
rect 12900 7964 12952 7973
rect 16488 8032 16540 8084
rect 19708 8032 19760 8084
rect 22008 8032 22060 8084
rect 23664 8075 23716 8084
rect 23664 8041 23673 8075
rect 23673 8041 23707 8075
rect 23707 8041 23716 8075
rect 23664 8032 23716 8041
rect 25872 8075 25924 8084
rect 25872 8041 25881 8075
rect 25881 8041 25915 8075
rect 25915 8041 25924 8075
rect 25872 8032 25924 8041
rect 27436 8075 27488 8084
rect 27436 8041 27445 8075
rect 27445 8041 27479 8075
rect 27479 8041 27488 8075
rect 27436 8032 27488 8041
rect 27988 8032 28040 8084
rect 28080 8075 28132 8084
rect 28080 8041 28089 8075
rect 28089 8041 28123 8075
rect 28123 8041 28132 8075
rect 28080 8032 28132 8041
rect 33508 8032 33560 8084
rect 34152 8032 34204 8084
rect 35532 8032 35584 8084
rect 36636 8075 36688 8084
rect 36636 8041 36645 8075
rect 36645 8041 36679 8075
rect 36679 8041 36688 8075
rect 36636 8032 36688 8041
rect 17132 7964 17184 8016
rect 17960 7964 18012 8016
rect 19156 7964 19208 8016
rect 21272 8007 21324 8016
rect 21272 7973 21281 8007
rect 21281 7973 21315 8007
rect 21315 7973 21324 8007
rect 21272 7964 21324 7973
rect 21824 8007 21876 8016
rect 21824 7973 21833 8007
rect 21833 7973 21867 8007
rect 21867 7973 21876 8007
rect 21824 7964 21876 7973
rect 22836 8007 22888 8016
rect 22836 7973 22845 8007
rect 22845 7973 22879 8007
rect 22879 7973 22888 8007
rect 22836 7964 22888 7973
rect 26792 7964 26844 8016
rect 28632 8007 28684 8016
rect 28632 7973 28641 8007
rect 28641 7973 28675 8007
rect 28675 7973 28684 8007
rect 28632 7964 28684 7973
rect 32220 7964 32272 8016
rect 34060 7964 34112 8016
rect 34704 7964 34756 8016
rect 9956 7896 10008 7905
rect 15200 7896 15252 7948
rect 18696 7896 18748 7948
rect 20720 7896 20772 7948
rect 24860 7939 24912 7948
rect 24860 7905 24869 7939
rect 24869 7905 24903 7939
rect 24903 7905 24912 7939
rect 24860 7896 24912 7905
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 30748 7939 30800 7948
rect 30748 7905 30757 7939
rect 30757 7905 30791 7939
rect 30791 7905 30800 7939
rect 30748 7896 30800 7905
rect 31300 7896 31352 7948
rect 33048 7939 33100 7948
rect 33048 7905 33057 7939
rect 33057 7905 33091 7939
rect 33091 7905 33100 7939
rect 33048 7896 33100 7905
rect 33876 7939 33928 7948
rect 33876 7905 33920 7939
rect 33920 7905 33928 7939
rect 36452 7939 36504 7948
rect 33876 7896 33928 7905
rect 36452 7905 36461 7939
rect 36461 7905 36495 7939
rect 36495 7905 36504 7939
rect 36452 7896 36504 7905
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 11704 7828 11756 7880
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 13544 7828 13596 7880
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 17500 7828 17552 7880
rect 17868 7828 17920 7880
rect 572 7760 624 7812
rect 21640 7828 21692 7880
rect 22468 7828 22520 7880
rect 24032 7828 24084 7880
rect 24952 7828 25004 7880
rect 27620 7828 27672 7880
rect 28540 7871 28592 7880
rect 28540 7837 28549 7871
rect 28549 7837 28583 7871
rect 28583 7837 28592 7871
rect 28540 7828 28592 7837
rect 29644 7828 29696 7880
rect 32128 7871 32180 7880
rect 32128 7837 32137 7871
rect 32137 7837 32171 7871
rect 32171 7837 32180 7871
rect 32128 7828 32180 7837
rect 35624 7871 35676 7880
rect 34796 7803 34848 7812
rect 34796 7769 34805 7803
rect 34805 7769 34839 7803
rect 34839 7769 34848 7803
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 35624 7828 35676 7837
rect 34796 7760 34848 7769
rect 36728 7760 36780 7812
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 5356 7692 5408 7744
rect 8668 7735 8720 7744
rect 8668 7701 8677 7735
rect 8677 7701 8711 7735
rect 8711 7701 8720 7735
rect 8668 7692 8720 7701
rect 16856 7735 16908 7744
rect 16856 7701 16865 7735
rect 16865 7701 16899 7735
rect 16899 7701 16908 7735
rect 16856 7692 16908 7701
rect 18512 7692 18564 7744
rect 18880 7692 18932 7744
rect 23572 7692 23624 7744
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 29460 7735 29512 7744
rect 29460 7701 29469 7735
rect 29469 7701 29503 7735
rect 29503 7701 29512 7735
rect 29460 7692 29512 7701
rect 34152 7692 34204 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 3516 7488 3568 7540
rect 4252 7488 4304 7540
rect 6460 7488 6512 7540
rect 6920 7488 6972 7540
rect 12808 7488 12860 7540
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 19248 7488 19300 7540
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 26976 7531 27028 7540
rect 26976 7497 26985 7531
rect 26985 7497 27019 7531
rect 27019 7497 27028 7531
rect 26976 7488 27028 7497
rect 27620 7531 27672 7540
rect 27620 7497 27629 7531
rect 27629 7497 27663 7531
rect 27663 7497 27672 7531
rect 27620 7488 27672 7497
rect 28632 7531 28684 7540
rect 28632 7497 28641 7531
rect 28641 7497 28675 7531
rect 28675 7497 28684 7531
rect 28632 7488 28684 7497
rect 32128 7488 32180 7540
rect 33048 7531 33100 7540
rect 33048 7497 33057 7531
rect 33057 7497 33091 7531
rect 33091 7497 33100 7531
rect 33048 7488 33100 7497
rect 33876 7488 33928 7540
rect 36452 7488 36504 7540
rect 2320 7420 2372 7472
rect 4344 7420 4396 7472
rect 7196 7420 7248 7472
rect 4620 7352 4672 7404
rect 4988 7352 5040 7404
rect 5540 7352 5592 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 6828 7395 6880 7404
rect 5632 7352 5684 7361
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 1676 7284 1728 7336
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 12900 7420 12952 7472
rect 21916 7420 21968 7472
rect 22468 7420 22520 7472
rect 23664 7420 23716 7472
rect 27528 7420 27580 7472
rect 10508 7352 10560 7404
rect 8760 7284 8812 7336
rect 8852 7284 8904 7336
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 15292 7352 15344 7404
rect 16488 7352 16540 7404
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 18144 7352 18196 7404
rect 19892 7352 19944 7404
rect 22008 7352 22060 7404
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 24492 7352 24544 7404
rect 25596 7352 25648 7404
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 29184 7352 29236 7404
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 33508 7352 33560 7404
rect 34796 7352 34848 7404
rect 35532 7420 35584 7472
rect 35624 7395 35676 7404
rect 35624 7361 35633 7395
rect 35633 7361 35667 7395
rect 35667 7361 35676 7395
rect 35624 7352 35676 7361
rect 36544 7395 36596 7404
rect 36544 7361 36553 7395
rect 36553 7361 36587 7395
rect 36587 7361 36596 7395
rect 36544 7352 36596 7361
rect 36728 7352 36780 7404
rect 28264 7327 28316 7336
rect 28264 7293 28273 7327
rect 28273 7293 28307 7327
rect 28307 7293 28316 7327
rect 28264 7284 28316 7293
rect 31300 7327 31352 7336
rect 2504 7216 2556 7268
rect 5356 7259 5408 7268
rect 5356 7225 5365 7259
rect 5365 7225 5399 7259
rect 5399 7225 5408 7259
rect 5356 7216 5408 7225
rect 7288 7216 7340 7268
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 8484 7148 8536 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 11980 7148 12032 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 15292 7216 15344 7268
rect 16120 7259 16172 7268
rect 16120 7225 16129 7259
rect 16129 7225 16163 7259
rect 16163 7225 16172 7259
rect 17868 7259 17920 7268
rect 16120 7216 16172 7225
rect 17868 7225 17877 7259
rect 17877 7225 17911 7259
rect 17911 7225 17920 7259
rect 17868 7216 17920 7225
rect 14740 7148 14792 7200
rect 17132 7191 17184 7200
rect 17132 7157 17141 7191
rect 17141 7157 17175 7191
rect 17175 7157 17184 7191
rect 17132 7148 17184 7157
rect 19156 7148 19208 7200
rect 20628 7216 20680 7268
rect 22468 7259 22520 7268
rect 22468 7225 22477 7259
rect 22477 7225 22511 7259
rect 22511 7225 22520 7259
rect 22468 7216 22520 7225
rect 24860 7259 24912 7268
rect 22836 7191 22888 7200
rect 22836 7157 22845 7191
rect 22845 7157 22879 7191
rect 22879 7157 22888 7191
rect 22836 7148 22888 7157
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 24860 7225 24869 7259
rect 24869 7225 24903 7259
rect 24903 7225 24912 7259
rect 24860 7216 24912 7225
rect 25964 7259 26016 7268
rect 25964 7225 25973 7259
rect 25973 7225 26007 7259
rect 26007 7225 26016 7259
rect 25964 7216 26016 7225
rect 26792 7216 26844 7268
rect 25320 7191 25372 7200
rect 23480 7148 23532 7157
rect 25320 7157 25329 7191
rect 25329 7157 25363 7191
rect 25363 7157 25372 7191
rect 25320 7148 25372 7157
rect 29460 7259 29512 7268
rect 29460 7225 29469 7259
rect 29469 7225 29503 7259
rect 29503 7225 29512 7259
rect 29460 7216 29512 7225
rect 29828 7216 29880 7268
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 33048 7216 33100 7268
rect 27528 7148 27580 7200
rect 30748 7148 30800 7200
rect 32220 7191 32272 7200
rect 32220 7157 32229 7191
rect 32229 7157 32263 7191
rect 32263 7157 32272 7191
rect 32220 7148 32272 7157
rect 34704 7191 34756 7200
rect 34704 7157 34713 7191
rect 34713 7157 34747 7191
rect 34747 7157 34756 7191
rect 34704 7148 34756 7157
rect 34796 7148 34848 7200
rect 35900 7191 35952 7200
rect 35900 7157 35909 7191
rect 35909 7157 35943 7191
rect 35943 7157 35952 7191
rect 35900 7148 35952 7157
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 4160 6944 4212 6996
rect 10508 6944 10560 6996
rect 11980 6944 12032 6996
rect 14096 6944 14148 6996
rect 14740 6944 14792 6996
rect 15200 6944 15252 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 18696 6944 18748 6996
rect 19892 6944 19944 6996
rect 20812 6944 20864 6996
rect 21916 6944 21968 6996
rect 22468 6944 22520 6996
rect 26056 6987 26108 6996
rect 26056 6953 26065 6987
rect 26065 6953 26099 6987
rect 26099 6953 26108 6987
rect 26056 6944 26108 6953
rect 28540 6944 28592 6996
rect 28632 6944 28684 6996
rect 29184 6944 29236 6996
rect 29460 6944 29512 6996
rect 36544 6944 36596 6996
rect 2504 6876 2556 6928
rect 4712 6876 4764 6928
rect 6276 6876 6328 6928
rect 8024 6876 8076 6928
rect 12900 6876 12952 6928
rect 16948 6876 17000 6928
rect 17868 6876 17920 6928
rect 18880 6919 18932 6928
rect 18880 6885 18889 6919
rect 18889 6885 18923 6919
rect 18923 6885 18932 6919
rect 18880 6876 18932 6885
rect 20628 6876 20680 6928
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 2872 6808 2924 6860
rect 5356 6808 5408 6860
rect 9588 6808 9640 6860
rect 10784 6808 10836 6860
rect 11888 6808 11940 6860
rect 15752 6808 15804 6860
rect 16396 6808 16448 6860
rect 20076 6808 20128 6860
rect 21272 6808 21324 6860
rect 22008 6808 22060 6860
rect 22928 6808 22980 6860
rect 23480 6876 23532 6928
rect 34152 6919 34204 6928
rect 24676 6808 24728 6860
rect 24952 6851 25004 6860
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 26792 6851 26844 6860
rect 26792 6817 26836 6851
rect 26836 6817 26844 6851
rect 26792 6808 26844 6817
rect 27436 6808 27488 6860
rect 27528 6808 27580 6860
rect 28080 6808 28132 6860
rect 30380 6808 30432 6860
rect 30472 6808 30524 6860
rect 31576 6808 31628 6860
rect 32128 6851 32180 6860
rect 32128 6817 32137 6851
rect 32137 6817 32171 6851
rect 32171 6817 32180 6851
rect 32128 6808 32180 6817
rect 1952 6740 2004 6792
rect 2596 6740 2648 6792
rect 3056 6740 3108 6792
rect 4804 6740 4856 6792
rect 5540 6740 5592 6792
rect 6368 6740 6420 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 6920 6740 6972 6792
rect 7472 6740 7524 6792
rect 5632 6672 5684 6724
rect 12716 6740 12768 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 16212 6740 16264 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 22376 6740 22428 6792
rect 27804 6783 27856 6792
rect 8208 6672 8260 6724
rect 18604 6672 18656 6724
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 8116 6604 8168 6656
rect 8852 6647 8904 6656
rect 8852 6613 8861 6647
rect 8861 6613 8895 6647
rect 8895 6613 8904 6647
rect 8852 6604 8904 6613
rect 9772 6604 9824 6656
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 17132 6604 17184 6656
rect 17868 6604 17920 6656
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 27804 6749 27813 6783
rect 27813 6749 27847 6783
rect 27847 6749 27856 6783
rect 27804 6740 27856 6749
rect 29552 6783 29604 6792
rect 29552 6749 29561 6783
rect 29561 6749 29595 6783
rect 29595 6749 29604 6783
rect 29552 6740 29604 6749
rect 32772 6808 32824 6860
rect 34152 6885 34155 6919
rect 34155 6885 34189 6919
rect 34189 6885 34204 6919
rect 34152 6876 34204 6885
rect 34704 6876 34756 6928
rect 35900 6919 35952 6928
rect 33692 6808 33744 6860
rect 35348 6851 35400 6860
rect 35348 6817 35357 6851
rect 35357 6817 35391 6851
rect 35391 6817 35400 6851
rect 35348 6808 35400 6817
rect 35900 6885 35903 6919
rect 35903 6885 35937 6919
rect 35937 6885 35952 6919
rect 35900 6876 35952 6885
rect 23848 6604 23900 6613
rect 27068 6604 27120 6656
rect 30932 6604 30984 6656
rect 31300 6604 31352 6656
rect 35440 6740 35492 6792
rect 34612 6672 34664 6724
rect 35808 6672 35860 6724
rect 33324 6647 33376 6656
rect 33324 6613 33333 6647
rect 33333 6613 33367 6647
rect 33367 6613 33376 6647
rect 33324 6604 33376 6613
rect 34796 6604 34848 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 2596 6400 2648 6452
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 5448 6400 5500 6452
rect 6368 6400 6420 6452
rect 8760 6400 8812 6452
rect 9588 6443 9640 6452
rect 4620 6332 4672 6384
rect 6276 6332 6328 6384
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 6552 6264 6604 6316
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 7012 6196 7064 6248
rect 9588 6409 9597 6443
rect 9597 6409 9631 6443
rect 9631 6409 9640 6443
rect 9588 6400 9640 6409
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 11980 6400 12032 6452
rect 12624 6400 12676 6452
rect 12808 6400 12860 6452
rect 12900 6400 12952 6452
rect 16212 6400 16264 6452
rect 18880 6400 18932 6452
rect 19616 6400 19668 6452
rect 21272 6443 21324 6452
rect 11704 6332 11756 6384
rect 13176 6332 13228 6384
rect 18788 6332 18840 6384
rect 12532 6307 12584 6316
rect 12532 6273 12541 6307
rect 12541 6273 12575 6307
rect 12575 6273 12584 6307
rect 12532 6264 12584 6273
rect 12624 6264 12676 6316
rect 10140 6239 10192 6248
rect 10140 6205 10149 6239
rect 10149 6205 10183 6239
rect 10183 6205 10192 6239
rect 10140 6196 10192 6205
rect 16396 6264 16448 6316
rect 21272 6409 21281 6443
rect 21281 6409 21315 6443
rect 21315 6409 21324 6443
rect 21272 6400 21324 6409
rect 28080 6443 28132 6452
rect 28080 6409 28089 6443
rect 28089 6409 28123 6443
rect 28123 6409 28132 6443
rect 28080 6400 28132 6409
rect 30840 6400 30892 6452
rect 32128 6443 32180 6452
rect 20076 6375 20128 6384
rect 20076 6341 20085 6375
rect 20085 6341 20119 6375
rect 20119 6341 20128 6375
rect 20076 6332 20128 6341
rect 21824 6332 21876 6384
rect 26792 6375 26844 6384
rect 26792 6341 26801 6375
rect 26801 6341 26835 6375
rect 26835 6341 26844 6375
rect 26792 6332 26844 6341
rect 27436 6332 27488 6384
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 22928 6307 22980 6316
rect 22928 6273 22937 6307
rect 22937 6273 22971 6307
rect 22971 6273 22980 6307
rect 22928 6264 22980 6273
rect 24676 6264 24728 6316
rect 24860 6264 24912 6316
rect 25228 6307 25280 6316
rect 25228 6273 25237 6307
rect 25237 6273 25271 6307
rect 25271 6273 25280 6307
rect 25228 6264 25280 6273
rect 27252 6264 27304 6316
rect 29000 6307 29052 6316
rect 29000 6273 29009 6307
rect 29009 6273 29043 6307
rect 29043 6273 29052 6307
rect 29000 6264 29052 6273
rect 2136 6128 2188 6180
rect 4160 6128 4212 6180
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 6276 6128 6328 6180
rect 8024 6128 8076 6180
rect 8300 6171 8352 6180
rect 8300 6137 8309 6171
rect 8309 6137 8343 6171
rect 8343 6137 8352 6171
rect 8300 6128 8352 6137
rect 10048 6128 10100 6180
rect 12348 6128 12400 6180
rect 14004 6171 14056 6180
rect 3148 6060 3200 6112
rect 3884 6060 3936 6112
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 6920 6060 6972 6112
rect 9680 6060 9732 6112
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 14004 6137 14013 6171
rect 14013 6137 14047 6171
rect 14047 6137 14056 6171
rect 14004 6128 14056 6137
rect 16948 6128 17000 6180
rect 17868 6171 17920 6180
rect 17868 6137 17877 6171
rect 17877 6137 17911 6171
rect 17911 6137 17920 6171
rect 18788 6171 18840 6180
rect 17868 6128 17920 6137
rect 12164 6060 12216 6069
rect 15752 6060 15804 6112
rect 18788 6137 18797 6171
rect 18797 6137 18831 6171
rect 18831 6137 18840 6171
rect 18788 6128 18840 6137
rect 19432 6171 19484 6180
rect 19432 6137 19441 6171
rect 19441 6137 19475 6171
rect 19475 6137 19484 6171
rect 19432 6128 19484 6137
rect 20444 6171 20496 6180
rect 20444 6137 20453 6171
rect 20453 6137 20487 6171
rect 20487 6137 20496 6171
rect 20996 6171 21048 6180
rect 20444 6128 20496 6137
rect 20996 6137 21005 6171
rect 21005 6137 21039 6171
rect 21039 6137 21048 6171
rect 20996 6128 21048 6137
rect 21916 6196 21968 6248
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 21640 6103 21692 6112
rect 21640 6069 21649 6103
rect 21649 6069 21683 6103
rect 21683 6069 21692 6103
rect 21640 6060 21692 6069
rect 23112 6060 23164 6112
rect 23940 6196 23992 6248
rect 25320 6196 25372 6248
rect 29736 6239 29788 6248
rect 29736 6205 29745 6239
rect 29745 6205 29779 6239
rect 29779 6205 29788 6239
rect 29736 6196 29788 6205
rect 32128 6409 32137 6443
rect 32137 6409 32171 6443
rect 32171 6409 32180 6443
rect 32128 6400 32180 6409
rect 32220 6400 32272 6452
rect 34152 6400 34204 6452
rect 35900 6443 35952 6452
rect 35900 6409 35909 6443
rect 35909 6409 35943 6443
rect 35943 6409 35952 6443
rect 35900 6400 35952 6409
rect 35348 6264 35400 6316
rect 35624 6264 35676 6316
rect 31576 6239 31628 6248
rect 31576 6205 31585 6239
rect 31585 6205 31619 6239
rect 31619 6205 31628 6239
rect 31576 6196 31628 6205
rect 34428 6196 34480 6248
rect 35808 6196 35860 6248
rect 24400 6171 24452 6180
rect 24400 6137 24409 6171
rect 24409 6137 24443 6171
rect 24443 6137 24452 6171
rect 24400 6128 24452 6137
rect 24676 6128 24728 6180
rect 24860 6128 24912 6180
rect 25964 6128 26016 6180
rect 27068 6171 27120 6180
rect 27068 6137 27077 6171
rect 27077 6137 27111 6171
rect 27111 6137 27120 6171
rect 27068 6128 27120 6137
rect 26056 6060 26108 6112
rect 26884 6060 26936 6112
rect 27804 6128 27856 6180
rect 31852 6171 31904 6180
rect 31852 6137 31861 6171
rect 31861 6137 31895 6171
rect 31895 6137 31904 6171
rect 31852 6128 31904 6137
rect 33324 6171 33376 6180
rect 33324 6137 33333 6171
rect 33333 6137 33367 6171
rect 33367 6137 33376 6171
rect 33324 6128 33376 6137
rect 30472 6060 30524 6112
rect 30932 6060 30984 6112
rect 33140 6103 33192 6112
rect 33140 6069 33149 6103
rect 33149 6069 33183 6103
rect 33183 6069 33192 6103
rect 35992 6128 36044 6180
rect 36544 6171 36596 6180
rect 36544 6137 36553 6171
rect 36553 6137 36587 6171
rect 36587 6137 36596 6171
rect 36544 6128 36596 6137
rect 33140 6060 33192 6069
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 4620 5856 4672 5908
rect 5356 5856 5408 5908
rect 7472 5899 7524 5908
rect 2136 5788 2188 5840
rect 4160 5788 4212 5840
rect 1860 5720 1912 5772
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 3976 5720 4028 5772
rect 5264 5788 5316 5840
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 8300 5856 8352 5908
rect 12624 5856 12676 5908
rect 12716 5856 12768 5908
rect 14648 5899 14700 5908
rect 14648 5865 14657 5899
rect 14657 5865 14691 5899
rect 14691 5865 14700 5899
rect 14648 5856 14700 5865
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 22376 5899 22428 5908
rect 22376 5865 22385 5899
rect 22385 5865 22419 5899
rect 22419 5865 22428 5899
rect 22376 5856 22428 5865
rect 23940 5856 23992 5908
rect 25228 5899 25280 5908
rect 25228 5865 25237 5899
rect 25237 5865 25271 5899
rect 25271 5865 25280 5899
rect 25228 5856 25280 5865
rect 29552 5856 29604 5908
rect 31208 5899 31260 5908
rect 31208 5865 31217 5899
rect 31217 5865 31251 5899
rect 31251 5865 31260 5899
rect 31208 5856 31260 5865
rect 33048 5899 33100 5908
rect 33048 5865 33057 5899
rect 33057 5865 33091 5899
rect 33091 5865 33100 5899
rect 33048 5856 33100 5865
rect 33692 5899 33744 5908
rect 33692 5865 33701 5899
rect 33701 5865 33735 5899
rect 33735 5865 33744 5899
rect 33692 5856 33744 5865
rect 34796 5899 34848 5908
rect 34796 5865 34805 5899
rect 34805 5865 34839 5899
rect 34839 5865 34848 5899
rect 34796 5856 34848 5865
rect 35072 5899 35124 5908
rect 35072 5865 35081 5899
rect 35081 5865 35115 5899
rect 35115 5865 35124 5899
rect 35072 5856 35124 5865
rect 36544 5856 36596 5908
rect 6276 5831 6328 5840
rect 6276 5797 6285 5831
rect 6285 5797 6319 5831
rect 6319 5797 6328 5831
rect 6276 5788 6328 5797
rect 7288 5788 7340 5840
rect 8116 5788 8168 5840
rect 7196 5720 7248 5772
rect 8484 5720 8536 5772
rect 10416 5788 10468 5840
rect 11980 5788 12032 5840
rect 14004 5788 14056 5840
rect 16396 5788 16448 5840
rect 16948 5788 17000 5840
rect 14832 5720 14884 5772
rect 15200 5720 15252 5772
rect 20444 5788 20496 5840
rect 20812 5788 20864 5840
rect 21732 5788 21784 5840
rect 22284 5788 22336 5840
rect 23848 5788 23900 5840
rect 24860 5788 24912 5840
rect 26332 5788 26384 5840
rect 28264 5831 28316 5840
rect 28264 5797 28273 5831
rect 28273 5797 28307 5831
rect 28307 5797 28316 5831
rect 28264 5788 28316 5797
rect 30472 5788 30524 5840
rect 32220 5788 32272 5840
rect 34152 5788 34204 5840
rect 35440 5831 35492 5840
rect 35440 5797 35449 5831
rect 35449 5797 35483 5831
rect 35483 5797 35492 5831
rect 35440 5788 35492 5797
rect 35808 5831 35860 5840
rect 35808 5797 35817 5831
rect 35817 5797 35851 5831
rect 35851 5797 35860 5831
rect 35808 5788 35860 5797
rect 4804 5652 4856 5704
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 10048 5695 10100 5704
rect 5632 5584 5684 5636
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 572 5516 624 5568
rect 8392 5516 8444 5568
rect 10508 5516 10560 5568
rect 11428 5559 11480 5568
rect 11428 5525 11437 5559
rect 11437 5525 11471 5559
rect 11471 5525 11480 5559
rect 12072 5652 12124 5704
rect 15292 5652 15344 5704
rect 18972 5695 19024 5704
rect 12532 5584 12584 5636
rect 13452 5584 13504 5636
rect 18972 5661 18981 5695
rect 18981 5661 19015 5695
rect 19015 5661 19024 5695
rect 18972 5652 19024 5661
rect 20720 5652 20772 5704
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 21916 5652 21968 5704
rect 33140 5720 33192 5772
rect 34060 5720 34112 5772
rect 23112 5652 23164 5704
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 26240 5652 26292 5704
rect 27252 5695 27304 5704
rect 27252 5661 27261 5695
rect 27261 5661 27295 5695
rect 27295 5661 27304 5695
rect 27252 5652 27304 5661
rect 28172 5695 28224 5704
rect 28172 5661 28181 5695
rect 28181 5661 28215 5695
rect 28215 5661 28224 5695
rect 28172 5652 28224 5661
rect 28356 5652 28408 5704
rect 29276 5695 29328 5704
rect 19064 5584 19116 5636
rect 26332 5584 26384 5636
rect 29276 5661 29285 5695
rect 29285 5661 29319 5695
rect 29319 5661 29328 5695
rect 29276 5652 29328 5661
rect 29736 5652 29788 5704
rect 30288 5695 30340 5704
rect 30288 5661 30297 5695
rect 30297 5661 30331 5695
rect 30331 5661 30340 5695
rect 30288 5652 30340 5661
rect 31944 5652 31996 5704
rect 33048 5652 33100 5704
rect 35072 5652 35124 5704
rect 35992 5695 36044 5704
rect 35992 5661 36001 5695
rect 36001 5661 36035 5695
rect 36035 5661 36044 5695
rect 35992 5652 36044 5661
rect 11428 5516 11480 5525
rect 13820 5516 13872 5568
rect 15844 5559 15896 5568
rect 15844 5525 15853 5559
rect 15853 5525 15887 5559
rect 15887 5525 15896 5559
rect 15844 5516 15896 5525
rect 16856 5516 16908 5568
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 20628 5516 20680 5568
rect 28172 5516 28224 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2688 5312 2740 5364
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 6276 5312 6328 5364
rect 7196 5355 7248 5364
rect 7196 5321 7205 5355
rect 7205 5321 7239 5355
rect 7239 5321 7248 5355
rect 7196 5312 7248 5321
rect 8300 5312 8352 5364
rect 2412 5244 2464 5296
rect 3056 5176 3108 5228
rect 3884 5176 3936 5228
rect 4712 5176 4764 5228
rect 6184 5176 6236 5228
rect 9588 5312 9640 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 17040 5355 17092 5364
rect 17040 5321 17049 5355
rect 17049 5321 17083 5355
rect 17083 5321 17092 5355
rect 17040 5312 17092 5321
rect 22284 5312 22336 5364
rect 24860 5355 24912 5364
rect 24860 5321 24869 5355
rect 24869 5321 24903 5355
rect 24903 5321 24912 5355
rect 24860 5312 24912 5321
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 28264 5312 28316 5364
rect 28356 5312 28408 5364
rect 33140 5312 33192 5364
rect 34060 5312 34112 5364
rect 34612 5312 34664 5364
rect 34980 5312 35032 5364
rect 35624 5312 35676 5364
rect 35900 5355 35952 5364
rect 35900 5321 35909 5355
rect 35909 5321 35943 5355
rect 35943 5321 35952 5355
rect 35900 5312 35952 5321
rect 12716 5244 12768 5296
rect 13084 5244 13136 5296
rect 18236 5287 18288 5296
rect 11980 5176 12032 5228
rect 13728 5176 13780 5228
rect 6828 5108 6880 5160
rect 9588 5151 9640 5160
rect 8116 5040 8168 5092
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 12532 5108 12584 5160
rect 12992 5108 13044 5160
rect 11520 5083 11572 5092
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 18236 5253 18245 5287
rect 18245 5253 18279 5287
rect 18279 5253 18288 5287
rect 18236 5244 18288 5253
rect 22100 5287 22152 5296
rect 22100 5253 22109 5287
rect 22109 5253 22143 5287
rect 22143 5253 22152 5287
rect 22100 5244 22152 5253
rect 26056 5244 26108 5296
rect 15384 5176 15436 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 20720 5176 20772 5228
rect 21732 5219 21784 5228
rect 21732 5185 21741 5219
rect 21741 5185 21775 5219
rect 21775 5185 21784 5219
rect 21732 5176 21784 5185
rect 26976 5219 27028 5228
rect 26976 5185 26985 5219
rect 26985 5185 27019 5219
rect 27019 5185 27028 5219
rect 26976 5176 27028 5185
rect 27252 5219 27304 5228
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 27252 5176 27304 5185
rect 28172 5176 28224 5228
rect 32220 5244 32272 5296
rect 34704 5244 34756 5296
rect 36636 5244 36688 5296
rect 31852 5176 31904 5228
rect 32956 5176 33008 5228
rect 34980 5219 35032 5228
rect 34980 5185 34989 5219
rect 34989 5185 35023 5219
rect 35023 5185 35032 5219
rect 34980 5176 35032 5185
rect 35256 5219 35308 5228
rect 35256 5185 35265 5219
rect 35265 5185 35299 5219
rect 35299 5185 35308 5219
rect 35256 5176 35308 5185
rect 35992 5176 36044 5228
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19156 5151 19208 5160
rect 19156 5117 19165 5151
rect 19165 5117 19199 5151
rect 19199 5117 19208 5151
rect 19156 5108 19208 5117
rect 19708 5108 19760 5160
rect 24308 5108 24360 5160
rect 30472 5108 30524 5160
rect 30840 5151 30892 5160
rect 30840 5117 30849 5151
rect 30849 5117 30883 5151
rect 30883 5117 30892 5151
rect 30840 5108 30892 5117
rect 15384 5083 15436 5092
rect 15384 5049 15393 5083
rect 15393 5049 15427 5083
rect 15427 5049 15436 5083
rect 15384 5040 15436 5049
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 15844 5040 15896 5092
rect 16948 4972 17000 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 20536 4972 20588 5024
rect 20812 5015 20864 5024
rect 20812 4981 20821 5015
rect 20821 4981 20855 5015
rect 20855 4981 20864 5015
rect 20812 4972 20864 4981
rect 24860 5040 24912 5092
rect 25412 5083 25464 5092
rect 25412 5049 25421 5083
rect 25421 5049 25455 5083
rect 25455 5049 25464 5083
rect 25412 5040 25464 5049
rect 29368 5083 29420 5092
rect 22560 5015 22612 5024
rect 22560 4981 22569 5015
rect 22569 4981 22603 5015
rect 22603 4981 22612 5015
rect 22560 4972 22612 4981
rect 23112 5015 23164 5024
rect 23112 4981 23121 5015
rect 23121 4981 23155 5015
rect 23155 4981 23164 5015
rect 23112 4972 23164 4981
rect 24584 5015 24636 5024
rect 24584 4981 24593 5015
rect 24593 4981 24627 5015
rect 24627 4981 24636 5015
rect 24584 4972 24636 4981
rect 29368 5049 29377 5083
rect 29377 5049 29411 5083
rect 29411 5049 29420 5083
rect 29368 5040 29420 5049
rect 32220 5040 32272 5092
rect 33692 5040 33744 5092
rect 35072 5083 35124 5092
rect 35072 5049 35081 5083
rect 35081 5049 35115 5083
rect 35115 5049 35124 5083
rect 35072 5040 35124 5049
rect 36360 5040 36412 5092
rect 36636 5083 36688 5092
rect 36636 5049 36645 5083
rect 36645 5049 36679 5083
rect 36679 5049 36688 5083
rect 36636 5040 36688 5049
rect 30380 4972 30432 5024
rect 30932 4972 30984 5024
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 1860 4768 1912 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 6092 4768 6144 4820
rect 12164 4811 12216 4820
rect 12164 4777 12173 4811
rect 12173 4777 12207 4811
rect 12207 4777 12216 4811
rect 12164 4768 12216 4777
rect 12624 4768 12676 4820
rect 14004 4811 14056 4820
rect 2412 4700 2464 4752
rect 3608 4700 3660 4752
rect 3976 4700 4028 4752
rect 8116 4700 8168 4752
rect 6644 4632 6696 4684
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 9220 4700 9272 4752
rect 10508 4700 10560 4752
rect 11980 4700 12032 4752
rect 12808 4743 12860 4752
rect 12808 4709 12817 4743
rect 12817 4709 12851 4743
rect 12851 4709 12860 4743
rect 12808 4700 12860 4709
rect 13084 4743 13136 4752
rect 13084 4709 13093 4743
rect 13093 4709 13127 4743
rect 13127 4709 13136 4743
rect 13084 4700 13136 4709
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 20536 4768 20588 4820
rect 21916 4811 21968 4820
rect 21916 4777 21925 4811
rect 21925 4777 21959 4811
rect 21959 4777 21968 4811
rect 21916 4768 21968 4777
rect 23572 4768 23624 4820
rect 24308 4811 24360 4820
rect 24308 4777 24317 4811
rect 24317 4777 24351 4811
rect 24351 4777 24360 4811
rect 24308 4768 24360 4777
rect 26332 4811 26384 4820
rect 26332 4777 26341 4811
rect 26341 4777 26375 4811
rect 26375 4777 26384 4811
rect 26332 4768 26384 4777
rect 29368 4811 29420 4820
rect 29368 4777 29377 4811
rect 29377 4777 29411 4811
rect 29411 4777 29420 4811
rect 29368 4768 29420 4777
rect 32956 4811 33008 4820
rect 32956 4777 32965 4811
rect 32965 4777 32999 4811
rect 32999 4777 33008 4811
rect 32956 4768 33008 4777
rect 34980 4811 35032 4820
rect 34980 4777 34989 4811
rect 34989 4777 35023 4811
rect 35023 4777 35032 4811
rect 34980 4768 35032 4777
rect 35072 4768 35124 4820
rect 36360 4768 36412 4820
rect 13544 4700 13596 4752
rect 14188 4700 14240 4752
rect 19156 4700 19208 4752
rect 19892 4743 19944 4752
rect 19892 4709 19901 4743
rect 19901 4709 19935 4743
rect 19935 4709 19944 4743
rect 19892 4700 19944 4709
rect 20812 4700 20864 4752
rect 21732 4700 21784 4752
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 15844 4675 15896 4684
rect 15844 4641 15853 4675
rect 15853 4641 15887 4675
rect 15887 4641 15896 4675
rect 15844 4632 15896 4641
rect 2596 4564 2648 4616
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 7472 4564 7524 4616
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 17776 4632 17828 4684
rect 18328 4632 18380 4684
rect 24032 4743 24084 4752
rect 24032 4709 24041 4743
rect 24041 4709 24075 4743
rect 24075 4709 24084 4743
rect 24032 4700 24084 4709
rect 26240 4700 26292 4752
rect 28264 4743 28316 4752
rect 28264 4709 28273 4743
rect 28273 4709 28307 4743
rect 28307 4709 28316 4743
rect 28264 4700 28316 4709
rect 31208 4743 31260 4752
rect 31208 4709 31217 4743
rect 31217 4709 31251 4743
rect 31251 4709 31260 4743
rect 31208 4700 31260 4709
rect 33692 4700 33744 4752
rect 35900 4700 35952 4752
rect 23756 4675 23808 4684
rect 23756 4641 23765 4675
rect 23765 4641 23799 4675
rect 23799 4641 23808 4675
rect 23756 4632 23808 4641
rect 24952 4675 25004 4684
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 16672 4564 16724 4616
rect 21272 4564 21324 4616
rect 22560 4564 22612 4616
rect 25136 4564 25188 4616
rect 30380 4632 30432 4684
rect 30932 4675 30984 4684
rect 30932 4641 30941 4675
rect 30941 4641 30975 4675
rect 30975 4641 30984 4675
rect 30932 4632 30984 4641
rect 26148 4564 26200 4616
rect 27252 4564 27304 4616
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 28816 4607 28868 4616
rect 28816 4573 28825 4607
rect 28825 4573 28859 4607
rect 28859 4573 28868 4607
rect 28816 4564 28868 4573
rect 32128 4607 32180 4616
rect 32128 4573 32137 4607
rect 32137 4573 32171 4607
rect 32171 4573 32180 4607
rect 32128 4564 32180 4573
rect 33968 4564 34020 4616
rect 35164 4607 35216 4616
rect 35164 4573 35173 4607
rect 35173 4573 35207 4607
rect 35207 4573 35216 4607
rect 35164 4564 35216 4573
rect 8300 4496 8352 4548
rect 8852 4496 8904 4548
rect 9588 4496 9640 4548
rect 18052 4539 18104 4548
rect 18052 4505 18061 4539
rect 18061 4505 18095 4539
rect 18095 4505 18104 4539
rect 18052 4496 18104 4505
rect 27160 4539 27212 4548
rect 27160 4505 27169 4539
rect 27169 4505 27203 4539
rect 27203 4505 27212 4539
rect 32588 4539 32640 4548
rect 27160 4496 27212 4505
rect 32588 4505 32597 4539
rect 32597 4505 32631 4539
rect 32631 4505 32640 4539
rect 32588 4496 32640 4505
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 8116 4428 8168 4480
rect 8208 4428 8260 4480
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 15108 4471 15160 4480
rect 15108 4437 15117 4471
rect 15117 4437 15151 4471
rect 15151 4437 15160 4471
rect 15108 4428 15160 4437
rect 16304 4428 16356 4480
rect 16948 4428 17000 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 18236 4428 18288 4480
rect 22652 4428 22704 4480
rect 28356 4428 28408 4480
rect 28724 4428 28776 4480
rect 31484 4471 31536 4480
rect 31484 4437 31493 4471
rect 31493 4437 31527 4471
rect 31527 4437 31536 4471
rect 31484 4428 31536 4437
rect 34612 4428 34664 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 2412 4267 2464 4276
rect 2412 4233 2421 4267
rect 2421 4233 2455 4267
rect 2455 4233 2464 4267
rect 2412 4224 2464 4233
rect 3976 4267 4028 4276
rect 3976 4233 3985 4267
rect 3985 4233 4019 4267
rect 4019 4233 4028 4267
rect 3976 4224 4028 4233
rect 6828 4224 6880 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 11980 4224 12032 4276
rect 13912 4224 13964 4276
rect 18052 4224 18104 4276
rect 20812 4224 20864 4276
rect 21272 4267 21324 4276
rect 21272 4233 21281 4267
rect 21281 4233 21315 4267
rect 21315 4233 21324 4267
rect 21272 4224 21324 4233
rect 21364 4224 21416 4276
rect 22284 4224 22336 4276
rect 23480 4224 23532 4276
rect 28264 4224 28316 4276
rect 30380 4224 30432 4276
rect 32220 4224 32272 4276
rect 33692 4267 33744 4276
rect 33692 4233 33701 4267
rect 33701 4233 33735 4267
rect 33735 4233 33744 4267
rect 33692 4224 33744 4233
rect 35900 4267 35952 4276
rect 35900 4233 35909 4267
rect 35909 4233 35943 4267
rect 35943 4233 35952 4267
rect 35900 4224 35952 4233
rect 35992 4224 36044 4276
rect 3240 4156 3292 4208
rect 2964 4088 3016 4140
rect 4804 4156 4856 4208
rect 6644 4156 6696 4208
rect 16580 4199 16632 4208
rect 16580 4165 16589 4199
rect 16589 4165 16623 4199
rect 16623 4165 16632 4199
rect 16580 4156 16632 4165
rect 17132 4156 17184 4208
rect 17592 4156 17644 4208
rect 4252 4088 4304 4140
rect 4712 4088 4764 4140
rect 7472 4088 7524 4140
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 11428 4088 11480 4140
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 6092 4020 6144 4072
rect 2504 3952 2556 4004
rect 4252 3995 4304 4004
rect 1952 3884 2004 3936
rect 4252 3961 4261 3995
rect 4261 3961 4295 3995
rect 4295 3961 4304 3995
rect 4252 3952 4304 3961
rect 2872 3884 2924 3936
rect 5816 3952 5868 4004
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6460 3884 6512 3936
rect 7288 3952 7340 4004
rect 7748 3995 7800 4004
rect 7748 3961 7757 3995
rect 7757 3961 7791 3995
rect 7791 3961 7800 3995
rect 7748 3952 7800 3961
rect 9588 3995 9640 4004
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 8116 3884 8168 3936
rect 9588 3961 9597 3995
rect 9597 3961 9631 3995
rect 9631 3961 9640 3995
rect 9588 3952 9640 3961
rect 10784 3952 10836 4004
rect 11060 3952 11112 4004
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 15292 4088 15344 4140
rect 16304 4088 16356 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 13820 4020 13872 4029
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 18236 4020 18288 4072
rect 19892 4088 19944 4140
rect 20628 4088 20680 4140
rect 23388 4088 23440 4140
rect 23756 4156 23808 4208
rect 24952 4156 25004 4208
rect 30932 4131 30984 4140
rect 30932 4097 30941 4131
rect 30941 4097 30975 4131
rect 30975 4097 30984 4131
rect 30932 4088 30984 4097
rect 34612 4131 34664 4140
rect 18788 4063 18840 4072
rect 18788 4029 18797 4063
rect 18797 4029 18831 4063
rect 18831 4029 18840 4063
rect 18788 4020 18840 4029
rect 21824 4063 21876 4072
rect 21824 4029 21833 4063
rect 21833 4029 21867 4063
rect 21867 4029 21876 4063
rect 21824 4020 21876 4029
rect 22192 4063 22244 4072
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 25504 4020 25556 4072
rect 26240 4020 26292 4072
rect 26332 4020 26384 4072
rect 29552 4063 29604 4072
rect 29552 4029 29561 4063
rect 29561 4029 29595 4063
rect 29595 4029 29604 4063
rect 29552 4020 29604 4029
rect 29920 4063 29972 4072
rect 29920 4029 29929 4063
rect 29929 4029 29963 4063
rect 29963 4029 29972 4063
rect 29920 4020 29972 4029
rect 32588 4063 32640 4072
rect 32588 4029 32597 4063
rect 32597 4029 32631 4063
rect 32631 4029 32640 4063
rect 32588 4020 32640 4029
rect 34612 4097 34621 4131
rect 34621 4097 34655 4131
rect 34655 4097 34664 4131
rect 34612 4088 34664 4097
rect 35256 4131 35308 4140
rect 35256 4097 35265 4131
rect 35265 4097 35299 4131
rect 35299 4097 35308 4131
rect 35256 4088 35308 4097
rect 36452 4063 36504 4072
rect 36452 4029 36461 4063
rect 36461 4029 36495 4063
rect 36495 4029 36504 4063
rect 37004 4063 37056 4072
rect 36452 4020 36504 4029
rect 37004 4029 37013 4063
rect 37013 4029 37047 4063
rect 37047 4029 37056 4063
rect 37004 4020 37056 4029
rect 37556 4063 37608 4072
rect 37556 4029 37600 4063
rect 37600 4029 37608 4063
rect 37556 4020 37608 4029
rect 12808 3952 12860 4004
rect 15200 3952 15252 4004
rect 16488 3952 16540 4004
rect 17040 3995 17092 4004
rect 17040 3961 17049 3995
rect 17049 3961 17083 3995
rect 17083 3961 17092 3995
rect 17040 3952 17092 3961
rect 17776 3952 17828 4004
rect 19156 3995 19208 4004
rect 19156 3961 19165 3995
rect 19165 3961 19199 3995
rect 19199 3961 19208 3995
rect 19156 3952 19208 3961
rect 25044 3952 25096 4004
rect 28724 3952 28776 4004
rect 30104 3995 30156 4004
rect 30104 3961 30113 3995
rect 30113 3961 30147 3995
rect 30147 3961 30156 3995
rect 30104 3952 30156 3961
rect 31116 3995 31168 4004
rect 31116 3961 31125 3995
rect 31125 3961 31159 3995
rect 31159 3961 31168 3995
rect 31116 3952 31168 3961
rect 31484 3952 31536 4004
rect 31576 3952 31628 4004
rect 33324 3995 33376 4004
rect 33324 3961 33333 3995
rect 33333 3961 33367 3995
rect 33367 3961 33376 3995
rect 33324 3952 33376 3961
rect 10232 3884 10284 3893
rect 13728 3884 13780 3936
rect 14924 3884 14976 3936
rect 16580 3884 16632 3936
rect 19800 3927 19852 3936
rect 19800 3893 19809 3927
rect 19809 3893 19843 3927
rect 19843 3893 19852 3927
rect 19800 3884 19852 3893
rect 22192 3884 22244 3936
rect 24216 3884 24268 3936
rect 26332 3884 26384 3936
rect 27344 3884 27396 3936
rect 28172 3884 28224 3936
rect 33968 3927 34020 3936
rect 33968 3893 33977 3927
rect 33977 3893 34011 3927
rect 34011 3893 34020 3927
rect 33968 3884 34020 3893
rect 34612 3884 34664 3936
rect 36820 3884 36872 3936
rect 37280 3884 37332 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 2780 3680 2832 3732
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 5356 3680 5408 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 8024 3680 8076 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 10140 3680 10192 3732
rect 11244 3680 11296 3732
rect 12440 3680 12492 3732
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 15108 3680 15160 3732
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 15844 3680 15896 3732
rect 17868 3723 17920 3732
rect 17868 3689 17877 3723
rect 17877 3689 17911 3723
rect 17911 3689 17920 3723
rect 17868 3680 17920 3689
rect 1768 3612 1820 3664
rect 2412 3612 2464 3664
rect 2872 3655 2924 3664
rect 2872 3621 2881 3655
rect 2881 3621 2915 3655
rect 2915 3621 2924 3655
rect 2872 3612 2924 3621
rect 4252 3612 4304 3664
rect 3700 3544 3752 3596
rect 1676 3476 1728 3528
rect 4160 3544 4212 3596
rect 5816 3587 5868 3596
rect 5816 3553 5825 3587
rect 5825 3553 5859 3587
rect 5859 3553 5868 3587
rect 5816 3544 5868 3553
rect 6276 3544 6328 3596
rect 8116 3612 8168 3664
rect 8760 3612 8812 3664
rect 10876 3612 10928 3664
rect 12808 3655 12860 3664
rect 12808 3621 12817 3655
rect 12817 3621 12851 3655
rect 12851 3621 12860 3655
rect 12808 3612 12860 3621
rect 13636 3612 13688 3664
rect 16396 3655 16448 3664
rect 16396 3621 16405 3655
rect 16405 3621 16439 3655
rect 16439 3621 16448 3655
rect 16396 3612 16448 3621
rect 17500 3612 17552 3664
rect 17776 3612 17828 3664
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 11060 3587 11112 3596
rect 11060 3553 11069 3587
rect 11069 3553 11103 3587
rect 11103 3553 11112 3587
rect 11060 3544 11112 3553
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 12992 3587 13044 3596
rect 12992 3553 12998 3587
rect 12998 3553 13044 3587
rect 12992 3544 13044 3553
rect 16488 3544 16540 3596
rect 16948 3544 17000 3596
rect 17960 3544 18012 3596
rect 22192 3723 22244 3732
rect 22192 3689 22201 3723
rect 22201 3689 22235 3723
rect 22235 3689 22244 3723
rect 22192 3680 22244 3689
rect 19892 3655 19944 3664
rect 19892 3621 19901 3655
rect 19901 3621 19935 3655
rect 19935 3621 19944 3655
rect 19892 3612 19944 3621
rect 21272 3612 21324 3664
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 19616 3587 19668 3596
rect 5908 3476 5960 3528
rect 8208 3476 8260 3528
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 13268 3476 13320 3528
rect 14096 3476 14148 3528
rect 15016 3476 15068 3528
rect 16672 3476 16724 3528
rect 17132 3476 17184 3528
rect 19616 3553 19625 3587
rect 19625 3553 19659 3587
rect 19659 3553 19668 3587
rect 19616 3544 19668 3553
rect 20076 3544 20128 3596
rect 20812 3544 20864 3596
rect 23480 3680 23532 3732
rect 25136 3723 25188 3732
rect 23112 3612 23164 3664
rect 24216 3655 24268 3664
rect 24216 3621 24225 3655
rect 24225 3621 24259 3655
rect 24259 3621 24268 3655
rect 24216 3612 24268 3621
rect 25136 3689 25145 3723
rect 25145 3689 25179 3723
rect 25179 3689 25188 3723
rect 25136 3680 25188 3689
rect 26240 3723 26292 3732
rect 26240 3689 26249 3723
rect 26249 3689 26283 3723
rect 26283 3689 26292 3723
rect 26240 3680 26292 3689
rect 28080 3723 28132 3732
rect 28080 3689 28089 3723
rect 28089 3689 28123 3723
rect 28123 3689 28132 3723
rect 28080 3680 28132 3689
rect 30104 3723 30156 3732
rect 30104 3689 30113 3723
rect 30113 3689 30147 3723
rect 30147 3689 30156 3723
rect 30104 3680 30156 3689
rect 26148 3612 26200 3664
rect 26884 3612 26936 3664
rect 27344 3655 27396 3664
rect 27344 3621 27353 3655
rect 27353 3621 27387 3655
rect 27387 3621 27396 3655
rect 27344 3612 27396 3621
rect 28724 3612 28776 3664
rect 31484 3680 31536 3732
rect 30472 3612 30524 3664
rect 33784 3612 33836 3664
rect 36268 3612 36320 3664
rect 31116 3544 31168 3596
rect 31576 3544 31628 3596
rect 32220 3587 32272 3596
rect 32220 3553 32229 3587
rect 32229 3553 32263 3587
rect 32263 3553 32272 3587
rect 32220 3544 32272 3553
rect 20628 3476 20680 3528
rect 24032 3476 24084 3528
rect 24492 3519 24544 3528
rect 24492 3485 24501 3519
rect 24501 3485 24535 3519
rect 24535 3485 24544 3519
rect 24492 3476 24544 3485
rect 24860 3476 24912 3528
rect 26332 3476 26384 3528
rect 26792 3476 26844 3528
rect 28172 3519 28224 3528
rect 28172 3485 28181 3519
rect 28181 3485 28215 3519
rect 28215 3485 28224 3519
rect 28172 3476 28224 3485
rect 31484 3476 31536 3528
rect 31668 3476 31720 3528
rect 33324 3544 33376 3596
rect 35164 3519 35216 3528
rect 35164 3485 35173 3519
rect 35173 3485 35207 3519
rect 35207 3485 35216 3519
rect 35164 3476 35216 3485
rect 35900 3476 35952 3528
rect 35992 3519 36044 3528
rect 35992 3485 36001 3519
rect 36001 3485 36035 3519
rect 36035 3485 36044 3519
rect 35992 3476 36044 3485
rect 7748 3408 7800 3460
rect 13912 3408 13964 3460
rect 18236 3408 18288 3460
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 8760 3340 8812 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 14004 3340 14056 3392
rect 15752 3340 15804 3392
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 21824 3383 21876 3392
rect 21824 3349 21833 3383
rect 21833 3349 21867 3383
rect 21867 3349 21876 3383
rect 21824 3340 21876 3349
rect 25504 3383 25556 3392
rect 25504 3349 25513 3383
rect 25513 3349 25547 3383
rect 25547 3349 25556 3383
rect 25504 3340 25556 3349
rect 28908 3340 28960 3392
rect 29368 3340 29420 3392
rect 29552 3340 29604 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 1768 3136 1820 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 4160 3136 4212 3188
rect 2964 3068 3016 3120
rect 1492 3000 1544 3052
rect 5448 3136 5500 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 8116 3179 8168 3188
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 9496 3136 9548 3188
rect 9956 3136 10008 3188
rect 10232 3136 10284 3188
rect 12164 3179 12216 3188
rect 5264 3111 5316 3120
rect 5264 3077 5273 3111
rect 5273 3077 5307 3111
rect 5307 3077 5316 3111
rect 5264 3068 5316 3077
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 13268 3136 13320 3188
rect 12532 3111 12584 3120
rect 12532 3077 12541 3111
rect 12541 3077 12575 3111
rect 12575 3077 12584 3111
rect 15108 3136 15160 3188
rect 15752 3136 15804 3188
rect 16304 3136 16356 3188
rect 17132 3136 17184 3188
rect 17592 3136 17644 3188
rect 20812 3136 20864 3188
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 21640 3136 21692 3188
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 24216 3179 24268 3188
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 26884 3136 26936 3188
rect 28172 3136 28224 3188
rect 28724 3179 28776 3188
rect 28724 3145 28733 3179
rect 28733 3145 28767 3179
rect 28767 3145 28776 3179
rect 28724 3136 28776 3145
rect 30472 3136 30524 3188
rect 32220 3136 32272 3188
rect 33324 3136 33376 3188
rect 34704 3179 34756 3188
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 35900 3179 35952 3188
rect 35900 3145 35909 3179
rect 35909 3145 35943 3179
rect 35943 3145 35952 3179
rect 35900 3136 35952 3145
rect 36268 3179 36320 3188
rect 36268 3145 36277 3179
rect 36277 3145 36311 3179
rect 36311 3145 36320 3179
rect 36268 3136 36320 3145
rect 37372 3136 37424 3188
rect 12532 3068 12584 3077
rect 13084 3043 13136 3052
rect 4712 2932 4764 2984
rect 5080 2932 5132 2984
rect 5448 2975 5500 2984
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 5816 2932 5868 2984
rect 6000 2932 6052 2984
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2504 2864 2556 2916
rect 5908 2907 5960 2916
rect 5908 2873 5917 2907
rect 5917 2873 5951 2907
rect 5951 2873 5960 2907
rect 5908 2864 5960 2873
rect 7104 2932 7156 2984
rect 7932 2932 7984 2984
rect 8852 2932 8904 2984
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 11612 2864 11664 2916
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 16028 3043 16080 3052
rect 14004 2975 14056 2984
rect 12164 2864 12216 2916
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 14188 2932 14240 2984
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 18420 3000 18472 3052
rect 27160 3111 27212 3120
rect 27160 3077 27169 3111
rect 27169 3077 27203 3111
rect 27203 3077 27212 3111
rect 27160 3068 27212 3077
rect 33692 3111 33744 3120
rect 33692 3077 33701 3111
rect 33701 3077 33735 3111
rect 33735 3077 33744 3111
rect 33692 3068 33744 3077
rect 22744 3043 22796 3052
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 17960 2932 18012 2984
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 18604 2932 18656 2984
rect 19800 2932 19852 2984
rect 22744 3009 22753 3043
rect 22753 3009 22787 3043
rect 22787 3009 22796 3043
rect 22744 3000 22796 3009
rect 29368 3000 29420 3052
rect 29644 3043 29696 3052
rect 29644 3009 29653 3043
rect 29653 3009 29687 3043
rect 29687 3009 29696 3043
rect 29644 3000 29696 3009
rect 30104 3000 30156 3052
rect 31944 3000 31996 3052
rect 33968 3000 34020 3052
rect 34980 3043 35032 3052
rect 34980 3009 34989 3043
rect 34989 3009 35023 3043
rect 35023 3009 35032 3043
rect 34980 3000 35032 3009
rect 35072 3000 35124 3052
rect 17776 2864 17828 2916
rect 19616 2864 19668 2916
rect 23388 2932 23440 2984
rect 24768 2975 24820 2984
rect 24768 2941 24777 2975
rect 24777 2941 24811 2975
rect 24811 2941 24820 2975
rect 24768 2932 24820 2941
rect 28080 2932 28132 2984
rect 30748 2975 30800 2984
rect 30748 2941 30757 2975
rect 30757 2941 30791 2975
rect 30791 2941 30800 2975
rect 30748 2932 30800 2941
rect 31300 2932 31352 2984
rect 31484 2932 31536 2984
rect 32312 2975 32364 2984
rect 32312 2941 32321 2975
rect 32321 2941 32355 2975
rect 32355 2941 32364 2975
rect 32312 2932 32364 2941
rect 32864 2975 32916 2984
rect 32864 2941 32873 2975
rect 32873 2941 32907 2975
rect 32907 2941 32916 2975
rect 32864 2932 32916 2941
rect 37004 2932 37056 2984
rect 23112 2907 23164 2916
rect 23112 2873 23121 2907
rect 23121 2873 23155 2907
rect 23155 2873 23164 2907
rect 23112 2864 23164 2873
rect 25044 2864 25096 2916
rect 2044 2796 2096 2805
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 13912 2796 13964 2848
rect 15016 2839 15068 2848
rect 15016 2805 15025 2839
rect 15025 2805 15059 2839
rect 15059 2805 15068 2839
rect 15016 2796 15068 2805
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 29460 2907 29512 2916
rect 29460 2873 29469 2907
rect 29469 2873 29503 2907
rect 29503 2873 29512 2907
rect 29460 2864 29512 2873
rect 34704 2864 34756 2916
rect 29736 2796 29788 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 2044 2592 2096 2601
rect 4712 2592 4764 2644
rect 6000 2592 6052 2644
rect 8024 2592 8076 2644
rect 8576 2592 8628 2644
rect 9496 2635 9548 2644
rect 4068 2524 4120 2576
rect 7932 2567 7984 2576
rect 1952 2388 2004 2440
rect 3424 2252 3476 2304
rect 5080 2456 5132 2508
rect 7932 2533 7941 2567
rect 7941 2533 7975 2567
rect 7975 2533 7984 2567
rect 8852 2567 8904 2576
rect 7932 2524 7984 2533
rect 5356 2456 5408 2508
rect 5816 2456 5868 2508
rect 6092 2456 6144 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8852 2533 8861 2567
rect 8861 2533 8895 2567
rect 8895 2533 8904 2567
rect 8852 2524 8904 2533
rect 8668 2388 8720 2440
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 12716 2592 12768 2644
rect 13268 2635 13320 2644
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 16580 2635 16632 2644
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 16580 2592 16632 2601
rect 9956 2567 10008 2576
rect 9956 2533 9965 2567
rect 9965 2533 9999 2567
rect 9999 2533 10008 2567
rect 9956 2524 10008 2533
rect 10508 2567 10560 2576
rect 10508 2533 10517 2567
rect 10517 2533 10551 2567
rect 10551 2533 10560 2567
rect 10508 2524 10560 2533
rect 11060 2524 11112 2576
rect 12900 2524 12952 2576
rect 11888 2388 11940 2440
rect 12624 2388 12676 2440
rect 14096 2456 14148 2508
rect 17316 2592 17368 2644
rect 17500 2635 17552 2644
rect 17500 2601 17509 2635
rect 17509 2601 17543 2635
rect 17543 2601 17552 2635
rect 17500 2592 17552 2601
rect 17592 2592 17644 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 18328 2567 18380 2576
rect 18328 2533 18337 2567
rect 18337 2533 18371 2567
rect 18371 2533 18380 2567
rect 18328 2524 18380 2533
rect 19800 2592 19852 2644
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 21364 2635 21416 2644
rect 21364 2601 21373 2635
rect 21373 2601 21407 2635
rect 21407 2601 21416 2635
rect 21364 2592 21416 2601
rect 23388 2635 23440 2644
rect 23388 2601 23397 2635
rect 23397 2601 23431 2635
rect 23431 2601 23440 2635
rect 23388 2592 23440 2601
rect 23572 2592 23624 2644
rect 24860 2592 24912 2644
rect 26332 2635 26384 2644
rect 20628 2567 20680 2576
rect 20628 2533 20637 2567
rect 20637 2533 20671 2567
rect 20671 2533 20680 2567
rect 20628 2524 20680 2533
rect 19984 2456 20036 2508
rect 24768 2524 24820 2576
rect 22652 2499 22704 2508
rect 22652 2465 22661 2499
rect 22661 2465 22695 2499
rect 22695 2465 22704 2499
rect 22652 2456 22704 2465
rect 15016 2320 15068 2372
rect 12808 2252 12860 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 15660 2388 15712 2440
rect 23572 2456 23624 2508
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 27252 2635 27304 2644
rect 27252 2601 27261 2635
rect 27261 2601 27295 2635
rect 27295 2601 27304 2635
rect 27252 2592 27304 2601
rect 28908 2592 28960 2644
rect 29460 2635 29512 2644
rect 29460 2601 29469 2635
rect 29469 2601 29503 2635
rect 29503 2601 29512 2635
rect 29460 2592 29512 2601
rect 29920 2592 29972 2644
rect 28172 2567 28224 2576
rect 26700 2499 26752 2508
rect 23388 2388 23440 2440
rect 26700 2465 26709 2499
rect 26709 2465 26743 2499
rect 26743 2465 26752 2499
rect 27712 2499 27764 2508
rect 26700 2456 26752 2465
rect 27712 2465 27721 2499
rect 27721 2465 27755 2499
rect 27755 2465 27764 2499
rect 27712 2456 27764 2465
rect 28172 2533 28181 2567
rect 28181 2533 28215 2567
rect 28215 2533 28224 2567
rect 28172 2524 28224 2533
rect 31300 2592 31352 2644
rect 31760 2592 31812 2644
rect 32864 2592 32916 2644
rect 34060 2635 34112 2644
rect 34060 2601 34069 2635
rect 34069 2601 34103 2635
rect 34103 2601 34112 2635
rect 34060 2592 34112 2601
rect 34980 2635 35032 2644
rect 34980 2601 34989 2635
rect 34989 2601 35023 2635
rect 35023 2601 35032 2635
rect 34980 2592 35032 2601
rect 35992 2635 36044 2644
rect 35992 2601 36001 2635
rect 36001 2601 36035 2635
rect 36035 2601 36044 2635
rect 35992 2592 36044 2601
rect 30104 2524 30156 2576
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 36360 2456 36412 2508
rect 30288 2431 30340 2440
rect 30288 2397 30297 2431
rect 30297 2397 30331 2431
rect 30331 2397 30340 2431
rect 30288 2388 30340 2397
rect 35900 2388 35952 2440
rect 17776 2320 17828 2372
rect 36360 2320 36412 2372
rect 20076 2295 20128 2304
rect 14832 2252 14884 2261
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 25964 2252 26016 2304
rect 31668 2252 31720 2304
rect 33140 2252 33192 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 22100 552 22152 604
rect 22284 552 22336 604
<< metal2 >>
rect 1398 15600 1454 15609
rect 1398 15535 1454 15544
rect 1412 10810 1440 15535
rect 6642 15520 6698 16000
rect 19982 15520 20038 16000
rect 33322 15520 33378 16000
rect 35530 15600 35586 15609
rect 35530 15535 35586 15544
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1504 12442 1532 14583
rect 1582 13832 1638 13841
rect 1582 13767 1638 13776
rect 1596 12986 1624 13767
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 2962 12880 3018 12889
rect 2962 12815 3018 12824
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11558 1716 12242
rect 1676 11552 1728 11558
rect 1674 11520 1676 11529
rect 1728 11520 1730 11529
rect 1674 11455 1730 11464
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 11014 1900 11154
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1872 10130 1900 10950
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1688 9518 1716 10066
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 570 8528 626 8537
rect 570 8463 626 8472
rect 584 7818 612 8463
rect 572 7812 624 7818
rect 572 7754 624 7760
rect 572 5568 624 5574
rect 572 5510 624 5516
rect 584 4865 612 5510
rect 570 4856 626 4865
rect 570 4791 626 4800
rect 1122 3768 1178 3777
rect 1122 3703 1178 3712
rect 1136 480 1164 3703
rect 1504 3058 1532 8774
rect 1688 7750 1716 8978
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7342 1716 7686
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1872 5778 1900 9930
rect 1964 8498 1992 12582
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2056 11694 2084 12038
rect 2424 11694 2452 12038
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2056 10742 2084 11630
rect 2424 11218 2452 11630
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 2044 10464 2096 10470
rect 2042 10432 2044 10441
rect 2096 10432 2098 10441
rect 2042 10367 2098 10376
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1964 6798 1992 8434
rect 2056 6866 2084 9386
rect 2134 8936 2190 8945
rect 2134 8871 2190 8880
rect 2148 8498 2176 8871
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2240 7954 2268 11086
rect 2424 10266 2452 11154
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2332 8838 2360 10066
rect 2516 9926 2544 10542
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2320 8832 2372 8838
rect 2318 8800 2320 8809
rect 2372 8800 2374 8809
rect 2318 8735 2374 8744
rect 2424 8566 2452 9454
rect 2516 9382 2544 9862
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9178 2544 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2516 8673 2544 9114
rect 2502 8664 2558 8673
rect 2502 8599 2558 8608
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2228 7948 2280 7954
rect 2280 7908 2360 7936
rect 2228 7890 2280 7896
rect 2332 7478 2360 7908
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2516 7274 2544 7958
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2056 6322 2084 6802
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2148 6186 2176 7142
rect 2516 6934 2544 7210
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2608 6798 2636 11562
rect 2700 11121 2728 12038
rect 2884 11898 2912 12242
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2792 9654 2820 10134
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2688 8968 2740 8974
rect 2740 8916 2820 8922
rect 2688 8910 2820 8916
rect 2700 8894 2820 8910
rect 2792 8294 2820 8894
rect 2884 8362 2912 9046
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2688 8084 2740 8090
rect 2884 8072 2912 8298
rect 2740 8044 2912 8072
rect 2688 8026 2740 8032
rect 2884 6866 2912 8044
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6458 2636 6734
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2148 5846 2176 6122
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1582 5400 1638 5409
rect 1582 5335 1584 5344
rect 1636 5335 1638 5344
rect 1584 5306 1636 5312
rect 1872 4826 1900 5714
rect 2778 5536 2834 5545
rect 2778 5471 2834 5480
rect 2688 5364 2740 5370
rect 2792 5352 2820 5471
rect 2976 5409 3004 12815
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 12646 5488 12718
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3344 11393 3372 11494
rect 3330 11384 3386 11393
rect 3330 11319 3386 11328
rect 3516 11008 3568 11014
rect 3422 10976 3478 10985
rect 3516 10950 3568 10956
rect 3422 10911 3478 10920
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3054 10160 3110 10169
rect 3054 10095 3056 10104
rect 3108 10095 3110 10104
rect 3056 10066 3108 10072
rect 3068 9722 3096 10066
rect 3240 9920 3292 9926
rect 3344 9897 3372 10542
rect 3240 9862 3292 9868
rect 3330 9888 3386 9897
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3054 8528 3110 8537
rect 3054 8463 3056 8472
rect 3108 8463 3110 8472
rect 3056 8434 3108 8440
rect 3068 6798 3096 8434
rect 3160 8362 3188 8570
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3160 8090 3188 8298
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5953 3188 6054
rect 3146 5944 3202 5953
rect 3146 5879 3202 5888
rect 3252 5778 3280 9862
rect 3330 9823 3386 9832
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 2740 5324 2820 5352
rect 2962 5400 3018 5409
rect 2962 5335 3018 5344
rect 2688 5306 2740 5312
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2424 4758 2452 5238
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2424 4282 2452 4694
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1768 3664 1820 3670
rect 1768 3606 1820 3612
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1688 2961 1716 3470
rect 1780 3194 1808 3606
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1674 2952 1730 2961
rect 1674 2887 1730 2896
rect 1688 2650 1716 2887
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1964 2446 1992 3878
rect 2424 3670 2452 4218
rect 2502 4040 2558 4049
rect 2502 3975 2504 3984
rect 2556 3975 2558 3984
rect 2504 3946 2556 3952
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2516 3482 2544 3946
rect 2608 3618 2636 4558
rect 3068 4486 3096 5170
rect 2688 4480 2740 4486
rect 3056 4480 3108 4486
rect 2688 4422 2740 4428
rect 3054 4448 3056 4457
rect 3108 4448 3110 4457
rect 2700 4026 2728 4422
rect 3054 4383 3110 4392
rect 3252 4214 3280 5714
rect 3344 5545 3372 9658
rect 3330 5536 3386 5545
rect 3330 5471 3386 5480
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2700 3998 2912 4026
rect 2884 3942 2912 3998
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2792 3618 2820 3674
rect 2884 3670 2912 3878
rect 2608 3590 2820 3618
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2516 3454 2820 3482
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2922 2544 3334
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2650 2084 2790
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2792 513 2820 3454
rect 2976 3126 3004 4082
rect 2964 3120 3016 3126
rect 3436 3097 3464 10911
rect 3528 10266 3556 10950
rect 3620 10305 3648 11494
rect 3606 10296 3662 10305
rect 3516 10260 3568 10266
rect 3606 10231 3662 10240
rect 3516 10202 3568 10208
rect 3528 9586 3556 10202
rect 3712 9602 3740 12582
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3988 11801 4016 12242
rect 4160 12096 4212 12102
rect 4066 12064 4122 12073
rect 4160 12038 4212 12044
rect 4066 11999 4122 12008
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 4080 10810 4108 11999
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3620 9574 3740 9602
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3528 8838 3556 9386
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 7546 3556 8774
rect 3620 8129 3648 9574
rect 3698 9480 3754 9489
rect 3698 9415 3700 9424
rect 3752 9415 3754 9424
rect 3700 9386 3752 9392
rect 3712 9110 3740 9386
rect 3882 9208 3938 9217
rect 3882 9143 3884 9152
rect 3936 9143 3938 9152
rect 3884 9114 3936 9120
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3712 8498 3740 9046
rect 3896 8566 3924 9114
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3790 8392 3846 8401
rect 3790 8327 3846 8336
rect 3804 8294 3832 8327
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3606 8120 3662 8129
rect 3804 8090 3832 8230
rect 3606 8055 3662 8064
rect 3792 8084 3844 8090
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3620 7426 3648 8055
rect 3792 8026 3844 8032
rect 3528 7398 3648 7426
rect 3528 4049 3556 7398
rect 3790 6896 3846 6905
rect 3790 6831 3846 6840
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3620 4758 3648 4966
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3514 4040 3570 4049
rect 3514 3975 3570 3984
rect 3804 3913 3832 6831
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5234 3924 6054
rect 3988 5778 4016 10474
rect 4080 7585 4108 10610
rect 4172 8022 4200 12038
rect 4264 11626 4292 12242
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4908 11257 4936 11630
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4894 11248 4950 11257
rect 4252 11212 4304 11218
rect 4894 11183 4950 11192
rect 4252 11154 4304 11160
rect 4264 10713 4292 11154
rect 4802 11112 4858 11121
rect 4712 11076 4764 11082
rect 4802 11047 4858 11056
rect 4712 11018 4764 11024
rect 4250 10704 4306 10713
rect 4250 10639 4252 10648
rect 4304 10639 4306 10648
rect 4252 10610 4304 10616
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4264 9217 4292 10066
rect 4540 9722 4568 10066
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4342 9344 4398 9353
rect 4342 9279 4398 9288
rect 4250 9208 4306 9217
rect 4250 9143 4306 9152
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4264 8634 4292 9046
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4172 7002 4200 7958
rect 4264 7546 4292 7958
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 7478 4384 9279
rect 4436 8968 4488 8974
rect 4434 8936 4436 8945
rect 4488 8936 4490 8945
rect 4434 8871 4490 8880
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4540 8634 4568 8842
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4526 7984 4582 7993
rect 4526 7919 4582 7928
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4540 7342 4568 7919
rect 4632 7410 4660 9998
rect 4724 8401 4752 11018
rect 4710 8392 4766 8401
rect 4710 8327 4766 8336
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4724 6780 4752 6870
rect 4816 6798 4844 11047
rect 4632 6752 4752 6780
rect 4804 6792 4856 6798
rect 4632 6390 4660 6752
rect 4804 6734 4856 6740
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4172 5846 4200 6122
rect 4632 6118 4660 6326
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5914 4660 6054
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3988 5409 4016 5714
rect 3974 5400 4030 5409
rect 4172 5370 4200 5782
rect 4816 5710 4844 6734
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 3974 5335 4030 5344
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 3896 4826 3924 5170
rect 4158 4856 4214 4865
rect 3884 4820 3936 4826
rect 4158 4791 4214 4800
rect 3884 4762 3936 4768
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3988 4282 4016 4694
rect 4172 4622 4200 4791
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 4724 4185 4752 5170
rect 4804 4616 4856 4622
rect 4802 4584 4804 4593
rect 4856 4584 4858 4593
rect 4802 4519 4858 4528
rect 4816 4214 4844 4519
rect 4804 4208 4856 4214
rect 4710 4176 4766 4185
rect 4252 4140 4304 4146
rect 4080 4100 4252 4128
rect 3790 3904 3846 3913
rect 3790 3839 3846 3848
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3712 3194 3740 3538
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 2964 3062 3016 3068
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 4080 2582 4108 4100
rect 4804 4150 4856 4156
rect 4710 4111 4712 4120
rect 4252 4082 4304 4088
rect 4764 4111 4766 4120
rect 4712 4082 4764 4088
rect 4724 4051 4752 4082
rect 4250 4040 4306 4049
rect 4250 3975 4252 3984
rect 4304 3975 4306 3984
rect 4252 3946 4304 3952
rect 4264 3670 4292 3946
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3194 4200 3538
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2650 4752 2926
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 3424 2304 3476 2310
rect 4908 2281 4936 11183
rect 5000 7410 5028 11494
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10606 5212 11154
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10470 5212 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10033 5212 10406
rect 5170 10024 5226 10033
rect 5170 9959 5226 9968
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5092 8498 5120 8910
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 8022 5120 8434
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5184 3738 5212 9454
rect 5276 6322 5304 12582
rect 5460 11801 5488 12582
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5446 11792 5502 11801
rect 5446 11727 5502 11736
rect 5448 11620 5500 11626
rect 5500 11580 5580 11608
rect 5448 11562 5500 11568
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 8906 5488 11018
rect 5552 10577 5580 11580
rect 5920 11558 5948 12242
rect 6182 11656 6238 11665
rect 6182 11591 6238 11600
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5816 10600 5868 10606
rect 5538 10568 5594 10577
rect 5816 10542 5868 10548
rect 5538 10503 5594 10512
rect 5722 10432 5778 10441
rect 5722 10367 5778 10376
rect 5736 10130 5764 10367
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5552 8537 5580 9862
rect 5736 9382 5764 10066
rect 5828 9586 5856 10542
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8634 5672 8978
rect 5736 8945 5764 9318
rect 5722 8936 5778 8945
rect 5722 8871 5778 8880
rect 5632 8628 5684 8634
rect 5684 8588 5764 8616
rect 5632 8570 5684 8576
rect 5538 8528 5594 8537
rect 5538 8463 5594 8472
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 7750 5396 8298
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 6866 5396 7210
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5846 5304 6258
rect 5368 6186 5396 6802
rect 5460 6458 5488 7890
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5552 6798 5580 7346
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5644 6730 5672 7346
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 5914 5396 6122
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5644 5642 5672 6666
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5538 5400 5594 5409
rect 5538 5335 5540 5344
rect 5592 5335 5594 5344
rect 5540 5306 5592 5312
rect 5736 4570 5764 8588
rect 5828 8566 5856 9522
rect 5920 9353 5948 11494
rect 6196 11218 6224 11591
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10470 6224 11154
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 5906 9344 5962 9353
rect 5906 9279 5962 9288
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5920 6633 5948 9279
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 8498 6040 8842
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5906 6624 5962 6633
rect 5906 6559 5962 6568
rect 5552 4542 5764 4570
rect 5264 3936 5316 3942
rect 5552 3913 5580 4542
rect 5722 4448 5778 4457
rect 5722 4383 5778 4392
rect 5264 3878 5316 3884
rect 5538 3904 5594 3913
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3126 5304 3878
rect 5538 3839 5594 3848
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5368 3641 5396 3674
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5092 2514 5120 2926
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 3424 2246 3476 2252
rect 4894 2272 4950 2281
rect 2778 504 2834 513
rect 1122 0 1178 480
rect 3436 480 3464 2246
rect 4894 2207 4950 2216
rect 5276 2009 5304 3062
rect 5368 2972 5396 3567
rect 5552 3210 5580 3839
rect 5736 3738 5764 4383
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5828 3602 5856 3946
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5460 3194 5580 3210
rect 5448 3188 5580 3194
rect 5500 3182 5580 3188
rect 5448 3130 5500 3136
rect 5828 2990 5856 3538
rect 5920 3534 5948 3878
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 6012 3074 6040 8434
rect 6104 4826 6132 8910
rect 6196 7041 6224 10406
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 6288 9042 6316 9386
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 7886 6316 8978
rect 6276 7880 6328 7886
rect 6274 7848 6276 7857
rect 6328 7848 6330 7857
rect 6274 7783 6330 7792
rect 6182 7032 6238 7041
rect 6182 6967 6238 6976
rect 6276 6928 6328 6934
rect 6182 6896 6238 6905
rect 6276 6870 6328 6876
rect 6182 6831 6238 6840
rect 6196 5710 6224 6831
rect 6288 6390 6316 6870
rect 6380 6798 6408 11018
rect 6656 10810 6684 15520
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11348 12306 11376 12650
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6458 10568 6514 10577
rect 6458 10503 6514 10512
rect 6472 7954 6500 10503
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9722 6684 10066
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6550 9072 6606 9081
rect 6550 9007 6606 9016
rect 6564 8809 6592 9007
rect 6550 8800 6606 8809
rect 6550 8735 6606 8744
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6472 7546 6500 7890
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6564 7426 6592 8735
rect 6472 7398 6592 7426
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 6458 6408 6734
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6288 5953 6316 6122
rect 6274 5944 6330 5953
rect 6274 5879 6330 5888
rect 6288 5846 6316 5879
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6196 5234 6224 5646
rect 6288 5370 6316 5782
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6104 4078 6132 4762
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6472 3942 6500 7398
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6564 6322 6592 6734
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6656 6225 6684 9658
rect 6748 6780 6776 12038
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11121 6960 11494
rect 6918 11112 6974 11121
rect 6918 11047 6974 11056
rect 7024 10985 7052 11630
rect 7102 11520 7158 11529
rect 7102 11455 7158 11464
rect 7116 11218 7144 11455
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7010 10976 7066 10985
rect 7010 10911 7066 10920
rect 7116 10810 7144 11154
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 8022 10976 8078 10985
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7194 10296 7250 10305
rect 6828 10260 6880 10266
rect 7194 10231 7250 10240
rect 6828 10202 6880 10208
rect 6840 8090 6868 10202
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9654 6960 10066
rect 7208 9897 7236 10231
rect 7194 9888 7250 9897
rect 7194 9823 7250 9832
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7102 9480 7158 9489
rect 7012 9444 7064 9450
rect 6932 9404 7012 9432
rect 6932 8838 6960 9404
rect 7102 9415 7158 9424
rect 7012 9386 7064 9392
rect 7116 9382 7144 9415
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7010 9208 7066 9217
rect 7208 9194 7236 9823
rect 7010 9143 7066 9152
rect 7116 9166 7236 9194
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8090 6960 8774
rect 7024 8401 7052 9143
rect 7010 8392 7066 8401
rect 7010 8327 7066 8336
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6918 7712 6974 7721
rect 6918 7647 6974 7656
rect 6932 7546 6960 7647
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6826 7440 6882 7449
rect 6826 7375 6828 7384
rect 6880 7375 6882 7384
rect 6828 7346 6880 7352
rect 6920 6792 6972 6798
rect 6748 6752 6920 6780
rect 6920 6734 6972 6740
rect 7010 6760 7066 6769
rect 7010 6695 7066 6704
rect 7024 6254 7052 6695
rect 7012 6248 7064 6254
rect 6642 6216 6698 6225
rect 7012 6190 7064 6196
rect 6642 6151 6698 6160
rect 6656 4690 6684 6151
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4690 6868 5102
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6656 4214 6684 4626
rect 6840 4282 6868 4626
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6840 3738 6868 4218
rect 6932 4049 6960 6054
rect 6918 4040 6974 4049
rect 6918 3975 6974 3984
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6288 3194 6316 3538
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6090 3088 6146 3097
rect 6012 3046 6090 3074
rect 6090 3023 6146 3032
rect 5448 2984 5500 2990
rect 5368 2944 5448 2972
rect 5368 2514 5396 2944
rect 5448 2926 5500 2932
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5920 2825 5948 2858
rect 5906 2816 5962 2825
rect 5906 2751 5962 2760
rect 6012 2650 6040 2926
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6104 2514 6132 3023
rect 6918 2952 6974 2961
rect 6918 2887 6974 2896
rect 6932 2854 6960 2887
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6918 2544 6974 2553
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6092 2508 6144 2514
rect 6918 2479 6920 2488
rect 6092 2450 6144 2456
rect 6972 2479 6974 2488
rect 6920 2450 6972 2456
rect 5262 2000 5318 2009
rect 5262 1935 5318 1944
rect 5828 480 5856 2450
rect 7024 1329 7052 6190
rect 7116 2990 7144 9166
rect 7300 8974 7328 10406
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7194 8664 7250 8673
rect 7194 8599 7250 8608
rect 7208 7478 7236 8599
rect 7300 8566 7328 8910
rect 7392 8634 7420 9046
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7378 8392 7434 8401
rect 7378 8327 7434 8336
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8022 7328 8230
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7300 7274 7328 7958
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 6662 7328 7210
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 5846 7328 6598
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5370 7236 5714
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7392 4978 7420 8327
rect 7484 6905 7512 10950
rect 7622 10908 7918 10928
rect 8022 10911 8078 10920
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 8036 10810 8064 10911
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8128 10690 8156 11630
rect 10060 11626 10088 12242
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 10428 11665 10456 12038
rect 10508 11688 10560 11694
rect 10414 11656 10470 11665
rect 10048 11620 10100 11626
rect 10508 11630 10560 11636
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 10414 11591 10470 11600
rect 10048 11562 10100 11568
rect 8206 11384 8262 11393
rect 8206 11319 8262 11328
rect 8220 11218 8248 11319
rect 8208 11212 8260 11218
rect 9772 11212 9824 11218
rect 8260 11172 8340 11200
rect 8208 11154 8260 11160
rect 8312 10810 8340 11172
rect 9772 11154 9824 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9600 10810 9628 11086
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 8298 10704 8354 10713
rect 8128 10662 8298 10690
rect 8298 10639 8354 10648
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 8220 9722 8248 10406
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 8974 7604 9522
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8036 8090 8064 8570
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 8312 7449 8340 9318
rect 8404 8906 8432 9454
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8298 7440 8354 7449
rect 8298 7375 8354 7384
rect 8024 6928 8076 6934
rect 7470 6896 7526 6905
rect 8312 6916 8340 7375
rect 8404 7206 8432 7890
rect 8392 7200 8444 7206
rect 8390 7168 8392 7177
rect 8484 7200 8536 7206
rect 8444 7168 8446 7177
rect 8484 7142 8536 7148
rect 8390 7103 8446 7112
rect 8024 6870 8076 6876
rect 8128 6888 8340 6916
rect 8390 6896 8446 6905
rect 7470 6831 7526 6840
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 5914 7512 6734
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8036 6186 8064 6870
rect 8128 6662 8156 6888
rect 8390 6831 8446 6840
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8220 6322 8248 6666
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5914 8340 6122
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8128 5098 8156 5782
rect 8312 5370 8340 5850
rect 8404 5574 8432 6831
rect 8496 5778 8524 7142
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 7300 4950 7420 4978
rect 7300 4010 7328 4950
rect 8128 4758 8156 5034
rect 8116 4752 8168 4758
rect 7838 4720 7894 4729
rect 8116 4694 8168 4700
rect 7838 4655 7840 4664
rect 7892 4655 7894 4664
rect 7840 4626 7892 4632
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4146 7512 4558
rect 7852 4468 7880 4626
rect 8128 4486 8156 4694
rect 8206 4584 8262 4593
rect 8206 4519 8262 4528
rect 8300 4548 8352 4554
rect 8220 4486 8248 4519
rect 8300 4490 8352 4496
rect 8116 4480 8168 4486
rect 7852 4440 8064 4468
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3777 7420 3878
rect 7378 3768 7434 3777
rect 7378 3703 7434 3712
rect 7760 3466 7788 3946
rect 8036 3738 8064 4440
rect 8116 4422 8168 4428
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8128 3942 8156 4422
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 8128 3194 8156 3606
rect 8220 3534 8248 4422
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8312 3380 8340 4490
rect 8220 3352 8340 3380
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8220 3074 8248 3352
rect 8036 3046 8248 3074
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 2582 7972 2926
rect 8036 2650 8064 3046
rect 8114 2952 8170 2961
rect 8114 2887 8170 2896
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 7010 1320 7066 1329
rect 7010 1255 7066 1264
rect 8128 480 8156 2887
rect 8588 2650 8616 10474
rect 9784 10470 9812 11154
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9048 10033 9076 10066
rect 9034 10024 9090 10033
rect 9034 9959 9090 9968
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8680 8634 8708 9454
rect 9048 9382 9076 9959
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 7750 8708 8366
rect 8772 8242 8800 8842
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8430 8892 8774
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8944 8288 8996 8294
rect 8772 8214 8892 8242
rect 8944 8230 8996 8236
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 7449 8708 7686
rect 8666 7440 8722 7449
rect 8666 7375 8722 7384
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8680 2446 8708 7375
rect 8864 7342 8892 8214
rect 8956 8090 8984 8230
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8772 6458 8800 7278
rect 8864 6662 8892 7278
rect 8852 6656 8904 6662
rect 8850 6624 8852 6633
rect 8904 6624 8906 6633
rect 8850 6559 8906 6568
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8864 4554 8892 6559
rect 9048 5817 9076 9318
rect 9034 5808 9090 5817
rect 9034 5743 9090 5752
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 9232 4282 9260 4694
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9034 4176 9090 4185
rect 9034 4111 9090 4120
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3670 8800 3878
rect 9048 3738 9076 4111
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8760 3528 8812 3534
rect 8758 3496 8760 3505
rect 8812 3496 8814 3505
rect 8758 3431 8814 3440
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 2922 8800 3334
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8864 2582 8892 2926
rect 9416 2689 9444 10406
rect 9784 10305 9812 10406
rect 9770 10296 9826 10305
rect 9770 10231 9826 10240
rect 9784 10130 9812 10231
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9600 8129 9628 9862
rect 9784 9722 9812 10066
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9876 7177 9904 11018
rect 10060 9081 10088 11562
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 11121 10456 11494
rect 10414 11112 10470 11121
rect 10414 11047 10470 11056
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10046 9072 10102 9081
rect 10046 9007 10048 9016
rect 10100 9007 10102 9016
rect 10140 9036 10192 9042
rect 10048 8978 10100 8984
rect 10140 8978 10192 8984
rect 10060 8566 10088 8978
rect 10152 8634 10180 8978
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10336 7993 10364 10542
rect 10520 9518 10548 11630
rect 11256 11257 11284 11630
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11242 11248 11298 11257
rect 11242 11183 11298 11192
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10508 9512 10560 9518
rect 10560 9472 10640 9500
rect 10508 9454 10560 9460
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10322 7984 10378 7993
rect 9956 7948 10008 7954
rect 10322 7919 10378 7928
rect 9956 7890 10008 7896
rect 9968 7313 9996 7890
rect 10520 7410 10548 9318
rect 10612 9217 10640 9472
rect 10598 9208 10654 9217
rect 10598 9143 10600 9152
rect 10652 9143 10654 9152
rect 10600 9114 10652 9120
rect 10612 9083 10640 9114
rect 10704 9081 10732 10406
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10690 9072 10746 9081
rect 10690 9007 10746 9016
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8090 10640 8910
rect 10690 8256 10746 8265
rect 10690 8191 10746 8200
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10704 7993 10732 8191
rect 10690 7984 10746 7993
rect 10690 7919 10746 7928
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 9954 7304 10010 7313
rect 9954 7239 10010 7248
rect 9968 7206 9996 7239
rect 9956 7200 10008 7206
rect 9862 7168 9918 7177
rect 9956 7142 10008 7148
rect 9862 7103 9918 7112
rect 9586 6896 9642 6905
rect 9586 6831 9588 6840
rect 9640 6831 9642 6840
rect 9588 6802 9640 6808
rect 9600 6458 9628 6802
rect 9968 6769 9996 7142
rect 10520 7002 10548 7346
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10796 6866 10824 10202
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 9042 10916 9454
rect 10980 9217 11008 11018
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10470 11284 10950
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 10966 9208 11022 9217
rect 10966 9143 11022 9152
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 8090 11008 8298
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 9954 6760 10010 6769
rect 9954 6695 10010 6704
rect 10138 6760 10194 6769
rect 10138 6695 10194 6704
rect 10152 6662 10180 6695
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5364 9640 5370
rect 9692 5352 9720 6054
rect 9640 5324 9720 5352
rect 9588 5306 9640 5312
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 4554 9628 5102
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4729 9720 4966
rect 9784 4865 9812 6598
rect 10152 6254 10180 6598
rect 10796 6458 10824 6802
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10140 6248 10192 6254
rect 10138 6216 10140 6225
rect 11256 6225 11284 10406
rect 11440 9178 11468 11494
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10130 11560 10610
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9722 11560 10066
rect 11716 9926 11744 11154
rect 11704 9920 11756 9926
rect 11702 9888 11704 9897
rect 11756 9888 11758 9897
rect 11702 9823 11758 9832
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11532 9518 11560 9658
rect 11808 9654 11836 12038
rect 12176 11558 12204 12242
rect 12164 11552 12216 11558
rect 11978 11520 12034 11529
rect 11978 11455 12034 11464
rect 12162 11520 12164 11529
rect 12716 11552 12768 11558
rect 12216 11520 12218 11529
rect 12716 11494 12768 11500
rect 12162 11455 12218 11464
rect 11992 11257 12020 11455
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 9897 11928 10542
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11886 9888 11942 9897
rect 11886 9823 11942 9832
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11808 9382 11836 9590
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11336 8492 11388 8498
rect 11440 8480 11468 9114
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11388 8452 11468 8480
rect 11336 8434 11388 8440
rect 11716 7886 11744 8910
rect 11900 8362 11928 9046
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11900 6866 11928 8298
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11992 7206 12020 7958
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 7002 12020 7142
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11992 6458 12020 6938
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11704 6384 11756 6390
rect 11334 6352 11390 6361
rect 11704 6326 11756 6332
rect 11334 6287 11390 6296
rect 10192 6216 10194 6225
rect 10048 6180 10100 6186
rect 10138 6151 10194 6160
rect 11242 6216 11298 6225
rect 11242 6151 11298 6160
rect 10048 6122 10100 6128
rect 10060 5710 10088 6122
rect 10048 5704 10100 5710
rect 10046 5672 10048 5681
rect 10100 5672 10102 5681
rect 10046 5607 10102 5616
rect 9954 5264 10010 5273
rect 9954 5199 10010 5208
rect 9968 5166 9996 5199
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9770 4856 9826 4865
rect 9770 4791 9826 4800
rect 9678 4720 9734 4729
rect 9678 4655 9734 4664
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9784 4185 9812 4558
rect 9770 4176 9826 4185
rect 9770 4111 9826 4120
rect 9586 4040 9642 4049
rect 9586 3975 9588 3984
rect 9640 3975 9642 3984
rect 9588 3946 9640 3952
rect 10152 3738 10180 6151
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10428 5370 10456 5782
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10520 4758 10548 5510
rect 11152 5160 11204 5166
rect 10598 5128 10654 5137
rect 11152 5102 11204 5108
rect 10598 5063 10654 5072
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10232 3936 10284 3942
rect 10230 3904 10232 3913
rect 10284 3904 10286 3913
rect 10230 3839 10286 3848
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9494 2816 9550 2825
rect 9692 2802 9720 3538
rect 10244 3194 10272 3839
rect 10520 3505 10548 4694
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 9550 2774 9720 2802
rect 9494 2751 9550 2760
rect 9402 2680 9458 2689
rect 9508 2650 9536 2751
rect 9402 2615 9458 2624
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9968 2582 9996 3130
rect 10520 2582 10548 3431
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 10612 1442 10640 5063
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10796 4010 10824 4422
rect 11164 4185 11192 5102
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11150 4176 11206 4185
rect 11150 4111 11206 4120
rect 11256 4049 11284 4558
rect 11348 4146 11376 6287
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11440 4146 11468 5510
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4729 11560 5034
rect 11716 5001 11744 6326
rect 11992 5846 12020 6394
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11992 5234 12020 5782
rect 12084 5710 12112 10474
rect 12452 10062 12480 11086
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9450 12572 9862
rect 12532 9444 12584 9450
rect 12360 9404 12532 9432
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8566 12296 8842
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12360 8090 12388 9404
rect 12532 9386 12584 9392
rect 12636 9178 12664 9998
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12530 9072 12586 9081
rect 12530 9007 12586 9016
rect 12544 8498 12572 9007
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12176 6118 12204 7278
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6322 12572 6598
rect 12636 6458 12664 8570
rect 12728 6798 12756 11494
rect 13188 10826 13216 12582
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13464 11558 13492 12242
rect 17038 12200 17094 12209
rect 17038 12135 17094 12144
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14016 11558 14044 12038
rect 14292 11694 14320 12038
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13188 10798 13308 10826
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12820 9722 12848 9930
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9382 12848 9522
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12912 8634 12940 10406
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12806 8120 12862 8129
rect 12806 8055 12862 8064
rect 12820 7886 12848 8055
rect 12912 8022 12940 8230
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7546 12848 7822
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 7478 12940 7958
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6934 12940 7142
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12360 6066 12388 6122
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11888 5024 11940 5030
rect 11702 4992 11758 5001
rect 11888 4966 11940 4972
rect 11702 4927 11758 4936
rect 11518 4720 11574 4729
rect 11518 4655 11574 4664
rect 11900 4593 11928 4966
rect 11992 4758 12020 5170
rect 12176 4826 12204 6054
rect 12360 6038 12480 6066
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11886 4584 11942 4593
rect 11886 4519 11942 4528
rect 11992 4282 12020 4694
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11242 4040 11298 4049
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 11060 4004 11112 4010
rect 11242 3975 11298 3984
rect 11060 3946 11112 3952
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10888 2650 10916 3606
rect 11072 3602 11100 3946
rect 11256 3738 11284 3975
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11348 3602 11376 4082
rect 12452 3738 12480 6038
rect 12544 5642 12572 6258
rect 12636 5914 12664 6258
rect 12728 5914 12756 6734
rect 12912 6458 12940 6870
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12532 5160 12584 5166
rect 12530 5128 12532 5137
rect 12584 5128 12586 5137
rect 12530 5063 12586 5072
rect 12636 4826 12664 5850
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12728 4706 12756 5238
rect 12820 4758 12848 6394
rect 13004 5370 13032 10542
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13004 5166 13032 5306
rect 13096 5302 13124 9658
rect 13188 9586 13216 9862
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13280 9382 13308 10798
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13266 9208 13322 9217
rect 13176 9172 13228 9178
rect 13266 9143 13322 9152
rect 13176 9114 13228 9120
rect 13188 7834 13216 9114
rect 13280 8974 13308 9143
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8566 13308 8910
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13188 7806 13308 7834
rect 13174 7712 13230 7721
rect 13174 7647 13230 7656
rect 13188 6798 13216 7647
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6390 13216 6734
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13082 5128 13138 5137
rect 13082 5063 13138 5072
rect 13096 4758 13124 5063
rect 12636 4678 12756 4706
rect 12808 4752 12860 4758
rect 13084 4752 13136 4758
rect 12860 4712 13032 4740
rect 12808 4694 12860 4700
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12162 3632 12218 3641
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11612 3596 11664 3602
rect 12162 3567 12218 3576
rect 11612 3538 11664 3544
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11072 2582 11100 3538
rect 11624 2922 11652 3538
rect 12176 3194 12204 3567
rect 12532 3392 12584 3398
rect 12636 3369 12664 4678
rect 13004 4049 13032 4712
rect 13084 4694 13136 4700
rect 12990 4040 13046 4049
rect 12808 4004 12860 4010
rect 12990 3975 13046 3984
rect 12808 3946 12860 3952
rect 12820 3670 12848 3946
rect 12808 3664 12860 3670
rect 12728 3612 12808 3618
rect 12728 3606 12860 3612
rect 12728 3590 12848 3606
rect 13004 3602 13032 3975
rect 13082 3768 13138 3777
rect 13082 3703 13138 3712
rect 12992 3596 13044 3602
rect 12532 3334 12584 3340
rect 12622 3360 12678 3369
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12176 2922 12204 3130
rect 12544 3126 12572 3334
rect 12622 3295 12678 3304
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12544 2961 12572 3062
rect 12530 2952 12586 2961
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 12164 2916 12216 2922
rect 12530 2887 12586 2896
rect 12164 2858 12216 2864
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 12636 2446 12664 3295
rect 12728 2650 12756 3590
rect 12992 3538 13044 3544
rect 12806 3496 12862 3505
rect 12806 3431 12862 3440
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 11888 2440 11940 2446
rect 11886 2408 11888 2417
rect 12624 2440 12676 2446
rect 11940 2408 11942 2417
rect 12624 2382 12676 2388
rect 11886 2343 11942 2352
rect 12820 2310 12848 3431
rect 13096 3058 13124 3703
rect 13280 3534 13308 7806
rect 13372 6633 13400 10950
rect 13464 10266 13492 11494
rect 14016 11218 14044 11494
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14016 10674 14044 11154
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13740 9654 13768 10066
rect 14108 9926 14136 10542
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13728 9648 13780 9654
rect 13648 9608 13728 9636
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8634 13492 9046
rect 13556 8974 13584 9386
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13556 7886 13584 8910
rect 13544 7880 13596 7886
rect 13450 7848 13506 7857
rect 13544 7822 13596 7828
rect 13450 7783 13506 7792
rect 13358 6624 13414 6633
rect 13358 6559 13414 6568
rect 13464 5760 13492 7783
rect 13464 5732 13584 5760
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13464 4622 13492 5578
rect 13556 4758 13584 5732
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13556 3641 13584 4014
rect 13648 3670 13676 9608
rect 13728 9590 13780 9596
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 7857 13768 8434
rect 13726 7848 13782 7857
rect 13726 7783 13782 7792
rect 13832 6361 13860 9318
rect 13818 6352 13874 6361
rect 13818 6287 13874 6296
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 5228 13780 5234
rect 13832 5216 13860 5510
rect 13780 5188 13860 5216
rect 13728 5170 13780 5176
rect 13740 3942 13768 5170
rect 13818 4992 13874 5001
rect 13818 4927 13874 4936
rect 13832 4078 13860 4927
rect 13924 4282 13952 9522
rect 14108 7449 14136 9862
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14660 8498 14688 9454
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14094 7440 14150 7449
rect 14094 7375 14150 7384
rect 14554 7440 14610 7449
rect 14554 7375 14610 7384
rect 14568 7342 14596 7375
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14094 7168 14150 7177
rect 14094 7103 14150 7112
rect 14108 7002 14136 7103
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14016 5846 14044 6122
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14660 5914 14688 8298
rect 14752 7313 14780 8366
rect 14738 7304 14794 7313
rect 14738 7239 14794 7248
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 7002 14780 7142
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14844 6769 14872 11698
rect 15290 11656 15346 11665
rect 15016 11620 15068 11626
rect 15290 11591 15346 11600
rect 15016 11562 15068 11568
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14936 8498 14964 11086
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14830 6760 14886 6769
rect 14830 6695 14886 6704
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14016 4826 14044 5782
rect 14660 5137 14688 5850
rect 14844 5778 14872 6695
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14646 5128 14702 5137
rect 14646 5063 14702 5072
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13924 3738 13952 4218
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13636 3664 13688 3670
rect 13542 3632 13598 3641
rect 13636 3606 13688 3612
rect 13542 3567 13598 3576
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13280 3194 13308 3470
rect 13924 3466 13952 3674
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 14016 2990 14044 3334
rect 14004 2984 14056 2990
rect 14108 2961 14136 3470
rect 14200 2990 14228 4694
rect 14738 4584 14794 4593
rect 14738 4519 14794 4528
rect 14752 4146 14780 4519
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14936 3942 14964 8298
rect 15028 7970 15056 11562
rect 15304 10810 15332 11591
rect 17052 11354 17080 12135
rect 18326 11792 18382 11801
rect 18326 11727 18382 11736
rect 18340 11694 18368 11727
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 17130 11384 17186 11393
rect 17040 11348 17092 11354
rect 17130 11319 17186 11328
rect 17040 11290 17092 11296
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 15660 11144 15712 11150
rect 15382 11112 15438 11121
rect 15660 11086 15712 11092
rect 15382 11047 15438 11056
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15304 10606 15332 10746
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15120 9058 15148 10474
rect 15396 10130 15424 11047
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 9722 15424 10066
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15292 9648 15344 9654
rect 15396 9625 15424 9658
rect 15292 9590 15344 9596
rect 15382 9616 15438 9625
rect 15120 9042 15240 9058
rect 15120 9036 15252 9042
rect 15120 9030 15200 9036
rect 15120 8090 15148 9030
rect 15200 8978 15252 8984
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15028 7954 15240 7970
rect 15028 7948 15252 7954
rect 15028 7942 15200 7948
rect 15200 7890 15252 7896
rect 15212 7002 15240 7890
rect 15304 7410 15332 9590
rect 15672 9586 15700 11086
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 15382 9551 15438 9560
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 9178 16160 9386
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15396 8566 15424 9046
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15396 8362 15424 8502
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15396 8090 15424 8298
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15396 7546 15424 8026
rect 15750 7576 15806 7585
rect 15384 7540 15436 7546
rect 15750 7511 15806 7520
rect 15384 7482 15436 7488
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15212 5370 15240 5714
rect 15304 5710 15332 7210
rect 15764 6866 15792 7511
rect 16132 7274 16160 8230
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15396 5137 15424 5170
rect 15382 5128 15438 5137
rect 15382 5063 15384 5072
rect 15436 5063 15438 5072
rect 15384 5034 15436 5040
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 4264 15148 4422
rect 15120 4236 15240 4264
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14936 3505 14964 3878
rect 15120 3738 15148 4014
rect 15212 4010 15240 4236
rect 15304 4146 15332 4626
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15016 3528 15068 3534
rect 14922 3496 14978 3505
rect 15016 3470 15068 3476
rect 14922 3431 14978 3440
rect 14188 2984 14240 2990
rect 14004 2926 14056 2932
rect 14094 2952 14150 2961
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13266 2680 13322 2689
rect 13266 2615 13268 2624
rect 13320 2615 13322 2624
rect 13268 2586 13320 2592
rect 12900 2576 12952 2582
rect 13924 2553 13952 2790
rect 14016 2650 14044 2926
rect 14188 2926 14240 2932
rect 14094 2887 14150 2896
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 12900 2518 12952 2524
rect 13910 2544 13966 2553
rect 12808 2304 12860 2310
rect 12912 2281 12940 2518
rect 14108 2514 14136 2887
rect 15028 2854 15056 3470
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 13910 2479 13966 2488
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 15028 2378 15056 2790
rect 15120 2632 15148 3130
rect 15200 2644 15252 2650
rect 15120 2604 15200 2632
rect 15200 2586 15252 2592
rect 15304 2530 15332 4082
rect 15488 3641 15516 6598
rect 15764 6118 15792 6802
rect 16224 6798 16252 10406
rect 16316 10130 16344 10542
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16316 9654 16344 10066
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16316 9489 16344 9590
rect 16302 9480 16358 9489
rect 16302 9415 16358 9424
rect 16408 6866 16436 9998
rect 16500 9353 16528 10474
rect 16684 10470 16712 11154
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 9450 16712 10406
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16486 9344 16542 9353
rect 16486 9279 16542 9288
rect 16684 8906 16712 9386
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16500 8090 16528 8230
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16488 7880 16540 7886
rect 16486 7848 16488 7857
rect 16540 7848 16542 7857
rect 16486 7783 16542 7792
rect 16500 7410 16528 7783
rect 16684 7410 16712 8842
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16868 7750 16896 8366
rect 16856 7744 16908 7750
rect 16854 7712 16856 7721
rect 16908 7712 16910 7721
rect 16854 7647 16910 7656
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16960 6934 16988 8502
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6458 16252 6734
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16408 6322 16436 6802
rect 16854 6624 16910 6633
rect 16854 6559 16910 6568
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 15752 6112 15804 6118
rect 15566 6080 15622 6089
rect 15752 6054 15804 6060
rect 15566 6015 15622 6024
rect 15580 5914 15608 6015
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15658 5672 15714 5681
rect 15658 5607 15714 5616
rect 15672 5234 15700 5607
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15764 4593 15792 6054
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15856 5098 15884 5510
rect 16408 5370 16436 5782
rect 16868 5574 16896 6559
rect 16960 6186 16988 6870
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16960 5846 16988 6122
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16856 5568 16908 5574
rect 17052 5545 17080 9318
rect 17144 8634 17172 11319
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17682 9480 17738 9489
rect 17682 9415 17738 9424
rect 17696 9382 17724 9415
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17236 8362 17264 9046
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17144 7206 17172 7958
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17512 7546 17540 7822
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17144 6662 17172 7142
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 16856 5510 16908 5516
rect 17038 5536 17094 5545
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16868 5166 16896 5510
rect 17038 5471 17094 5480
rect 17052 5370 17080 5471
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 16948 5024 17000 5030
rect 16394 4992 16450 5001
rect 16948 4966 17000 4972
rect 16394 4927 16450 4936
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15750 4584 15806 4593
rect 15750 4519 15806 4528
rect 15856 3738 15884 4626
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4146 16344 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15474 3632 15530 3641
rect 15474 3567 15530 3576
rect 15580 2553 15608 3674
rect 15752 3392 15804 3398
rect 15750 3360 15752 3369
rect 15804 3360 15806 3369
rect 15750 3295 15806 3304
rect 15764 3194 15792 3295
rect 16316 3194 16344 4082
rect 16408 3670 16436 4927
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16500 3602 16528 3946
rect 16592 3942 16620 4150
rect 16684 4146 16712 4558
rect 16960 4486 16988 4966
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17144 4214 17172 4422
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16026 3088 16082 3097
rect 16500 3074 16528 3538
rect 16684 3534 16712 4082
rect 16946 4040 17002 4049
rect 16946 3975 17002 3984
rect 17040 4004 17092 4010
rect 16960 3602 16988 3975
rect 17040 3946 17092 3952
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16578 3088 16634 3097
rect 16500 3046 16578 3074
rect 16026 3023 16028 3032
rect 16080 3023 16082 3032
rect 16578 3023 16634 3032
rect 16028 2994 16080 3000
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15212 2502 15332 2530
rect 15566 2544 15622 2553
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14832 2304 14884 2310
rect 12808 2246 12860 2252
rect 12898 2272 12954 2281
rect 10520 1414 10640 1442
rect 10520 480 10548 1414
rect 12820 480 12848 2246
rect 14832 2246 14884 2252
rect 12898 2207 12954 2216
rect 14844 2009 14872 2246
rect 14830 2000 14886 2009
rect 14830 1935 14886 1944
rect 15212 480 15240 2502
rect 15566 2479 15622 2488
rect 15672 2446 15700 2926
rect 16592 2650 16620 3023
rect 17052 2689 17080 3946
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17144 3194 17172 3470
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17038 2680 17094 2689
rect 16580 2644 16632 2650
rect 17328 2650 17356 4422
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17512 2650 17540 3606
rect 17604 3194 17632 4150
rect 17696 3482 17724 9318
rect 17880 7886 17908 10406
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17972 9722 18000 10066
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17958 9616 18014 9625
rect 17958 9551 18014 9560
rect 17972 9518 18000 9551
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17972 9178 18000 9454
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17972 9081 18000 9114
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 18064 8945 18092 10542
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18248 9450 18276 10066
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18234 9344 18290 9353
rect 18050 8936 18106 8945
rect 18050 8871 18106 8880
rect 17960 8560 18012 8566
rect 18064 8537 18092 8871
rect 17960 8502 18012 8508
rect 18050 8528 18106 8537
rect 17972 8022 18000 8502
rect 18050 8463 18106 8472
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 18156 7410 18184 9318
rect 18234 9279 18290 9288
rect 18248 9042 18276 9279
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17880 6934 17908 7210
rect 18156 7002 18184 7346
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17880 6186 17908 6598
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 18236 5296 18288 5302
rect 18234 5264 18236 5273
rect 18288 5264 18290 5273
rect 18234 5199 18290 5208
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17776 5024 17828 5030
rect 18064 5001 18092 5102
rect 17776 4966 17828 4972
rect 18050 4992 18106 5001
rect 17788 4865 17816 4966
rect 18050 4927 18106 4936
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 17788 4690 17816 4791
rect 18340 4690 18368 9998
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 17788 4010 17816 4626
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 18064 4282 18092 4490
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18050 4176 18106 4185
rect 18050 4111 18106 4120
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17788 3670 17816 3946
rect 17866 3768 17922 3777
rect 17866 3703 17868 3712
rect 17920 3703 17922 3712
rect 17868 3674 17920 3680
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17696 3454 17816 3482
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17788 2922 17816 3454
rect 17972 2990 18000 3538
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17038 2615 17094 2624
rect 17316 2644 17368 2650
rect 16580 2586 16632 2592
rect 17316 2586 17368 2592
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 17604 480 17632 2586
rect 17788 2378 17816 2858
rect 18064 2650 18092 4111
rect 18248 4078 18276 4422
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18248 3466 18276 4014
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18432 3058 18460 12582
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18510 11248 18566 11257
rect 18510 11183 18512 11192
rect 18564 11183 18566 11192
rect 18512 11154 18564 11160
rect 18524 10810 18552 11154
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18524 9110 18552 9454
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18524 8634 18552 9046
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 7750 18552 8298
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18616 6730 18644 11018
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18708 7954 18736 9114
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7002 18736 7890
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18800 6798 18828 11494
rect 19338 10840 19394 10849
rect 19338 10775 19394 10784
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18984 9761 19012 10542
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18970 9752 19026 9761
rect 18970 9687 19026 9696
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 6934 18920 7686
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18616 6168 18644 6666
rect 18800 6390 18828 6734
rect 18892 6458 18920 6870
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18788 6180 18840 6186
rect 18616 6140 18788 6168
rect 18788 6122 18840 6128
rect 18984 5710 19012 8502
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 19076 5642 19104 10406
rect 19352 10130 19380 10775
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19352 9722 19380 10066
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19260 8634 19288 8910
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19352 8537 19380 8910
rect 19338 8528 19394 8537
rect 19338 8463 19394 8472
rect 19260 8362 19380 8378
rect 19260 8356 19392 8362
rect 19260 8350 19340 8356
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 19168 7206 19196 7958
rect 19260 7546 19288 8350
rect 19340 8298 19392 8304
rect 19444 8242 19472 11630
rect 19996 11393 20024 15520
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 33336 12209 33364 15520
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35440 12776 35492 12782
rect 35440 12718 35492 12724
rect 33322 12200 33378 12209
rect 33322 12135 33378 12144
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 20718 11792 20774 11801
rect 20718 11727 20774 11736
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19982 11384 20038 11393
rect 19982 11319 20038 11328
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19536 10713 19564 11154
rect 20088 11121 20116 11494
rect 20074 11112 20130 11121
rect 19616 11076 19668 11082
rect 20074 11047 20130 11056
rect 19616 11018 19668 11024
rect 19522 10704 19578 10713
rect 19522 10639 19524 10648
rect 19576 10639 19578 10648
rect 19524 10610 19576 10616
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19536 8838 19564 9454
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19352 8214 19472 8242
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 19076 5273 19104 5578
rect 19062 5264 19118 5273
rect 19062 5199 19118 5208
rect 19168 5166 19196 7142
rect 19352 5681 19380 8214
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6186 19472 6734
rect 19628 6458 19656 11018
rect 20626 10976 20682 10985
rect 20626 10911 20682 10920
rect 19798 10704 19854 10713
rect 19798 10639 19854 10648
rect 19708 9920 19760 9926
rect 19812 9897 19840 10639
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19892 9920 19944 9926
rect 19708 9862 19760 9868
rect 19798 9888 19854 9897
rect 19720 8498 19748 9862
rect 19892 9862 19944 9868
rect 19798 9823 19854 9832
rect 19904 9518 19932 9862
rect 19892 9512 19944 9518
rect 19812 9472 19892 9500
rect 19812 9042 19840 9472
rect 19892 9454 19944 9460
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19720 8090 19748 8434
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19812 7313 19840 8774
rect 19904 7410 19932 9318
rect 19996 8945 20024 10542
rect 20640 9994 20668 10911
rect 20732 10606 20760 11727
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 25502 11248 25558 11257
rect 22100 11212 22152 11218
rect 25502 11183 25558 11192
rect 26608 11212 26660 11218
rect 22100 11154 22152 11160
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 22112 10538 22140 11154
rect 22282 11112 22338 11121
rect 22282 11047 22338 11056
rect 24308 11076 24360 11082
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 22100 10532 22152 10538
rect 22100 10474 22152 10480
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19982 8936 20038 8945
rect 19982 8871 20038 8880
rect 20088 8498 20116 9114
rect 20548 8498 20576 9522
rect 20628 9172 20680 9178
rect 20732 9160 20760 10406
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 20824 9722 20852 9998
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20824 9625 20852 9658
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20680 9132 20760 9160
rect 20628 9114 20680 9120
rect 21284 9110 21312 9862
rect 21468 9450 21496 9862
rect 21560 9450 21588 9998
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21468 9353 21496 9386
rect 21454 9344 21510 9353
rect 21454 9279 21510 9288
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21364 9104 21416 9110
rect 21364 9046 21416 9052
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20732 7954 20760 8298
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19798 7304 19854 7313
rect 19798 7239 19854 7248
rect 19904 7002 19932 7346
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 20640 6934 20668 7210
rect 20824 7002 20852 8978
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21284 8634 21312 9046
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21376 8514 21404 9046
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21284 8486 21404 8514
rect 21468 8498 21496 8774
rect 21456 8492 21508 8498
rect 21284 8430 21312 8486
rect 21456 8434 21508 8440
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21560 8362 21588 9386
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21284 7546 21312 7958
rect 21652 7886 21680 9930
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 20088 6390 20116 6802
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21284 6458 21312 6802
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 20076 6384 20128 6390
rect 20074 6352 20076 6361
rect 20128 6352 20130 6361
rect 20074 6287 20130 6296
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19338 5672 19394 5681
rect 19338 5607 19394 5616
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19720 5166 19748 5510
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19168 4758 19196 5102
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 18788 4072 18840 4078
rect 18786 4040 18788 4049
rect 18840 4040 18842 4049
rect 19168 4010 19196 4694
rect 18786 3975 18842 3984
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19062 3632 19118 3641
rect 19062 3567 19064 3576
rect 19116 3567 19118 3576
rect 19616 3596 19668 3602
rect 19064 3538 19116 3544
rect 19616 3538 19668 3544
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18616 2990 18644 3334
rect 18328 2984 18380 2990
rect 18326 2952 18328 2961
rect 18604 2984 18656 2990
rect 18380 2952 18382 2961
rect 18604 2926 18656 2932
rect 19628 2922 19656 3538
rect 18326 2887 18382 2896
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19720 2854 19748 5102
rect 19892 4752 19944 4758
rect 19890 4720 19892 4729
rect 19944 4720 19946 4729
rect 19946 4678 20024 4706
rect 19890 4655 19946 4664
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 3482 19840 3878
rect 19904 3670 19932 4082
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19812 3454 19932 3482
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19812 2650 19840 2926
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 18328 2576 18380 2582
rect 18326 2544 18328 2553
rect 18380 2544 18382 2553
rect 18326 2479 18382 2488
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 19904 480 19932 3454
rect 19996 2514 20024 4678
rect 20088 3602 20116 6287
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 20456 5846 20484 6122
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4826 20576 4966
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20640 4146 20668 5510
rect 20732 5234 20760 5646
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20824 5030 20852 5782
rect 21008 5710 21036 6122
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 21284 4865 21312 6394
rect 21638 6352 21694 6361
rect 21638 6287 21694 6296
rect 21652 6118 21680 6287
rect 21640 6112 21692 6118
rect 21638 6080 21640 6089
rect 21692 6080 21694 6089
rect 21638 6015 21694 6024
rect 21270 4856 21326 4865
rect 21270 4791 21326 4800
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20824 4282 20852 4694
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21284 4282 21312 4558
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 2582 20668 3470
rect 20824 3194 20852 3538
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 21284 3194 21312 3606
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21284 3097 21312 3130
rect 21270 3088 21326 3097
rect 21270 3023 21326 3032
rect 20902 2680 20958 2689
rect 21376 2650 21404 4218
rect 21652 3194 21680 6015
rect 21744 5846 21772 10474
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 21836 9178 21864 10406
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8498 21864 8842
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21836 8129 21864 8434
rect 21822 8120 21878 8129
rect 21822 8055 21878 8064
rect 21836 8022 21864 8055
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21928 7478 21956 9522
rect 22020 8090 22048 10406
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 22020 7410 22048 8026
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22112 7290 22140 9386
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22020 7262 22140 7290
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 21836 6225 21864 6326
rect 21928 6254 21956 6938
rect 22020 6866 22048 7262
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 22204 6746 22232 9114
rect 22020 6718 22232 6746
rect 21916 6248 21968 6254
rect 21822 6216 21878 6225
rect 21916 6190 21968 6196
rect 21822 6151 21878 6160
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21744 5234 21772 5782
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21744 4758 21772 5170
rect 21928 4826 21956 5646
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21836 3398 21864 4014
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 20902 2615 20904 2624
rect 20956 2615 20958 2624
rect 21364 2644 21416 2650
rect 20904 2586 20956 2592
rect 21364 2586 21416 2592
rect 20628 2576 20680 2582
rect 20626 2544 20628 2553
rect 21836 2553 21864 3334
rect 22020 3097 22048 6718
rect 22296 6338 22324 11047
rect 24308 11018 24360 11024
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22388 10470 22416 10542
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22388 9897 22416 10406
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22374 9888 22430 9897
rect 22374 9823 22430 9832
rect 22480 9518 22508 9998
rect 22468 9512 22520 9518
rect 22466 9480 22468 9489
rect 22520 9480 22522 9489
rect 22940 9450 22968 10066
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 22466 9415 22522 9424
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 23478 9344 23534 9353
rect 23478 9279 23534 9288
rect 23492 9178 23520 9279
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22848 8809 22876 8978
rect 22834 8800 22890 8809
rect 22834 8735 22890 8744
rect 22848 8634 22876 8735
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22480 7478 22508 7822
rect 22468 7472 22520 7478
rect 22468 7414 22520 7420
rect 22480 7274 22508 7414
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22480 7002 22508 7210
rect 22848 7206 22876 7958
rect 23584 7750 23612 8502
rect 23662 8120 23718 8129
rect 23662 8055 23664 8064
rect 23716 8055 23718 8064
rect 23664 8026 23716 8032
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22848 6905 22876 7142
rect 23492 6934 23520 7142
rect 23480 6928 23532 6934
rect 22650 6896 22706 6905
rect 22650 6831 22706 6840
rect 22834 6896 22890 6905
rect 23480 6870 23532 6876
rect 22834 6831 22890 6840
rect 22928 6860 22980 6866
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22204 6310 22324 6338
rect 22388 6322 22416 6734
rect 22376 6316 22428 6322
rect 22100 5296 22152 5302
rect 22098 5264 22100 5273
rect 22152 5264 22154 5273
rect 22098 5199 22154 5208
rect 22204 4162 22232 6310
rect 22376 6258 22428 6264
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22296 5846 22324 6190
rect 22388 5914 22416 6258
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 22296 5370 22324 5782
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22296 4282 22324 5306
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22572 4622 22600 4966
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22664 4486 22692 6831
rect 22928 6802 22980 6808
rect 22940 6322 22968 6802
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23124 5710 23152 6054
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23124 5545 23152 5646
rect 23110 5536 23166 5545
rect 23110 5471 23166 5480
rect 23124 5030 23152 5471
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 23124 4729 23152 4966
rect 23584 4826 23612 7686
rect 23676 7478 23704 8026
rect 23664 7472 23716 7478
rect 23664 7414 23716 7420
rect 23572 4820 23624 4826
rect 23492 4780 23572 4808
rect 23110 4720 23166 4729
rect 23110 4655 23166 4664
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 23492 4282 23520 4780
rect 23572 4762 23624 4768
rect 23570 4720 23626 4729
rect 23768 4690 23796 9862
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23938 9208 23994 9217
rect 23938 9143 23994 9152
rect 23952 9042 23980 9143
rect 24044 9081 24072 9386
rect 24030 9072 24086 9081
rect 23940 9036 23992 9042
rect 24030 9007 24086 9016
rect 23940 8978 23992 8984
rect 23952 8634 23980 8978
rect 24136 8838 24164 10066
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24044 7410 24072 7822
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23860 5846 23888 6598
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23952 5914 23980 6190
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24044 4758 24072 5646
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 23570 4655 23626 4664
rect 23756 4684 23808 4690
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 22112 4134 22232 4162
rect 22006 3088 22062 3097
rect 22006 3023 22062 3032
rect 20680 2544 20682 2553
rect 19984 2508 20036 2514
rect 20626 2479 20682 2488
rect 21822 2544 21878 2553
rect 21822 2479 21878 2488
rect 19984 2450 20036 2456
rect 20076 2304 20128 2310
rect 20074 2272 20076 2281
rect 20128 2272 20130 2281
rect 20074 2207 20130 2216
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 22112 610 22140 4134
rect 22192 4072 22244 4078
rect 22296 4060 22324 4218
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 22244 4032 22324 4060
rect 22192 4014 22244 4020
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22204 3738 22232 3878
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 22742 3360 22798 3369
rect 22742 3295 22798 3304
rect 22756 3058 22784 3295
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23124 2922 23152 3606
rect 23400 2990 23428 4082
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23492 3194 23520 3674
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23112 2916 23164 2922
rect 23112 2858 23164 2864
rect 23400 2650 23428 2926
rect 23584 2650 23612 4655
rect 23756 4626 23808 4632
rect 23768 4214 23796 4626
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 24136 3777 24164 8774
rect 24320 5250 24348 11018
rect 25516 10849 25544 11183
rect 26608 11154 26660 11160
rect 34152 11212 34204 11218
rect 34152 11154 34204 11160
rect 35256 11212 35308 11218
rect 35256 11154 35308 11160
rect 26238 10976 26294 10985
rect 26238 10911 26294 10920
rect 25502 10840 25558 10849
rect 26252 10810 26280 10911
rect 25502 10775 25558 10784
rect 26240 10804 26292 10810
rect 25516 10130 25544 10775
rect 26240 10746 26292 10752
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 26148 10600 26200 10606
rect 26620 10577 26648 11154
rect 27526 11112 27582 11121
rect 27526 11047 27528 11056
rect 27580 11047 27582 11056
rect 29366 11112 29422 11121
rect 29366 11047 29422 11056
rect 27528 11018 27580 11024
rect 27158 10704 27214 10713
rect 27158 10639 27214 10648
rect 27172 10606 27200 10639
rect 26700 10600 26752 10606
rect 26148 10542 26200 10548
rect 26606 10568 26662 10577
rect 25700 10169 25728 10542
rect 25686 10160 25742 10169
rect 25504 10124 25556 10130
rect 25686 10095 25742 10104
rect 25504 10066 25556 10072
rect 24492 9920 24544 9926
rect 24492 9862 24544 9868
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24504 9518 24532 9862
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24596 9110 24624 9862
rect 25516 9722 25544 10066
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24412 7750 24440 8366
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24412 7585 24440 7686
rect 24398 7576 24454 7585
rect 24398 7511 24454 7520
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24398 6216 24454 6225
rect 24398 6151 24400 6160
rect 24452 6151 24454 6160
rect 24400 6122 24452 6128
rect 24320 5222 24434 5250
rect 24406 5216 24434 5222
rect 24406 5188 24440 5216
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 24320 4826 24348 5102
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 24122 3768 24178 3777
rect 24122 3703 24178 3712
rect 24228 3670 24256 3878
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24032 3528 24084 3534
rect 24030 3496 24032 3505
rect 24084 3496 24086 3505
rect 24030 3431 24086 3440
rect 24228 3194 24256 3606
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24412 2836 24440 5188
rect 24504 3534 24532 7346
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24688 6322 24716 6802
rect 24780 6338 24808 9522
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24872 9042 24900 9386
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24964 8430 24992 8978
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24872 7313 24900 7890
rect 24964 7886 24992 8366
rect 25424 8362 25452 8910
rect 25412 8356 25464 8362
rect 25412 8298 25464 8304
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24858 7304 24914 7313
rect 24858 7239 24860 7248
rect 24912 7239 24914 7248
rect 24860 7210 24912 7216
rect 24872 6474 24900 7210
rect 25332 7206 25360 7890
rect 25424 7857 25452 8298
rect 25410 7848 25466 7857
rect 25410 7783 25466 7792
rect 25608 7410 25636 8910
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25884 8090 25912 8366
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25976 7449 26004 9862
rect 25962 7440 26018 7449
rect 25596 7404 25648 7410
rect 25962 7375 26018 7384
rect 26056 7404 26108 7410
rect 25596 7346 25648 7352
rect 26056 7346 26108 7352
rect 25964 7268 26016 7274
rect 25964 7210 26016 7216
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 24950 6896 25006 6905
rect 24950 6831 24952 6840
rect 25004 6831 25006 6840
rect 24952 6802 25004 6808
rect 24950 6488 25006 6497
rect 24872 6446 24950 6474
rect 24950 6423 25006 6432
rect 24780 6322 24900 6338
rect 24676 6316 24728 6322
rect 24780 6316 24912 6322
rect 24780 6310 24860 6316
rect 24676 6258 24728 6264
rect 24860 6258 24912 6264
rect 24688 6186 24716 6258
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24872 5846 24900 6122
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 24872 5370 24900 5782
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24872 5098 24900 5306
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24584 5024 24636 5030
rect 24582 4992 24584 5001
rect 24636 4992 24638 5001
rect 24582 4927 24638 4936
rect 24964 4690 24992 6423
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 25240 5914 25268 6258
rect 25332 6254 25360 7142
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25332 5681 25360 6190
rect 25976 6186 26004 7210
rect 26068 7002 26096 7346
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 25964 6180 26016 6186
rect 25964 6122 26016 6128
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 25318 5672 25374 5681
rect 25318 5607 25374 5616
rect 26068 5302 26096 6054
rect 26160 5692 26188 10542
rect 26700 10542 26752 10548
rect 27160 10600 27212 10606
rect 28172 10600 28224 10606
rect 27160 10542 27212 10548
rect 28170 10568 28172 10577
rect 28224 10568 28226 10577
rect 26606 10503 26662 10512
rect 26620 10470 26648 10503
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26620 9654 26648 10406
rect 26712 10033 26740 10542
rect 27988 10532 28040 10538
rect 28170 10503 28226 10512
rect 27988 10474 28040 10480
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 27264 10266 27292 10406
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 26698 10024 26754 10033
rect 26698 9959 26754 9968
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 27264 9586 27292 10202
rect 27436 10192 27488 10198
rect 27436 10134 27488 10140
rect 27252 9580 27304 9586
rect 27252 9522 27304 9528
rect 26240 9512 26292 9518
rect 26238 9480 26240 9489
rect 26292 9480 26294 9489
rect 27448 9450 27476 10134
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 26238 9415 26294 9424
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26712 9178 26740 9318
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26804 8022 26832 8230
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26804 7274 26832 7958
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26804 6390 26832 6802
rect 26896 6769 26924 9318
rect 26976 9104 27028 9110
rect 26976 9046 27028 9052
rect 26988 8294 27016 9046
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26988 7546 27016 8230
rect 27448 8090 27476 9386
rect 27540 8838 27568 9998
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 28000 9110 28028 10474
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28262 9480 28318 9489
rect 28080 9444 28132 9450
rect 28262 9415 28318 9424
rect 28080 9386 28132 9392
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 27988 9104 28040 9110
rect 27988 9046 28040 9052
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27632 8838 27660 8910
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27434 7712 27490 7721
rect 27434 7647 27490 7656
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 27448 6866 27476 7647
rect 27540 7478 27568 8774
rect 27724 8498 27752 9046
rect 28092 8974 28120 9386
rect 28276 9217 28304 9415
rect 28262 9208 28318 9217
rect 28262 9143 28318 9152
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28080 8832 28132 8838
rect 28080 8774 28132 8780
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27816 8362 27844 8570
rect 27804 8356 27856 8362
rect 27804 8298 27856 8304
rect 27988 8356 28040 8362
rect 27988 8298 28040 8304
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 28000 8090 28028 8298
rect 28092 8090 28120 8774
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27632 7546 27660 7822
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 28170 7440 28226 7449
rect 28170 7375 28226 7384
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27540 6866 27568 7142
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 27804 6792 27856 6798
rect 26882 6760 26938 6769
rect 27804 6734 27856 6740
rect 26882 6695 26938 6704
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 26792 6384 26844 6390
rect 26792 6326 26844 6332
rect 27080 6186 27108 6598
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 27068 6180 27120 6186
rect 27068 6122 27120 6128
rect 26884 6112 26936 6118
rect 26884 6054 26936 6060
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 26240 5704 26292 5710
rect 26160 5664 26240 5692
rect 26240 5646 26292 5652
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 26252 5250 26280 5646
rect 26344 5642 26372 5782
rect 26332 5636 26384 5642
rect 26332 5578 26384 5584
rect 26344 5370 26372 5578
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26252 5222 26372 5250
rect 25410 5128 25466 5137
rect 25410 5063 25412 5072
rect 25464 5063 25466 5072
rect 25412 5034 25464 5040
rect 26344 4826 26372 5222
rect 26896 5001 26924 6054
rect 26974 5264 27030 5273
rect 26974 5199 26976 5208
rect 27028 5199 27030 5208
rect 26976 5170 27028 5176
rect 26882 4992 26938 5001
rect 26882 4927 26938 4936
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24964 4214 24992 4626
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 26148 4616 26200 4622
rect 26148 4558 26200 4564
rect 24952 4208 25004 4214
rect 24952 4150 25004 4156
rect 25044 4004 25096 4010
rect 25044 3946 25096 3952
rect 24674 3904 24730 3913
rect 24674 3839 24730 3848
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24412 2808 24532 2836
rect 24504 2666 24532 2808
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23572 2644 23624 2650
rect 24504 2638 24624 2666
rect 23572 2586 23624 2592
rect 22650 2544 22706 2553
rect 22650 2479 22652 2488
rect 22704 2479 22706 2488
rect 22652 2450 22704 2456
rect 23400 2446 23428 2586
rect 23584 2514 23612 2586
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 22100 604 22152 610
rect 22100 546 22152 552
rect 22284 604 22336 610
rect 22284 546 22336 552
rect 22296 480 22324 546
rect 24596 480 24624 2638
rect 24688 2446 24716 3839
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 24780 2582 24808 2926
rect 24872 2650 24900 3470
rect 25056 2922 25084 3946
rect 25148 3738 25176 4558
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25516 3398 25544 4014
rect 26160 3670 26188 4558
rect 26252 4078 26280 4694
rect 26790 4448 26846 4457
rect 26790 4383 26846 4392
rect 26240 4072 26292 4078
rect 26240 4014 26292 4020
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26252 3738 26280 4014
rect 26344 3942 26372 4014
rect 26332 3936 26384 3942
rect 26330 3904 26332 3913
rect 26384 3904 26386 3913
rect 26330 3839 26386 3848
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26148 3664 26200 3670
rect 26148 3606 26200 3612
rect 26804 3534 26832 4383
rect 26896 3670 26924 4927
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 25504 3392 25556 3398
rect 25502 3360 25504 3369
rect 25556 3360 25558 3369
rect 25502 3295 25558 3304
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 26344 2650 26372 3470
rect 26896 3194 26924 3606
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 26698 2544 26754 2553
rect 26698 2479 26700 2488
rect 26752 2479 26754 2488
rect 26700 2450 26752 2456
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 25964 2304 26016 2310
rect 25962 2272 25964 2281
rect 26016 2272 26018 2281
rect 25962 2207 26018 2216
rect 27080 2145 27108 6122
rect 27264 5710 27292 6258
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 27342 5672 27398 5681
rect 27264 5234 27292 5646
rect 27342 5607 27398 5616
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 27264 4622 27292 5170
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 27160 4548 27212 4554
rect 27160 4490 27212 4496
rect 27172 3126 27200 4490
rect 27356 4434 27384 5607
rect 27264 4406 27384 4434
rect 27160 3120 27212 3126
rect 27160 3062 27212 3068
rect 27264 2650 27292 4406
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27356 3670 27384 3878
rect 27344 3664 27396 3670
rect 27344 3606 27396 3612
rect 27252 2644 27304 2650
rect 27252 2586 27304 2592
rect 27066 2136 27122 2145
rect 27066 2071 27122 2080
rect 26974 2000 27030 2009
rect 26974 1935 27030 1944
rect 26988 480 27016 1935
rect 27448 1465 27476 6326
rect 27816 6186 27844 6734
rect 28092 6458 28120 6802
rect 28080 6452 28132 6458
rect 28080 6394 28132 6400
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28184 5710 28212 7375
rect 28276 7342 28304 9143
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 28264 5840 28316 5846
rect 28264 5782 28316 5788
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28184 5234 28212 5510
rect 28276 5370 28304 5782
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 28368 5370 28396 5646
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28356 5364 28408 5370
rect 28356 5306 28408 5312
rect 28460 5273 28488 9862
rect 28632 9648 28684 9654
rect 28632 9590 28684 9596
rect 28540 8968 28592 8974
rect 28644 8945 28672 9590
rect 28920 9382 28948 10066
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28908 9376 28960 9382
rect 28908 9318 28960 9324
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 28540 8910 28592 8916
rect 28630 8936 28686 8945
rect 28552 8362 28580 8910
rect 28630 8871 28686 8880
rect 28540 8356 28592 8362
rect 28540 8298 28592 8304
rect 28552 7886 28580 8298
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28552 7002 28580 7822
rect 28644 7546 28672 7958
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28644 7002 28672 7482
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 28632 6996 28684 7002
rect 28632 6938 28684 6944
rect 28446 5264 28502 5273
rect 28172 5228 28224 5234
rect 28446 5199 28502 5208
rect 28172 5170 28224 5176
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28184 4622 28212 5170
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28078 4040 28134 4049
rect 28078 3975 28134 3984
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28092 3738 28120 3975
rect 28184 3942 28212 4558
rect 28276 4282 28304 4694
rect 28736 4486 28764 9318
rect 28908 9172 28960 9178
rect 28908 9114 28960 9120
rect 28920 9081 28948 9114
rect 29000 9104 29052 9110
rect 28906 9072 28962 9081
rect 29104 9081 29132 9318
rect 29000 9046 29052 9052
rect 29090 9072 29146 9081
rect 28906 9007 28962 9016
rect 29012 8634 29040 9046
rect 29090 9007 29146 9016
rect 29196 8974 29224 9998
rect 29184 8968 29236 8974
rect 29184 8910 29236 8916
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29196 8566 29224 8910
rect 29184 8560 29236 8566
rect 29184 8502 29236 8508
rect 29196 7410 29224 8502
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29196 7002 29224 7346
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 28998 6352 29054 6361
rect 28998 6287 29000 6296
rect 29052 6287 29054 6296
rect 29000 6258 29052 6264
rect 29276 5704 29328 5710
rect 29274 5672 29276 5681
rect 29328 5672 29330 5681
rect 29274 5607 29330 5616
rect 29380 5098 29408 11047
rect 34060 11008 34112 11014
rect 34164 10985 34192 11154
rect 34060 10950 34112 10956
rect 34150 10976 34206 10985
rect 33414 10840 33470 10849
rect 33414 10775 33470 10784
rect 32310 10704 32366 10713
rect 32310 10639 32366 10648
rect 32324 9654 32352 10639
rect 33428 10606 33456 10775
rect 33416 10600 33468 10606
rect 33416 10542 33468 10548
rect 33428 10130 33456 10542
rect 33600 10464 33652 10470
rect 33600 10406 33652 10412
rect 33784 10464 33836 10470
rect 33784 10406 33836 10412
rect 33416 10124 33468 10130
rect 33416 10066 33468 10072
rect 33428 9722 33456 10066
rect 33416 9716 33468 9722
rect 33416 9658 33468 9664
rect 32312 9648 32364 9654
rect 32312 9590 32364 9596
rect 32586 9616 32642 9625
rect 32586 9551 32588 9560
rect 32640 9551 32642 9560
rect 32588 9522 32640 9528
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 29828 9376 29880 9382
rect 29826 9344 29828 9353
rect 29880 9344 29882 9353
rect 29826 9279 29882 9288
rect 29840 8906 29868 9279
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29472 7750 29500 8434
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29460 7744 29512 7750
rect 29458 7712 29460 7721
rect 29512 7712 29514 7721
rect 29458 7647 29514 7656
rect 29656 7410 29684 7822
rect 29826 7576 29882 7585
rect 29826 7511 29882 7520
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29460 7268 29512 7274
rect 29460 7210 29512 7216
rect 29472 7002 29500 7210
rect 29460 6996 29512 7002
rect 29460 6938 29512 6944
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 29564 6225 29592 6734
rect 29550 6216 29606 6225
rect 29550 6151 29606 6160
rect 29564 5914 29592 6151
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29368 5092 29420 5098
rect 29368 5034 29420 5040
rect 29380 4826 29408 5034
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 28816 4616 28868 4622
rect 28816 4558 28868 4564
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 28724 4480 28776 4486
rect 28724 4422 28776 4428
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28172 3936 28224 3942
rect 28368 3913 28396 4422
rect 28828 4321 28856 4558
rect 28814 4312 28870 4321
rect 28814 4247 28870 4256
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 28724 4004 28776 4010
rect 28724 3946 28776 3952
rect 28172 3878 28224 3884
rect 28354 3904 28410 3913
rect 28354 3839 28410 3848
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 28092 2990 28120 3674
rect 28736 3670 28764 3946
rect 28724 3664 28776 3670
rect 28724 3606 28776 3612
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 28184 3194 28212 3470
rect 28736 3194 28764 3606
rect 29564 3398 29592 4014
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 29368 3392 29420 3398
rect 29552 3392 29604 3398
rect 29420 3352 29500 3380
rect 29368 3334 29420 3340
rect 28172 3188 28224 3194
rect 28172 3130 28224 3136
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 28184 2582 28212 3130
rect 28920 2650 28948 3334
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 28172 2576 28224 2582
rect 27710 2544 27766 2553
rect 28172 2518 28224 2524
rect 27710 2479 27712 2488
rect 27764 2479 27766 2488
rect 27712 2450 27764 2456
rect 27434 1456 27490 1465
rect 27434 1391 27490 1400
rect 29380 480 29408 2994
rect 29472 2922 29500 3352
rect 29552 3334 29604 3340
rect 29460 2916 29512 2922
rect 29460 2858 29512 2864
rect 29458 2816 29514 2825
rect 29458 2751 29514 2760
rect 29472 2650 29500 2751
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29564 2553 29592 3334
rect 29656 3058 29684 7346
rect 29840 7274 29868 7511
rect 29828 7268 29880 7274
rect 29828 7210 29880 7216
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 29748 5710 29776 6190
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29734 4176 29790 4185
rect 29734 4111 29790 4120
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29748 2854 29776 4111
rect 29736 2848 29788 2854
rect 29840 2825 29868 7210
rect 29920 4072 29972 4078
rect 29920 4014 29972 4020
rect 29736 2790 29788 2796
rect 29826 2816 29882 2825
rect 29826 2751 29882 2760
rect 29932 2650 29960 4014
rect 30104 4004 30156 4010
rect 30104 3946 30156 3952
rect 30116 3738 30144 3946
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30208 3641 30236 9454
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 32680 9376 32732 9382
rect 32680 9318 32732 9324
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33508 9376 33560 9382
rect 33508 9318 33560 9324
rect 30380 9036 30432 9042
rect 30380 8978 30432 8984
rect 30392 8362 30420 8978
rect 30380 8356 30432 8362
rect 30380 8298 30432 8304
rect 30392 7993 30420 8298
rect 30378 7984 30434 7993
rect 30378 7919 30434 7928
rect 30484 6866 30512 9318
rect 32312 9036 32364 9042
rect 32312 8978 32364 8984
rect 30564 8832 30616 8838
rect 30564 8774 30616 8780
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30392 6100 30420 6802
rect 30472 6112 30524 6118
rect 30392 6072 30472 6100
rect 30472 6054 30524 6060
rect 30484 5846 30512 6054
rect 30472 5840 30524 5846
rect 30472 5782 30524 5788
rect 30288 5704 30340 5710
rect 30288 5646 30340 5652
rect 30300 4978 30328 5646
rect 30484 5166 30512 5782
rect 30472 5160 30524 5166
rect 30472 5102 30524 5108
rect 30380 5024 30432 5030
rect 30300 4972 30380 4978
rect 30300 4966 30432 4972
rect 30300 4950 30420 4966
rect 30194 3632 30250 3641
rect 30194 3567 30250 3576
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 29920 2644 29972 2650
rect 29920 2586 29972 2592
rect 30116 2582 30144 2994
rect 30104 2576 30156 2582
rect 29550 2544 29606 2553
rect 30104 2518 30156 2524
rect 29550 2479 29606 2488
rect 30300 2446 30328 4950
rect 30378 4720 30434 4729
rect 30378 4655 30380 4664
rect 30432 4655 30434 4664
rect 30380 4626 30432 4632
rect 30392 4282 30420 4626
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30484 3670 30512 5102
rect 30576 4457 30604 8774
rect 31404 8430 31432 8774
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 30748 7948 30800 7954
rect 30748 7890 30800 7896
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 30760 7857 30788 7890
rect 30746 7848 30802 7857
rect 30746 7783 30802 7792
rect 30760 7206 30788 7783
rect 31312 7342 31340 7890
rect 31404 7410 31432 8366
rect 32324 8362 32352 8978
rect 32692 8401 32720 9318
rect 32772 9036 32824 9042
rect 32772 8978 32824 8984
rect 32678 8392 32734 8401
rect 32312 8356 32364 8362
rect 32784 8362 32812 8978
rect 33336 8974 33364 9318
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 32678 8327 32734 8336
rect 32772 8356 32824 8362
rect 32312 8298 32364 8304
rect 32772 8298 32824 8304
rect 32220 8288 32272 8294
rect 32220 8230 32272 8236
rect 32232 8022 32260 8230
rect 32220 8016 32272 8022
rect 32220 7958 32272 7964
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32140 7546 32168 7822
rect 32128 7540 32180 7546
rect 32128 7482 32180 7488
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 30748 7200 30800 7206
rect 30748 7142 30800 7148
rect 30562 4448 30618 4457
rect 30562 4383 30618 4392
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30484 3194 30512 3606
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30760 2990 30788 7142
rect 31312 6662 31340 7278
rect 32232 7206 32260 7958
rect 32220 7200 32272 7206
rect 32220 7142 32272 7148
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 30932 6656 30984 6662
rect 30932 6598 30984 6604
rect 31300 6656 31352 6662
rect 31300 6598 31352 6604
rect 30838 6488 30894 6497
rect 30838 6423 30840 6432
rect 30892 6423 30894 6432
rect 30840 6394 30892 6400
rect 30944 6118 30972 6598
rect 31588 6254 31616 6802
rect 32140 6458 32168 6802
rect 32232 6458 32260 7142
rect 32128 6452 32180 6458
rect 32128 6394 32180 6400
rect 32220 6452 32272 6458
rect 32220 6394 32272 6400
rect 31576 6248 31628 6254
rect 31576 6190 31628 6196
rect 30932 6112 30984 6118
rect 30932 6054 30984 6060
rect 31206 6080 31262 6089
rect 30840 5160 30892 5166
rect 30840 5102 30892 5108
rect 30852 3505 30880 5102
rect 30944 5030 30972 6054
rect 31206 6015 31262 6024
rect 31220 5914 31248 6015
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31206 5808 31262 5817
rect 31206 5743 31262 5752
rect 30932 5024 30984 5030
rect 30932 4966 30984 4972
rect 30944 4690 30972 4966
rect 31220 4758 31248 5743
rect 31208 4752 31260 4758
rect 31208 4694 31260 4700
rect 30932 4684 30984 4690
rect 30932 4626 30984 4632
rect 30944 4146 30972 4626
rect 31484 4480 31536 4486
rect 31484 4422 31536 4428
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 31496 4010 31524 4422
rect 31588 4162 31616 6190
rect 31852 6180 31904 6186
rect 31852 6122 31904 6128
rect 31864 5234 31892 6122
rect 32232 5846 32260 6394
rect 32324 6361 32352 8298
rect 32784 6866 32812 8298
rect 32772 6860 32824 6866
rect 32772 6802 32824 6808
rect 32310 6352 32366 6361
rect 32310 6287 32366 6296
rect 32220 5840 32272 5846
rect 32220 5782 32272 5788
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 31852 5228 31904 5234
rect 31852 5170 31904 5176
rect 31588 4134 31708 4162
rect 31574 4040 31630 4049
rect 31116 4004 31168 4010
rect 31116 3946 31168 3952
rect 31484 4004 31536 4010
rect 31574 3975 31576 3984
rect 31484 3946 31536 3952
rect 31628 3975 31630 3984
rect 31576 3946 31628 3952
rect 31128 3602 31156 3946
rect 31496 3738 31524 3946
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31116 3596 31168 3602
rect 31116 3538 31168 3544
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31484 3528 31536 3534
rect 30838 3496 30894 3505
rect 31484 3470 31536 3476
rect 30838 3431 30894 3440
rect 31496 2990 31524 3470
rect 31588 3346 31616 3538
rect 31680 3534 31708 4134
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 31588 3318 31800 3346
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31312 2650 31340 2926
rect 31772 2650 31800 3318
rect 31956 3058 31984 5646
rect 32232 5302 32260 5782
rect 32220 5296 32272 5302
rect 32220 5238 32272 5244
rect 32232 5098 32260 5238
rect 32220 5092 32272 5098
rect 32220 5034 32272 5040
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32140 4185 32168 4558
rect 32220 4276 32272 4282
rect 32220 4218 32272 4224
rect 32126 4176 32182 4185
rect 32126 4111 32182 4120
rect 32232 3602 32260 4218
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 32232 3194 32260 3538
rect 32220 3188 32272 3194
rect 32220 3130 32272 3136
rect 31944 3052 31996 3058
rect 31944 2994 31996 3000
rect 32324 2990 32352 6287
rect 32968 5794 32996 8910
rect 33324 8832 33376 8838
rect 33324 8774 33376 8780
rect 33336 8362 33364 8774
rect 33324 8356 33376 8362
rect 33324 8298 33376 8304
rect 33520 8090 33548 9318
rect 33612 9178 33640 10406
rect 33692 9512 33744 9518
rect 33692 9454 33744 9460
rect 33704 9217 33732 9454
rect 33690 9208 33746 9217
rect 33600 9172 33652 9178
rect 33690 9143 33746 9152
rect 33600 9114 33652 9120
rect 33612 8498 33640 9114
rect 33796 8809 33824 10406
rect 33874 10296 33930 10305
rect 33874 10231 33930 10240
rect 33888 9897 33916 10231
rect 33874 9888 33930 9897
rect 33874 9823 33930 9832
rect 34072 9217 34100 10950
rect 34150 10911 34206 10920
rect 34164 10470 34192 10911
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 35268 10606 35296 11154
rect 35452 10713 35480 12718
rect 35438 10704 35494 10713
rect 35438 10639 35494 10648
rect 35256 10600 35308 10606
rect 35256 10542 35308 10548
rect 35440 10600 35492 10606
rect 35440 10542 35492 10548
rect 34152 10464 34204 10470
rect 34152 10406 34204 10412
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34702 10160 34758 10169
rect 34702 10095 34704 10104
rect 34756 10095 34758 10104
rect 34704 10066 34756 10072
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 34058 9208 34114 9217
rect 34058 9143 34114 9152
rect 34060 9104 34112 9110
rect 34060 9046 34112 9052
rect 34164 9058 34192 9862
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34716 9382 34744 10066
rect 34808 9897 34836 10406
rect 35452 10305 35480 10542
rect 35438 10296 35494 10305
rect 35438 10231 35494 10240
rect 35256 9920 35308 9926
rect 34794 9888 34850 9897
rect 35256 9862 35308 9868
rect 35348 9920 35400 9926
rect 35348 9862 35400 9868
rect 35438 9888 35494 9897
rect 34794 9823 34850 9832
rect 35162 9616 35218 9625
rect 35162 9551 35164 9560
rect 35216 9551 35218 9560
rect 35164 9522 35216 9528
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 35164 9376 35216 9382
rect 35164 9318 35216 9324
rect 34886 9072 34942 9081
rect 33876 8900 33928 8906
rect 33876 8842 33928 8848
rect 33782 8800 33838 8809
rect 33782 8735 33838 8744
rect 33888 8566 33916 8842
rect 33966 8664 34022 8673
rect 34072 8634 34100 9046
rect 34164 9030 34376 9058
rect 34348 8974 34376 9030
rect 34886 9007 34942 9016
rect 34152 8968 34204 8974
rect 34152 8910 34204 8916
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 33966 8599 34022 8608
rect 34060 8628 34112 8634
rect 33876 8560 33928 8566
rect 33876 8502 33928 8508
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33980 8294 34008 8599
rect 34060 8570 34112 8576
rect 33968 8288 34020 8294
rect 33968 8230 34020 8236
rect 33508 8084 33560 8090
rect 33508 8026 33560 8032
rect 33048 7948 33100 7954
rect 33048 7890 33100 7896
rect 33060 7546 33088 7890
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 33060 7274 33088 7482
rect 33520 7410 33548 8026
rect 33874 7984 33930 7993
rect 33874 7919 33876 7928
rect 33928 7919 33930 7928
rect 33876 7890 33928 7896
rect 33888 7546 33916 7890
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33336 6186 33364 6598
rect 33324 6180 33376 6186
rect 33324 6122 33376 6128
rect 33140 6112 33192 6118
rect 33138 6080 33140 6089
rect 33192 6080 33194 6089
rect 33138 6015 33194 6024
rect 33046 5944 33102 5953
rect 33046 5879 33048 5888
rect 33100 5879 33102 5888
rect 33048 5850 33100 5856
rect 32968 5778 33180 5794
rect 32968 5772 33192 5778
rect 32968 5766 33140 5772
rect 33140 5714 33192 5720
rect 33048 5704 33100 5710
rect 33048 5646 33100 5652
rect 33060 5386 33088 5646
rect 33060 5370 33180 5386
rect 33060 5364 33192 5370
rect 33060 5358 33140 5364
rect 33140 5306 33192 5312
rect 33336 5273 33364 6122
rect 33704 5914 33732 6802
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 33322 5264 33378 5273
rect 32956 5228 33008 5234
rect 33980 5250 34008 8230
rect 34072 8022 34100 8570
rect 34164 8090 34192 8910
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34152 8084 34204 8090
rect 34152 8026 34204 8032
rect 34060 8016 34112 8022
rect 34060 7958 34112 7964
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 34164 7449 34192 7686
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34150 7440 34206 7449
rect 34150 7375 34206 7384
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 34164 6458 34192 6870
rect 34624 6730 34652 8298
rect 34704 8016 34756 8022
rect 34704 7958 34756 7964
rect 34716 7206 34744 7958
rect 34796 7812 34848 7818
rect 34796 7754 34848 7760
rect 34808 7410 34836 7754
rect 34900 7585 34928 9007
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34992 8498 35020 8774
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 35070 8392 35126 8401
rect 35070 8327 35126 8336
rect 34886 7576 34942 7585
rect 34886 7511 34942 7520
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 34704 7200 34756 7206
rect 34704 7142 34756 7148
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34716 6934 34744 7142
rect 34704 6928 34756 6934
rect 34704 6870 34756 6876
rect 34612 6724 34664 6730
rect 34612 6666 34664 6672
rect 34808 6662 34836 7142
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34152 6452 34204 6458
rect 34152 6394 34204 6400
rect 34164 5846 34192 6394
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34440 6100 34468 6190
rect 34440 6072 34652 6100
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 34060 5772 34112 5778
rect 34060 5714 34112 5720
rect 34072 5370 34100 5714
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34624 5370 34652 6072
rect 34808 5914 34836 6598
rect 35084 5914 35112 8327
rect 35176 6100 35204 9318
rect 35268 6225 35296 9862
rect 35360 6866 35388 9862
rect 35438 9823 35494 9832
rect 35452 7324 35480 9823
rect 35544 9654 35572 15535
rect 35714 14648 35770 14657
rect 35714 14583 35770 14592
rect 35622 13832 35678 13841
rect 35622 13767 35678 13776
rect 35636 12986 35664 13767
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35622 12064 35678 12073
rect 35622 11999 35678 12008
rect 35636 11354 35664 11999
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35622 11112 35678 11121
rect 35622 11047 35678 11056
rect 35636 10810 35664 11047
rect 35624 10804 35676 10810
rect 35624 10746 35676 10752
rect 35728 10266 35756 14583
rect 36818 12880 36874 12889
rect 36818 12815 36874 12824
rect 36266 10568 36322 10577
rect 36266 10503 36322 10512
rect 35716 10260 35768 10266
rect 35716 10202 35768 10208
rect 36280 10130 36308 10503
rect 36634 10296 36690 10305
rect 36634 10231 36690 10240
rect 35808 10124 35860 10130
rect 35808 10066 35860 10072
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 35532 9648 35584 9654
rect 35532 9590 35584 9596
rect 35820 9602 35848 10066
rect 36648 9654 36676 10231
rect 36636 9648 36688 9654
rect 35820 9574 35940 9602
rect 36636 9590 36688 9596
rect 35912 9382 35940 9574
rect 36452 9512 36504 9518
rect 36450 9480 36452 9489
rect 36504 9480 36506 9489
rect 36084 9444 36136 9450
rect 36450 9415 36506 9424
rect 36084 9386 36136 9392
rect 35900 9376 35952 9382
rect 35898 9344 35900 9353
rect 35952 9344 35954 9353
rect 35898 9279 35954 9288
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35636 8634 35664 9046
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35532 8560 35584 8566
rect 35532 8502 35584 8508
rect 35544 8090 35572 8502
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35544 7478 35572 8026
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35532 7472 35584 7478
rect 35532 7414 35584 7420
rect 35636 7410 35664 7822
rect 35624 7404 35676 7410
rect 35676 7364 35756 7392
rect 35624 7346 35676 7352
rect 35452 7296 35572 7324
rect 35348 6860 35400 6866
rect 35348 6802 35400 6808
rect 35360 6322 35388 6802
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 35254 6216 35310 6225
rect 35254 6151 35310 6160
rect 35176 6072 35388 6100
rect 34796 5908 34848 5914
rect 34796 5850 34848 5856
rect 35072 5908 35124 5914
rect 35072 5850 35124 5856
rect 35084 5710 35112 5850
rect 35072 5704 35124 5710
rect 35072 5646 35124 5652
rect 34060 5364 34112 5370
rect 34060 5306 34112 5312
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 34980 5364 35032 5370
rect 34980 5306 35032 5312
rect 34704 5296 34756 5302
rect 33980 5222 34100 5250
rect 34704 5238 34756 5244
rect 33322 5199 33378 5208
rect 32956 5170 33008 5176
rect 32968 4826 32996 5170
rect 33692 5092 33744 5098
rect 33692 5034 33744 5040
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 33704 4758 33732 5034
rect 33692 4752 33744 4758
rect 33692 4694 33744 4700
rect 32586 4584 32642 4593
rect 32586 4519 32588 4528
rect 32640 4519 32642 4528
rect 32588 4490 32640 4496
rect 32600 4078 32628 4490
rect 33704 4282 33732 4694
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 33692 4276 33744 4282
rect 33692 4218 33744 4224
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 33324 4004 33376 4010
rect 33324 3946 33376 3952
rect 33336 3602 33364 3946
rect 33704 3652 33732 4218
rect 33980 3942 34008 4558
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 33784 3664 33836 3670
rect 33704 3624 33784 3652
rect 33324 3596 33376 3602
rect 33324 3538 33376 3544
rect 33336 3194 33364 3538
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 33704 3126 33732 3624
rect 33784 3606 33836 3612
rect 33692 3120 33744 3126
rect 33692 3062 33744 3068
rect 33980 3058 34008 3878
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 32864 2984 32916 2990
rect 32864 2926 32916 2932
rect 32876 2650 32904 2926
rect 34072 2650 34100 5222
rect 34612 4480 34664 4486
rect 34612 4422 34664 4428
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 34624 4146 34652 4422
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34624 3942 34652 4082
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 34716 3194 34744 5238
rect 34992 5234 35020 5306
rect 34980 5228 35032 5234
rect 34980 5170 35032 5176
rect 35256 5228 35308 5234
rect 35256 5170 35308 5176
rect 34992 4826 35020 5170
rect 35072 5092 35124 5098
rect 35072 5034 35124 5040
rect 35084 4826 35112 5034
rect 34980 4820 35032 4826
rect 34980 4762 35032 4768
rect 35072 4820 35124 4826
rect 35072 4762 35124 4768
rect 34992 3380 35020 4762
rect 35164 4616 35216 4622
rect 35164 4558 35216 4564
rect 35176 3534 35204 4558
rect 35268 4146 35296 5170
rect 35256 4140 35308 4146
rect 35256 4082 35308 4088
rect 35268 4049 35296 4082
rect 35254 4040 35310 4049
rect 35254 3975 35310 3984
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 34992 3352 35112 3380
rect 34978 3224 35034 3233
rect 34704 3188 34756 3194
rect 34978 3159 35034 3168
rect 34704 3130 34756 3136
rect 34716 2922 34744 3130
rect 34992 3058 35020 3159
rect 35084 3058 35112 3352
rect 34980 3052 35032 3058
rect 34980 2994 35032 3000
rect 35072 3052 35124 3058
rect 35072 2994 35124 3000
rect 34704 2916 34756 2922
rect 34704 2858 34756 2864
rect 34992 2650 35020 2994
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 34060 2644 34112 2650
rect 34060 2586 34112 2592
rect 34980 2644 35032 2650
rect 34980 2586 35032 2592
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 34058 2272 34114 2281
rect 31680 480 31708 2246
rect 33152 2145 33180 2246
rect 34058 2207 34114 2216
rect 33138 2136 33194 2145
rect 33138 2071 33194 2080
rect 34072 480 34100 2207
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 35360 1329 35388 6072
rect 35452 5846 35480 6734
rect 35440 5840 35492 5846
rect 35438 5808 35440 5817
rect 35492 5808 35494 5817
rect 35438 5743 35494 5752
rect 35544 4865 35572 7296
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35636 5370 35664 6258
rect 35624 5364 35676 5370
rect 35624 5306 35676 5312
rect 35530 4856 35586 4865
rect 35530 4791 35586 4800
rect 35728 3618 35756 7364
rect 35900 7200 35952 7206
rect 35820 7148 35900 7154
rect 35820 7142 35952 7148
rect 35820 7126 35940 7142
rect 35820 6730 35848 7126
rect 35900 6928 35952 6934
rect 35900 6870 35952 6876
rect 35808 6724 35860 6730
rect 35808 6666 35860 6672
rect 35912 6458 35940 6870
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 35808 6248 35860 6254
rect 35808 6190 35860 6196
rect 35820 5953 35848 6190
rect 35992 6180 36044 6186
rect 35992 6122 36044 6128
rect 35806 5944 35862 5953
rect 35806 5879 35862 5888
rect 35820 5846 35848 5879
rect 35808 5840 35860 5846
rect 35860 5788 35940 5794
rect 35808 5782 35940 5788
rect 35820 5766 35940 5782
rect 35912 5370 35940 5766
rect 36004 5710 36032 6122
rect 35992 5704 36044 5710
rect 35992 5646 36044 5652
rect 35900 5364 35952 5370
rect 35900 5306 35952 5312
rect 36004 5234 36032 5646
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 35900 4752 35952 4758
rect 35900 4694 35952 4700
rect 35912 4282 35940 4694
rect 36004 4282 36032 5170
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 35728 3590 36032 3618
rect 36004 3534 36032 3590
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 35912 3194 35940 3470
rect 35900 3188 35952 3194
rect 35900 3130 35952 3136
rect 36004 2650 36032 3470
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 35900 2440 35952 2446
rect 35898 2408 35900 2417
rect 35952 2408 35954 2417
rect 35898 2343 35954 2352
rect 35346 1320 35402 1329
rect 35346 1255 35402 1264
rect 36096 513 36124 9386
rect 36634 9344 36690 9353
rect 36634 9279 36690 9288
rect 36358 9208 36414 9217
rect 36358 9143 36414 9152
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36280 8634 36308 8910
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36268 8424 36320 8430
rect 36268 8366 36320 8372
rect 36280 7313 36308 8366
rect 36266 7304 36322 7313
rect 36266 7239 36322 7248
rect 36372 5098 36400 9143
rect 36648 8634 36676 9279
rect 36728 8900 36780 8906
rect 36728 8842 36780 8848
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 36634 8528 36690 8537
rect 36634 8463 36690 8472
rect 36648 8090 36676 8463
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36452 7948 36504 7954
rect 36452 7890 36504 7896
rect 36464 7546 36492 7890
rect 36740 7818 36768 8842
rect 36728 7812 36780 7818
rect 36728 7754 36780 7760
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36542 7440 36598 7449
rect 36740 7410 36768 7754
rect 36542 7375 36544 7384
rect 36596 7375 36598 7384
rect 36728 7404 36780 7410
rect 36544 7346 36596 7352
rect 36728 7346 36780 7352
rect 36556 7002 36584 7346
rect 36544 6996 36596 7002
rect 36544 6938 36596 6944
rect 36542 6216 36598 6225
rect 36542 6151 36544 6160
rect 36596 6151 36598 6160
rect 36544 6122 36596 6128
rect 36556 5914 36584 6122
rect 36544 5908 36596 5914
rect 36544 5850 36596 5856
rect 36636 5296 36688 5302
rect 36636 5238 36688 5244
rect 36648 5098 36676 5238
rect 36360 5092 36412 5098
rect 36360 5034 36412 5040
rect 36636 5092 36688 5098
rect 36636 5034 36688 5040
rect 36372 4826 36400 5034
rect 36360 4820 36412 4826
rect 36360 4762 36412 4768
rect 36358 4176 36414 4185
rect 36358 4111 36414 4120
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 36280 3194 36308 3606
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 36372 2514 36400 4111
rect 36452 4072 36504 4078
rect 36452 4014 36504 4020
rect 36464 3913 36492 4014
rect 36832 3942 36860 12815
rect 37188 10124 37240 10130
rect 37188 10066 37240 10072
rect 37200 9330 37228 10066
rect 37280 9376 37332 9382
rect 37200 9324 37280 9330
rect 37200 9318 37332 9324
rect 37200 9302 37320 9318
rect 37200 5817 37228 9302
rect 38016 8424 38068 8430
rect 38016 8366 38068 8372
rect 37554 7304 37610 7313
rect 37554 7239 37610 7248
rect 37186 5808 37242 5817
rect 37186 5743 37242 5752
rect 37370 5264 37426 5273
rect 37370 5199 37426 5208
rect 37004 4072 37056 4078
rect 37004 4014 37056 4020
rect 36820 3936 36872 3942
rect 36450 3904 36506 3913
rect 36820 3878 36872 3884
rect 36450 3839 36506 3848
rect 37016 2990 37044 4014
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 37292 3233 37320 3878
rect 37278 3224 37334 3233
rect 37384 3194 37412 5199
rect 37568 4078 37596 7239
rect 37556 4072 37608 4078
rect 38028 4049 38056 8366
rect 37556 4014 37608 4020
rect 38014 4040 38070 4049
rect 38014 3975 38070 3984
rect 37278 3159 37334 3168
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 39394 3088 39450 3097
rect 39394 3023 39450 3032
rect 37004 2984 37056 2990
rect 39408 2961 39436 3023
rect 37004 2926 37056 2932
rect 39394 2952 39450 2961
rect 39394 2887 39450 2896
rect 38750 2680 38806 2689
rect 38750 2615 38806 2624
rect 36360 2508 36412 2514
rect 36360 2450 36412 2456
rect 36360 2372 36412 2378
rect 36360 2314 36412 2320
rect 36082 504 36138 513
rect 2778 439 2834 448
rect 3422 0 3478 480
rect 5814 0 5870 480
rect 8114 0 8170 480
rect 10506 0 10562 480
rect 12806 0 12862 480
rect 15198 0 15254 480
rect 17590 0 17646 480
rect 19890 0 19946 480
rect 22282 0 22338 480
rect 24582 0 24638 480
rect 26974 0 27030 480
rect 29366 0 29422 480
rect 31666 0 31722 480
rect 34058 0 34114 480
rect 36372 480 36400 2314
rect 38764 480 38792 2615
rect 36082 439 36138 448
rect 36358 0 36414 480
rect 38750 0 38806 480
<< via2 >>
rect 1398 15544 1454 15600
rect 35530 15544 35586 15600
rect 1490 14592 1546 14648
rect 1582 13776 1638 13832
rect 2962 12824 3018 12880
rect 1674 11500 1676 11520
rect 1676 11500 1728 11520
rect 1728 11500 1730 11520
rect 1674 11464 1730 11500
rect 570 8472 626 8528
rect 570 4800 626 4856
rect 1122 3712 1178 3768
rect 2042 10412 2044 10432
rect 2044 10412 2096 10432
rect 2096 10412 2098 10432
rect 2042 10376 2098 10412
rect 2134 8880 2190 8936
rect 2318 8780 2320 8800
rect 2320 8780 2372 8800
rect 2372 8780 2374 8800
rect 2318 8744 2374 8780
rect 2502 8608 2558 8664
rect 2686 11056 2742 11112
rect 1582 5364 1638 5400
rect 1582 5344 1584 5364
rect 1584 5344 1636 5364
rect 1636 5344 1638 5364
rect 2778 5480 2834 5536
rect 3330 11328 3386 11384
rect 3422 10920 3478 10976
rect 3054 10124 3110 10160
rect 3054 10104 3056 10124
rect 3056 10104 3108 10124
rect 3108 10104 3110 10124
rect 3054 8492 3110 8528
rect 3054 8472 3056 8492
rect 3056 8472 3108 8492
rect 3108 8472 3110 8492
rect 3146 5888 3202 5944
rect 3330 9832 3386 9888
rect 2962 5344 3018 5400
rect 1674 2896 1730 2952
rect 2502 4004 2558 4040
rect 2502 3984 2504 4004
rect 2504 3984 2556 4004
rect 2556 3984 2558 4004
rect 3054 4428 3056 4448
rect 3056 4428 3108 4448
rect 3108 4428 3110 4448
rect 3054 4392 3110 4428
rect 3330 5480 3386 5536
rect 3606 10240 3662 10296
rect 4066 12008 4122 12064
rect 3974 11736 4030 11792
rect 3698 9444 3754 9480
rect 3698 9424 3700 9444
rect 3700 9424 3752 9444
rect 3752 9424 3754 9444
rect 3882 9172 3938 9208
rect 3882 9152 3884 9172
rect 3884 9152 3936 9172
rect 3936 9152 3938 9172
rect 3790 8336 3846 8392
rect 3606 8064 3662 8120
rect 3790 6840 3846 6896
rect 3514 3984 3570 4040
rect 4894 11192 4950 11248
rect 4802 11056 4858 11112
rect 4250 10668 4306 10704
rect 4250 10648 4252 10668
rect 4252 10648 4304 10668
rect 4304 10648 4306 10668
rect 4342 9288 4398 9344
rect 4250 9152 4306 9208
rect 4066 7520 4122 7576
rect 4434 8916 4436 8936
rect 4436 8916 4488 8936
rect 4488 8916 4490 8936
rect 4434 8880 4490 8916
rect 4526 7928 4582 7984
rect 4710 8336 4766 8392
rect 3974 5344 4030 5400
rect 4158 4800 4214 4856
rect 4802 4564 4804 4584
rect 4804 4564 4856 4584
rect 4856 4564 4858 4584
rect 4802 4528 4858 4564
rect 3790 3848 3846 3904
rect 3422 3032 3478 3088
rect 4710 4140 4766 4176
rect 4710 4120 4712 4140
rect 4712 4120 4764 4140
rect 4764 4120 4766 4140
rect 4250 4004 4306 4040
rect 4250 3984 4252 4004
rect 4252 3984 4304 4004
rect 4304 3984 4306 4004
rect 5170 9968 5226 10024
rect 5446 11736 5502 11792
rect 6182 11600 6238 11656
rect 5538 10512 5594 10568
rect 5722 10376 5778 10432
rect 5722 8880 5778 8936
rect 5538 8472 5594 8528
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5538 5364 5594 5400
rect 5538 5344 5540 5364
rect 5540 5344 5592 5364
rect 5592 5344 5594 5364
rect 5906 9288 5962 9344
rect 5906 6568 5962 6624
rect 5722 4392 5778 4448
rect 5538 3848 5594 3904
rect 5354 3576 5410 3632
rect 2778 448 2834 504
rect 4894 2216 4950 2272
rect 6274 7828 6276 7848
rect 6276 7828 6328 7848
rect 6328 7828 6330 7848
rect 6274 7792 6330 7828
rect 6182 6976 6238 7032
rect 6182 6840 6238 6896
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 6458 10512 6514 10568
rect 6550 9016 6606 9072
rect 6550 8744 6606 8800
rect 6274 5888 6330 5944
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 6918 11056 6974 11112
rect 7102 11464 7158 11520
rect 7010 10920 7066 10976
rect 7194 10240 7250 10296
rect 7194 9832 7250 9888
rect 7102 9424 7158 9480
rect 7010 9152 7066 9208
rect 7010 8336 7066 8392
rect 6918 7656 6974 7712
rect 6826 7404 6882 7440
rect 6826 7384 6828 7404
rect 6828 7384 6880 7404
rect 6880 7384 6882 7404
rect 7010 6704 7066 6760
rect 6642 6160 6698 6216
rect 6918 3984 6974 4040
rect 6090 3032 6146 3088
rect 5906 2760 5962 2816
rect 6918 2896 6974 2952
rect 6918 2508 6974 2544
rect 6918 2488 6920 2508
rect 6920 2488 6972 2508
rect 6972 2488 6974 2508
rect 5262 1944 5318 2000
rect 7194 8608 7250 8664
rect 7378 8336 7434 8392
rect 8022 10920 8078 10976
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 10414 11600 10470 11656
rect 8206 11328 8262 11384
rect 8298 10648 8354 10704
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 8298 7384 8354 7440
rect 7470 6840 7526 6896
rect 8390 7148 8392 7168
rect 8392 7148 8444 7168
rect 8444 7148 8446 7168
rect 8390 7112 8446 7148
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 8390 6840 8446 6896
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7838 4684 7894 4720
rect 7838 4664 7840 4684
rect 7840 4664 7892 4684
rect 7892 4664 7894 4684
rect 8206 4528 8262 4584
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7378 3712 7434 3768
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 8114 2896 8170 2952
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 7010 1264 7066 1320
rect 9034 9968 9090 10024
rect 8666 7384 8722 7440
rect 8850 6604 8852 6624
rect 8852 6604 8904 6624
rect 8904 6604 8906 6624
rect 8850 6568 8906 6604
rect 9034 5752 9090 5808
rect 9034 4120 9090 4176
rect 8758 3476 8760 3496
rect 8760 3476 8812 3496
rect 8812 3476 8814 3496
rect 8758 3440 8814 3476
rect 9770 10240 9826 10296
rect 9586 8064 9642 8120
rect 10414 11056 10470 11112
rect 10046 9036 10102 9072
rect 10046 9016 10048 9036
rect 10048 9016 10100 9036
rect 10100 9016 10102 9036
rect 11242 11192 11298 11248
rect 10322 7928 10378 7984
rect 10598 9172 10654 9208
rect 10598 9152 10600 9172
rect 10600 9152 10652 9172
rect 10652 9152 10654 9172
rect 10690 9016 10746 9072
rect 10690 8200 10746 8256
rect 10690 7928 10746 7984
rect 9954 7248 10010 7304
rect 9862 7112 9918 7168
rect 9586 6860 9642 6896
rect 9586 6840 9588 6860
rect 9588 6840 9640 6860
rect 9640 6840 9642 6860
rect 10966 9152 11022 9208
rect 9954 6704 10010 6760
rect 10138 6704 10194 6760
rect 11702 9868 11704 9888
rect 11704 9868 11756 9888
rect 11756 9868 11758 9888
rect 11702 9832 11758 9868
rect 11978 11464 12034 11520
rect 12162 11500 12164 11520
rect 12164 11500 12216 11520
rect 12216 11500 12218 11520
rect 12162 11464 12218 11500
rect 11978 11192 12034 11248
rect 11886 9832 11942 9888
rect 11334 6296 11390 6352
rect 10138 6196 10140 6216
rect 10140 6196 10192 6216
rect 10192 6196 10194 6216
rect 10138 6160 10194 6196
rect 11242 6160 11298 6216
rect 10046 5652 10048 5672
rect 10048 5652 10100 5672
rect 10100 5652 10102 5672
rect 10046 5616 10102 5652
rect 9954 5208 10010 5264
rect 9770 4800 9826 4856
rect 9678 4664 9734 4720
rect 9770 4120 9826 4176
rect 9586 4004 9642 4040
rect 9586 3984 9588 4004
rect 9588 3984 9640 4004
rect 9640 3984 9642 4004
rect 10598 5072 10654 5128
rect 10230 3884 10232 3904
rect 10232 3884 10284 3904
rect 10284 3884 10286 3904
rect 10230 3848 10286 3884
rect 9494 2760 9550 2816
rect 10506 3440 10562 3496
rect 9402 2624 9458 2680
rect 11150 4120 11206 4176
rect 12530 9016 12586 9072
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 17038 12144 17094 12200
rect 12806 8064 12862 8120
rect 11702 4936 11758 4992
rect 11518 4664 11574 4720
rect 11886 4528 11942 4584
rect 11242 3984 11298 4040
rect 12530 5108 12532 5128
rect 12532 5108 12584 5128
rect 12584 5108 12586 5128
rect 12530 5072 12586 5108
rect 13266 9152 13322 9208
rect 13174 7656 13230 7712
rect 13082 5072 13138 5128
rect 12162 3576 12218 3632
rect 12990 3984 13046 4040
rect 13082 3712 13138 3768
rect 12622 3304 12678 3360
rect 12530 2896 12586 2952
rect 12806 3440 12862 3496
rect 11886 2388 11888 2408
rect 11888 2388 11940 2408
rect 11940 2388 11942 2408
rect 11886 2352 11942 2388
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 13450 7792 13506 7848
rect 13358 6568 13414 6624
rect 13726 7792 13782 7848
rect 13818 6296 13874 6352
rect 13818 4936 13874 4992
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14094 7384 14150 7440
rect 14554 7384 14610 7440
rect 14094 7112 14150 7168
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14738 7248 14794 7304
rect 15290 11600 15346 11656
rect 14830 6704 14886 6760
rect 14646 5072 14702 5128
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 13542 3576 13598 3632
rect 14738 4528 14794 4584
rect 18326 11736 18382 11792
rect 17130 11328 17186 11384
rect 15382 11056 15438 11112
rect 15382 9560 15438 9616
rect 15750 7520 15806 7576
rect 15382 5092 15438 5128
rect 15382 5072 15384 5092
rect 15384 5072 15436 5092
rect 15436 5072 15438 5092
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14922 3440 14978 3496
rect 13266 2644 13322 2680
rect 13266 2624 13268 2644
rect 13268 2624 13320 2644
rect 13320 2624 13322 2644
rect 14094 2896 14150 2952
rect 13910 2488 13966 2544
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 16302 9424 16358 9480
rect 16486 9288 16542 9344
rect 16486 7828 16488 7848
rect 16488 7828 16540 7848
rect 16540 7828 16542 7848
rect 16486 7792 16542 7828
rect 16854 7692 16856 7712
rect 16856 7692 16908 7712
rect 16908 7692 16910 7712
rect 16854 7656 16910 7692
rect 16854 6568 16910 6624
rect 15566 6024 15622 6080
rect 15658 5616 15714 5672
rect 17682 9424 17738 9480
rect 17038 5480 17094 5536
rect 16394 4936 16450 4992
rect 15750 4528 15806 4584
rect 15474 3576 15530 3632
rect 15750 3340 15752 3360
rect 15752 3340 15804 3360
rect 15804 3340 15806 3360
rect 15750 3304 15806 3340
rect 16026 3052 16082 3088
rect 16026 3032 16028 3052
rect 16028 3032 16080 3052
rect 16080 3032 16082 3052
rect 16946 3984 17002 4040
rect 16578 3032 16634 3088
rect 12898 2216 12954 2272
rect 14830 1944 14886 2000
rect 15566 2488 15622 2544
rect 17038 2624 17094 2680
rect 17958 9560 18014 9616
rect 17958 9016 18014 9072
rect 18050 8880 18106 8936
rect 18050 8472 18106 8528
rect 18234 9288 18290 9344
rect 18234 5244 18236 5264
rect 18236 5244 18288 5264
rect 18288 5244 18290 5264
rect 18234 5208 18290 5244
rect 18050 4936 18106 4992
rect 17774 4800 17830 4856
rect 18050 4120 18106 4176
rect 17866 3732 17922 3768
rect 17866 3712 17868 3732
rect 17868 3712 17920 3732
rect 17920 3712 17922 3732
rect 18510 11212 18566 11248
rect 18510 11192 18512 11212
rect 18512 11192 18564 11212
rect 18564 11192 18566 11212
rect 19338 10784 19394 10840
rect 18970 9696 19026 9752
rect 19338 8472 19394 8528
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 33322 12144 33378 12200
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 20718 11736 20774 11792
rect 19982 11328 20038 11384
rect 20074 11056 20130 11112
rect 19522 10668 19578 10704
rect 19522 10648 19524 10668
rect 19524 10648 19576 10668
rect 19576 10648 19578 10668
rect 19062 5208 19118 5264
rect 20626 10920 20682 10976
rect 19798 10648 19854 10704
rect 19798 9832 19854 9888
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 25502 11192 25558 11248
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 22282 11056 22338 11112
rect 19982 8880 20038 8936
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20810 9560 20866 9616
rect 21454 9288 21510 9344
rect 19798 7248 19854 7304
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20074 6332 20076 6352
rect 20076 6332 20128 6352
rect 20128 6332 20130 6352
rect 20074 6296 20130 6332
rect 19338 5616 19394 5672
rect 18786 4020 18788 4040
rect 18788 4020 18840 4040
rect 18840 4020 18842 4040
rect 18786 3984 18842 4020
rect 19062 3596 19118 3632
rect 19062 3576 19064 3596
rect 19064 3576 19116 3596
rect 19116 3576 19118 3596
rect 18326 2932 18328 2952
rect 18328 2932 18380 2952
rect 18380 2932 18382 2952
rect 18326 2896 18382 2932
rect 19890 4700 19892 4720
rect 19892 4700 19944 4720
rect 19944 4700 19946 4720
rect 19890 4664 19946 4700
rect 18326 2524 18328 2544
rect 18328 2524 18380 2544
rect 18380 2524 18382 2544
rect 18326 2488 18382 2524
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 21638 6296 21694 6352
rect 21638 6060 21640 6080
rect 21640 6060 21692 6080
rect 21692 6060 21694 6080
rect 21638 6024 21694 6060
rect 21270 4800 21326 4856
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 21270 3032 21326 3088
rect 20902 2644 20958 2680
rect 21822 8064 21878 8120
rect 21822 6160 21878 6216
rect 20902 2624 20904 2644
rect 20904 2624 20956 2644
rect 20956 2624 20958 2644
rect 22374 9832 22430 9888
rect 22466 9460 22468 9480
rect 22468 9460 22520 9480
rect 22520 9460 22522 9480
rect 22466 9424 22522 9460
rect 23478 9288 23534 9344
rect 22834 8744 22890 8800
rect 23662 8084 23718 8120
rect 23662 8064 23664 8084
rect 23664 8064 23716 8084
rect 23716 8064 23718 8084
rect 22650 6840 22706 6896
rect 22834 6840 22890 6896
rect 22098 5244 22100 5264
rect 22100 5244 22152 5264
rect 22152 5244 22154 5264
rect 22098 5208 22154 5244
rect 23110 5480 23166 5536
rect 23110 4664 23166 4720
rect 23570 4664 23626 4720
rect 23938 9152 23994 9208
rect 24030 9016 24086 9072
rect 22006 3032 22062 3088
rect 20626 2524 20628 2544
rect 20628 2524 20680 2544
rect 20680 2524 20682 2544
rect 20626 2488 20682 2524
rect 21822 2488 21878 2544
rect 20074 2252 20076 2272
rect 20076 2252 20128 2272
rect 20128 2252 20130 2272
rect 20074 2216 20130 2252
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 22742 3304 22798 3360
rect 26238 10920 26294 10976
rect 25502 10784 25558 10840
rect 27526 11076 27582 11112
rect 27526 11056 27528 11076
rect 27528 11056 27580 11076
rect 27580 11056 27582 11076
rect 29366 11056 29422 11112
rect 27158 10648 27214 10704
rect 25686 10104 25742 10160
rect 24398 7520 24454 7576
rect 24398 6180 24454 6216
rect 24398 6160 24400 6180
rect 24400 6160 24452 6180
rect 24452 6160 24454 6180
rect 24122 3712 24178 3768
rect 24030 3476 24032 3496
rect 24032 3476 24084 3496
rect 24084 3476 24086 3496
rect 24030 3440 24086 3476
rect 24858 7268 24914 7304
rect 24858 7248 24860 7268
rect 24860 7248 24912 7268
rect 24912 7248 24914 7268
rect 25410 7792 25466 7848
rect 25962 7384 26018 7440
rect 24950 6860 25006 6896
rect 24950 6840 24952 6860
rect 24952 6840 25004 6860
rect 25004 6840 25006 6860
rect 24950 6432 25006 6488
rect 24582 4972 24584 4992
rect 24584 4972 24636 4992
rect 24636 4972 24638 4992
rect 24582 4936 24638 4972
rect 25318 5616 25374 5672
rect 26606 10512 26662 10568
rect 28170 10548 28172 10568
rect 28172 10548 28224 10568
rect 28224 10548 28226 10568
rect 28170 10512 28226 10548
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 26698 9968 26754 10024
rect 26238 9460 26240 9480
rect 26240 9460 26292 9480
rect 26292 9460 26294 9480
rect 26238 9424 26294 9460
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 28262 9424 28318 9480
rect 27434 7656 27490 7712
rect 28262 9152 28318 9208
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 28170 7384 28226 7440
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 26882 6704 26938 6760
rect 25410 5092 25466 5128
rect 25410 5072 25412 5092
rect 25412 5072 25464 5092
rect 25464 5072 25466 5092
rect 26974 5228 27030 5264
rect 26974 5208 26976 5228
rect 26976 5208 27028 5228
rect 27028 5208 27030 5228
rect 26882 4936 26938 4992
rect 24674 3848 24730 3904
rect 22650 2508 22706 2544
rect 22650 2488 22652 2508
rect 22652 2488 22704 2508
rect 22704 2488 22706 2508
rect 26790 4392 26846 4448
rect 26330 3884 26332 3904
rect 26332 3884 26384 3904
rect 26384 3884 26386 3904
rect 26330 3848 26386 3884
rect 25502 3340 25504 3360
rect 25504 3340 25556 3360
rect 25556 3340 25558 3360
rect 25502 3304 25558 3340
rect 26698 2508 26754 2544
rect 26698 2488 26700 2508
rect 26700 2488 26752 2508
rect 26752 2488 26754 2508
rect 25962 2252 25964 2272
rect 25964 2252 26016 2272
rect 26016 2252 26018 2272
rect 25962 2216 26018 2252
rect 27342 5616 27398 5672
rect 27066 2080 27122 2136
rect 26974 1944 27030 2000
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 28630 8880 28686 8936
rect 28446 5208 28502 5264
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 28078 3984 28134 4040
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 28906 9016 28962 9072
rect 29090 9016 29146 9072
rect 28998 6316 29054 6352
rect 28998 6296 29000 6316
rect 29000 6296 29052 6316
rect 29052 6296 29054 6316
rect 29274 5652 29276 5672
rect 29276 5652 29328 5672
rect 29328 5652 29330 5672
rect 29274 5616 29330 5652
rect 33414 10784 33470 10840
rect 32310 10648 32366 10704
rect 32586 9580 32642 9616
rect 32586 9560 32588 9580
rect 32588 9560 32640 9580
rect 32640 9560 32642 9580
rect 29826 9324 29828 9344
rect 29828 9324 29880 9344
rect 29880 9324 29882 9344
rect 29826 9288 29882 9324
rect 29458 7692 29460 7712
rect 29460 7692 29512 7712
rect 29512 7692 29514 7712
rect 29458 7656 29514 7692
rect 29826 7520 29882 7576
rect 29550 6160 29606 6216
rect 28814 4256 28870 4312
rect 28354 3848 28410 3904
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 27710 2508 27766 2544
rect 27710 2488 27712 2508
rect 27712 2488 27764 2508
rect 27764 2488 27766 2508
rect 27434 1400 27490 1456
rect 29458 2760 29514 2816
rect 29734 4120 29790 4176
rect 29826 2760 29882 2816
rect 30378 7928 30434 7984
rect 30194 3576 30250 3632
rect 29550 2488 29606 2544
rect 30378 4684 30434 4720
rect 30378 4664 30380 4684
rect 30380 4664 30432 4684
rect 30432 4664 30434 4684
rect 30746 7792 30802 7848
rect 32678 8336 32734 8392
rect 30562 4392 30618 4448
rect 30838 6452 30894 6488
rect 30838 6432 30840 6452
rect 30840 6432 30892 6452
rect 30892 6432 30894 6452
rect 31206 6024 31262 6080
rect 31206 5752 31262 5808
rect 32310 6296 32366 6352
rect 31574 4004 31630 4040
rect 31574 3984 31576 4004
rect 31576 3984 31628 4004
rect 31628 3984 31630 4004
rect 30838 3440 30894 3496
rect 32126 4120 32182 4176
rect 33690 9152 33746 9208
rect 33874 10240 33930 10296
rect 33874 9832 33930 9888
rect 34150 10920 34206 10976
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 35438 10648 35494 10704
rect 34702 10124 34758 10160
rect 34702 10104 34704 10124
rect 34704 10104 34756 10124
rect 34756 10104 34758 10124
rect 34058 9152 34114 9208
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 35438 10240 35494 10296
rect 34794 9832 34850 9888
rect 35162 9580 35218 9616
rect 35162 9560 35164 9580
rect 35164 9560 35216 9580
rect 35216 9560 35218 9580
rect 33782 8744 33838 8800
rect 33966 8608 34022 8664
rect 34886 9016 34942 9072
rect 33874 7948 33930 7984
rect 33874 7928 33876 7948
rect 33876 7928 33928 7948
rect 33928 7928 33930 7948
rect 33138 6060 33140 6080
rect 33140 6060 33192 6080
rect 33192 6060 33194 6080
rect 33138 6024 33194 6060
rect 33046 5908 33102 5944
rect 33046 5888 33048 5908
rect 33048 5888 33100 5908
rect 33100 5888 33102 5908
rect 33322 5208 33378 5264
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34150 7384 34206 7440
rect 35070 8336 35126 8392
rect 34886 7520 34942 7576
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 35438 9832 35494 9888
rect 35714 14592 35770 14648
rect 35622 13776 35678 13832
rect 35622 12008 35678 12064
rect 35622 11056 35678 11112
rect 36818 12824 36874 12880
rect 36266 10512 36322 10568
rect 36634 10240 36690 10296
rect 36450 9460 36452 9480
rect 36452 9460 36504 9480
rect 36504 9460 36506 9480
rect 36450 9424 36506 9460
rect 35898 9324 35900 9344
rect 35900 9324 35952 9344
rect 35952 9324 35954 9344
rect 35898 9288 35954 9324
rect 35254 6160 35310 6216
rect 32586 4548 32642 4584
rect 32586 4528 32588 4548
rect 32588 4528 32640 4548
rect 32640 4528 32642 4548
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 35254 3984 35310 4040
rect 34978 3168 35034 3224
rect 34058 2216 34114 2272
rect 33138 2080 33194 2136
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 35438 5788 35440 5808
rect 35440 5788 35492 5808
rect 35492 5788 35494 5808
rect 35438 5752 35494 5788
rect 35530 4800 35586 4856
rect 35806 5888 35862 5944
rect 35898 2388 35900 2408
rect 35900 2388 35952 2408
rect 35952 2388 35954 2408
rect 35898 2352 35954 2388
rect 35346 1264 35402 1320
rect 36634 9288 36690 9344
rect 36358 9152 36414 9208
rect 36266 7248 36322 7304
rect 36634 8472 36690 8528
rect 36542 7404 36598 7440
rect 36542 7384 36544 7404
rect 36544 7384 36596 7404
rect 36596 7384 36598 7404
rect 36542 6180 36598 6216
rect 36542 6160 36544 6180
rect 36544 6160 36596 6180
rect 36596 6160 36598 6180
rect 36358 4120 36414 4176
rect 37554 7248 37610 7304
rect 37186 5752 37242 5808
rect 37370 5208 37426 5264
rect 36450 3848 36506 3904
rect 37278 3168 37334 3224
rect 38014 3984 38070 4040
rect 39394 3032 39450 3088
rect 39394 2896 39450 2952
rect 38750 2624 38806 2680
rect 36082 448 36138 504
<< metal3 >>
rect 0 15602 480 15632
rect 1393 15602 1459 15605
rect 0 15600 1459 15602
rect 0 15544 1398 15600
rect 1454 15544 1459 15600
rect 0 15542 1459 15544
rect 0 15512 480 15542
rect 1393 15539 1459 15542
rect 35525 15602 35591 15605
rect 39520 15602 40000 15632
rect 35525 15600 40000 15602
rect 35525 15544 35530 15600
rect 35586 15544 40000 15600
rect 35525 15542 40000 15544
rect 35525 15539 35591 15542
rect 39520 15512 40000 15542
rect 0 14650 480 14680
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 480 14590
rect 1485 14587 1551 14590
rect 35709 14650 35775 14653
rect 39520 14650 40000 14680
rect 35709 14648 40000 14650
rect 35709 14592 35714 14648
rect 35770 14592 40000 14648
rect 35709 14590 40000 14592
rect 35709 14587 35775 14590
rect 39520 14560 40000 14590
rect 0 13834 480 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 480 13774
rect 1577 13771 1643 13774
rect 35617 13834 35683 13837
rect 39520 13834 40000 13864
rect 35617 13832 40000 13834
rect 35617 13776 35622 13832
rect 35678 13776 40000 13832
rect 35617 13774 40000 13776
rect 35617 13771 35683 13774
rect 39520 13744 40000 13774
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12882 480 12912
rect 2957 12882 3023 12885
rect 0 12880 3023 12882
rect 0 12824 2962 12880
rect 3018 12824 3023 12880
rect 0 12822 3023 12824
rect 0 12792 480 12822
rect 2957 12819 3023 12822
rect 36813 12882 36879 12885
rect 39520 12882 40000 12912
rect 36813 12880 40000 12882
rect 36813 12824 36818 12880
rect 36874 12824 40000 12880
rect 36813 12822 40000 12824
rect 36813 12819 36879 12822
rect 39520 12792 40000 12822
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 17033 12202 17099 12205
rect 33317 12202 33383 12205
rect 17033 12200 33383 12202
rect 17033 12144 17038 12200
rect 17094 12144 33322 12200
rect 33378 12144 33383 12200
rect 17033 12142 33383 12144
rect 17033 12139 17099 12142
rect 33317 12139 33383 12142
rect 0 12066 480 12096
rect 4061 12066 4127 12069
rect 0 12064 4127 12066
rect 0 12008 4066 12064
rect 4122 12008 4127 12064
rect 0 12006 4127 12008
rect 0 11976 480 12006
rect 4061 12003 4127 12006
rect 35617 12066 35683 12069
rect 39520 12066 40000 12096
rect 35617 12064 40000 12066
rect 35617 12008 35622 12064
rect 35678 12008 40000 12064
rect 35617 12006 40000 12008
rect 35617 12003 35683 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12006
rect 34277 11935 34597 11936
rect 3969 11794 4035 11797
rect 5441 11794 5507 11797
rect 18321 11794 18387 11797
rect 20713 11794 20779 11797
rect 3969 11792 20779 11794
rect 3969 11736 3974 11792
rect 4030 11736 5446 11792
rect 5502 11736 18326 11792
rect 18382 11736 20718 11792
rect 20774 11736 20779 11792
rect 3969 11734 20779 11736
rect 3969 11731 4035 11734
rect 5441 11731 5507 11734
rect 18321 11731 18387 11734
rect 20713 11731 20779 11734
rect 6177 11658 6243 11661
rect 10409 11658 10475 11661
rect 15285 11658 15351 11661
rect 6177 11656 10242 11658
rect 6177 11600 6182 11656
rect 6238 11600 10242 11656
rect 6177 11598 10242 11600
rect 6177 11595 6243 11598
rect 1669 11522 1735 11525
rect 7097 11522 7163 11525
rect 1669 11520 7163 11522
rect 1669 11464 1674 11520
rect 1730 11464 7102 11520
rect 7158 11464 7163 11520
rect 1669 11462 7163 11464
rect 10182 11522 10242 11598
rect 10409 11656 15351 11658
rect 10409 11600 10414 11656
rect 10470 11600 15290 11656
rect 15346 11600 15351 11656
rect 10409 11598 15351 11600
rect 10409 11595 10475 11598
rect 15285 11595 15351 11598
rect 11973 11522 12039 11525
rect 12157 11524 12223 11525
rect 12157 11522 12204 11524
rect 10182 11520 12039 11522
rect 10182 11464 11978 11520
rect 12034 11464 12039 11520
rect 10182 11462 12039 11464
rect 12112 11520 12204 11522
rect 12112 11464 12162 11520
rect 12112 11462 12204 11464
rect 1669 11459 1735 11462
rect 7097 11459 7163 11462
rect 11973 11459 12039 11462
rect 12157 11460 12204 11462
rect 12268 11460 12274 11524
rect 12157 11459 12223 11460
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 3325 11386 3391 11389
rect 8201 11386 8267 11389
rect 3325 11384 8267 11386
rect 3325 11328 3330 11384
rect 3386 11328 8206 11384
rect 8262 11328 8267 11384
rect 3325 11326 8267 11328
rect 3325 11323 3391 11326
rect 8201 11323 8267 11326
rect 17125 11386 17191 11389
rect 19977 11386 20043 11389
rect 17125 11384 20043 11386
rect 17125 11328 17130 11384
rect 17186 11328 19982 11384
rect 20038 11328 20043 11384
rect 17125 11326 20043 11328
rect 17125 11323 17191 11326
rect 19977 11323 20043 11326
rect 4889 11250 4955 11253
rect 11237 11252 11303 11253
rect 11237 11250 11284 11252
rect 4889 11248 11284 11250
rect 11348 11250 11354 11252
rect 11973 11250 12039 11253
rect 18505 11250 18571 11253
rect 25497 11250 25563 11253
rect 4889 11192 4894 11248
rect 4950 11192 11242 11248
rect 4889 11190 11284 11192
rect 4889 11187 4955 11190
rect 11237 11188 11284 11190
rect 11348 11190 11430 11250
rect 11973 11248 25563 11250
rect 11973 11192 11978 11248
rect 12034 11192 18510 11248
rect 18566 11192 25502 11248
rect 25558 11192 25563 11248
rect 11973 11190 25563 11192
rect 11348 11188 11354 11190
rect 11237 11187 11303 11188
rect 11973 11187 12039 11190
rect 18505 11187 18571 11190
rect 25497 11187 25563 11190
rect 0 11114 480 11144
rect 2681 11114 2747 11117
rect 0 11112 2747 11114
rect 0 11056 2686 11112
rect 2742 11056 2747 11112
rect 0 11054 2747 11056
rect 0 11024 480 11054
rect 2681 11051 2747 11054
rect 4797 11114 4863 11117
rect 6913 11114 6979 11117
rect 4797 11112 6979 11114
rect 4797 11056 4802 11112
rect 4858 11056 6918 11112
rect 6974 11056 6979 11112
rect 4797 11054 6979 11056
rect 4797 11051 4863 11054
rect 6913 11051 6979 11054
rect 10409 11114 10475 11117
rect 15377 11114 15443 11117
rect 10409 11112 15443 11114
rect 10409 11056 10414 11112
rect 10470 11056 15382 11112
rect 15438 11056 15443 11112
rect 10409 11054 15443 11056
rect 10409 11051 10475 11054
rect 15377 11051 15443 11054
rect 20069 11114 20135 11117
rect 22277 11114 22343 11117
rect 20069 11112 22343 11114
rect 20069 11056 20074 11112
rect 20130 11056 22282 11112
rect 22338 11056 22343 11112
rect 20069 11054 22343 11056
rect 20069 11051 20135 11054
rect 22277 11051 22343 11054
rect 27521 11114 27587 11117
rect 29361 11114 29427 11117
rect 27521 11112 29427 11114
rect 27521 11056 27526 11112
rect 27582 11056 29366 11112
rect 29422 11056 29427 11112
rect 27521 11054 29427 11056
rect 27521 11051 27587 11054
rect 29361 11051 29427 11054
rect 35617 11114 35683 11117
rect 39520 11114 40000 11144
rect 35617 11112 40000 11114
rect 35617 11056 35622 11112
rect 35678 11056 40000 11112
rect 35617 11054 40000 11056
rect 35617 11051 35683 11054
rect 39520 11024 40000 11054
rect 3417 10978 3483 10981
rect 7005 10978 7071 10981
rect 3417 10976 7071 10978
rect 3417 10920 3422 10976
rect 3478 10920 7010 10976
rect 7066 10920 7071 10976
rect 3417 10918 7071 10920
rect 3417 10915 3483 10918
rect 7005 10915 7071 10918
rect 8017 10978 8083 10981
rect 20621 10978 20687 10981
rect 8017 10976 20687 10978
rect 8017 10920 8022 10976
rect 8078 10920 20626 10976
rect 20682 10920 20687 10976
rect 8017 10918 20687 10920
rect 8017 10915 8083 10918
rect 20621 10915 20687 10918
rect 26233 10978 26299 10981
rect 34145 10978 34211 10981
rect 26233 10976 34211 10978
rect 26233 10920 26238 10976
rect 26294 10920 34150 10976
rect 34206 10920 34211 10976
rect 26233 10918 34211 10920
rect 26233 10915 26299 10918
rect 34145 10915 34211 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 19333 10842 19399 10845
rect 8158 10840 19399 10842
rect 8158 10784 19338 10840
rect 19394 10784 19399 10840
rect 8158 10782 19399 10784
rect 4245 10706 4311 10709
rect 8158 10706 8218 10782
rect 19333 10779 19399 10782
rect 25497 10842 25563 10845
rect 33409 10842 33475 10845
rect 25497 10840 33475 10842
rect 25497 10784 25502 10840
rect 25558 10784 33414 10840
rect 33470 10784 33475 10840
rect 25497 10782 33475 10784
rect 25497 10779 25563 10782
rect 33409 10779 33475 10782
rect 4245 10704 8218 10706
rect 4245 10648 4250 10704
rect 4306 10648 8218 10704
rect 4245 10646 8218 10648
rect 8293 10706 8359 10709
rect 19517 10706 19583 10709
rect 8293 10704 19583 10706
rect 8293 10648 8298 10704
rect 8354 10648 19522 10704
rect 19578 10648 19583 10704
rect 8293 10646 19583 10648
rect 4245 10643 4311 10646
rect 8293 10643 8359 10646
rect 19517 10643 19583 10646
rect 19793 10706 19859 10709
rect 27153 10706 27219 10709
rect 32305 10706 32371 10709
rect 35433 10706 35499 10709
rect 19793 10704 26986 10706
rect 19793 10648 19798 10704
rect 19854 10648 26986 10704
rect 19793 10646 26986 10648
rect 19793 10643 19859 10646
rect 5533 10570 5599 10573
rect 6453 10570 6519 10573
rect 26601 10570 26667 10573
rect 5533 10568 26667 10570
rect 5533 10512 5538 10568
rect 5594 10512 6458 10568
rect 6514 10512 26606 10568
rect 26662 10512 26667 10568
rect 5533 10510 26667 10512
rect 5533 10507 5599 10510
rect 6453 10507 6519 10510
rect 26601 10507 26667 10510
rect 2037 10434 2103 10437
rect 5717 10434 5783 10437
rect 2037 10432 5783 10434
rect 2037 10376 2042 10432
rect 2098 10376 5722 10432
rect 5778 10376 5783 10432
rect 2037 10374 5783 10376
rect 2037 10371 2103 10374
rect 5717 10371 5783 10374
rect 14277 10368 14597 10369
rect 0 10298 480 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 3601 10298 3667 10301
rect 0 10296 3667 10298
rect 0 10240 3606 10296
rect 3662 10240 3667 10296
rect 0 10238 3667 10240
rect 0 10208 480 10238
rect 3601 10235 3667 10238
rect 7189 10298 7255 10301
rect 9765 10298 9831 10301
rect 7189 10296 9831 10298
rect 7189 10240 7194 10296
rect 7250 10240 9770 10296
rect 9826 10240 9831 10296
rect 7189 10238 9831 10240
rect 7189 10235 7255 10238
rect 9765 10235 9831 10238
rect 3049 10162 3115 10165
rect 25681 10162 25747 10165
rect 3049 10160 25747 10162
rect 3049 10104 3054 10160
rect 3110 10104 25686 10160
rect 25742 10104 25747 10160
rect 3049 10102 25747 10104
rect 26926 10162 26986 10646
rect 27153 10704 35499 10706
rect 27153 10648 27158 10704
rect 27214 10648 32310 10704
rect 32366 10648 35438 10704
rect 35494 10648 35499 10704
rect 27153 10646 35499 10648
rect 27153 10643 27219 10646
rect 32305 10643 32371 10646
rect 35433 10643 35499 10646
rect 28165 10572 28231 10573
rect 28165 10570 28212 10572
rect 28120 10568 28212 10570
rect 28276 10570 28282 10572
rect 36261 10570 36327 10573
rect 28276 10568 36327 10570
rect 28120 10512 28170 10568
rect 28276 10512 36266 10568
rect 36322 10512 36327 10568
rect 28120 10510 28212 10512
rect 28165 10508 28212 10510
rect 28276 10510 36327 10512
rect 28276 10508 28282 10510
rect 28165 10507 28231 10508
rect 36261 10507 36327 10510
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 33869 10298 33935 10301
rect 35433 10298 35499 10301
rect 33869 10296 35499 10298
rect 33869 10240 33874 10296
rect 33930 10240 35438 10296
rect 35494 10240 35499 10296
rect 33869 10238 35499 10240
rect 33869 10235 33935 10238
rect 35433 10235 35499 10238
rect 36629 10298 36695 10301
rect 39520 10298 40000 10328
rect 36629 10296 40000 10298
rect 36629 10240 36634 10296
rect 36690 10240 40000 10296
rect 36629 10238 40000 10240
rect 36629 10235 36695 10238
rect 39520 10208 40000 10238
rect 34697 10162 34763 10165
rect 26926 10160 34763 10162
rect 26926 10104 34702 10160
rect 34758 10104 34763 10160
rect 26926 10102 34763 10104
rect 3049 10099 3115 10102
rect 25681 10099 25747 10102
rect 34697 10099 34763 10102
rect 5165 10026 5231 10029
rect 9029 10026 9095 10029
rect 26693 10026 26759 10029
rect 5165 10024 8218 10026
rect 5165 9968 5170 10024
rect 5226 9968 8218 10024
rect 5165 9966 8218 9968
rect 5165 9963 5231 9966
rect 3325 9890 3391 9893
rect 7189 9890 7255 9893
rect 3325 9888 7255 9890
rect 3325 9832 3330 9888
rect 3386 9832 7194 9888
rect 7250 9832 7255 9888
rect 3325 9830 7255 9832
rect 3325 9827 3391 9830
rect 7189 9827 7255 9830
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 8158 9754 8218 9966
rect 9029 10024 26759 10026
rect 9029 9968 9034 10024
rect 9090 9968 26698 10024
rect 26754 9968 26759 10024
rect 9029 9966 26759 9968
rect 9029 9963 9095 9966
rect 26693 9963 26759 9966
rect 11697 9892 11763 9893
rect 11646 9890 11652 9892
rect 11606 9830 11652 9890
rect 11716 9888 11763 9892
rect 11758 9832 11763 9888
rect 11646 9828 11652 9830
rect 11716 9828 11763 9832
rect 11697 9827 11763 9828
rect 11881 9890 11947 9893
rect 19793 9890 19859 9893
rect 11881 9888 19859 9890
rect 11881 9832 11886 9888
rect 11942 9832 19798 9888
rect 19854 9832 19859 9888
rect 11881 9830 19859 9832
rect 11881 9827 11947 9830
rect 19793 9827 19859 9830
rect 22369 9890 22435 9893
rect 33869 9890 33935 9893
rect 22369 9888 33935 9890
rect 22369 9832 22374 9888
rect 22430 9832 33874 9888
rect 33930 9832 33935 9888
rect 22369 9830 33935 9832
rect 22369 9827 22435 9830
rect 33869 9827 33935 9830
rect 34789 9890 34855 9893
rect 35433 9890 35499 9893
rect 34789 9888 35499 9890
rect 34789 9832 34794 9888
rect 34850 9832 35438 9888
rect 35494 9832 35499 9888
rect 34789 9830 35499 9832
rect 34789 9827 34855 9830
rect 35433 9827 35499 9830
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 18965 9754 19031 9757
rect 8158 9752 19031 9754
rect 8158 9696 18970 9752
rect 19026 9696 19031 9752
rect 8158 9694 19031 9696
rect 18965 9691 19031 9694
rect 15377 9618 15443 9621
rect 17953 9618 18019 9621
rect 9584 9584 12266 9618
rect 12390 9584 14796 9618
rect 9584 9558 14796 9584
rect 9584 9516 9644 9558
rect 12206 9524 12450 9558
rect 3693 9482 3759 9485
rect 7097 9482 7163 9485
rect 3693 9480 7163 9482
rect 3693 9424 3698 9480
rect 3754 9424 7102 9480
rect 7158 9424 7163 9480
rect 3693 9422 7163 9424
rect 3693 9419 3759 9422
rect 7097 9419 7163 9422
rect 9446 9456 9644 9516
rect 0 9346 480 9376
rect 4337 9346 4403 9349
rect 0 9344 4403 9346
rect 0 9288 4342 9344
rect 4398 9288 4403 9344
rect 0 9286 4403 9288
rect 0 9256 480 9286
rect 4337 9283 4403 9286
rect 5901 9346 5967 9349
rect 9446 9346 9506 9456
rect 5901 9344 9506 9346
rect 5901 9288 5906 9344
rect 5962 9288 9506 9344
rect 5901 9286 9506 9288
rect 5901 9283 5967 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 3877 9210 3943 9213
rect 4245 9210 4311 9213
rect 7005 9210 7071 9213
rect 10593 9210 10659 9213
rect 3877 9208 10659 9210
rect 3877 9152 3882 9208
rect 3938 9152 4250 9208
rect 4306 9152 7010 9208
rect 7066 9152 10598 9208
rect 10654 9152 10659 9208
rect 3877 9150 10659 9152
rect 3877 9147 3943 9150
rect 4245 9147 4311 9150
rect 7005 9147 7071 9150
rect 10593 9147 10659 9150
rect 10961 9210 11027 9213
rect 13261 9210 13327 9213
rect 10961 9208 13327 9210
rect 10961 9152 10966 9208
rect 11022 9152 13266 9208
rect 13322 9152 13327 9208
rect 10961 9150 13327 9152
rect 14736 9210 14796 9558
rect 15377 9616 18019 9618
rect 15377 9560 15382 9616
rect 15438 9560 17958 9616
rect 18014 9560 18019 9616
rect 15377 9558 18019 9560
rect 15377 9555 15443 9558
rect 17953 9555 18019 9558
rect 20805 9618 20871 9621
rect 32581 9618 32647 9621
rect 35157 9618 35223 9621
rect 20805 9616 35223 9618
rect 20805 9560 20810 9616
rect 20866 9560 32586 9616
rect 32642 9560 35162 9616
rect 35218 9560 35223 9616
rect 20805 9558 35223 9560
rect 20805 9555 20871 9558
rect 32581 9555 32647 9558
rect 35157 9555 35223 9558
rect 16297 9482 16363 9485
rect 17677 9482 17743 9485
rect 16297 9480 17743 9482
rect 16297 9424 16302 9480
rect 16358 9424 17682 9480
rect 17738 9424 17743 9480
rect 16297 9422 17743 9424
rect 16297 9419 16363 9422
rect 17677 9419 17743 9422
rect 22461 9482 22527 9485
rect 26233 9482 26299 9485
rect 22461 9480 26299 9482
rect 22461 9424 22466 9480
rect 22522 9424 26238 9480
rect 26294 9424 26299 9480
rect 22461 9422 26299 9424
rect 22461 9419 22527 9422
rect 26233 9419 26299 9422
rect 28257 9482 28323 9485
rect 36445 9482 36511 9485
rect 28257 9480 36511 9482
rect 28257 9424 28262 9480
rect 28318 9424 36450 9480
rect 36506 9424 36511 9480
rect 28257 9422 36511 9424
rect 28257 9419 28323 9422
rect 36445 9419 36511 9422
rect 16481 9346 16547 9349
rect 18229 9346 18295 9349
rect 16481 9344 18295 9346
rect 16481 9288 16486 9344
rect 16542 9288 18234 9344
rect 18290 9288 18295 9344
rect 16481 9286 18295 9288
rect 16481 9283 16547 9286
rect 18229 9283 18295 9286
rect 21449 9346 21515 9349
rect 23473 9346 23539 9349
rect 21449 9344 23539 9346
rect 21449 9288 21454 9344
rect 21510 9288 23478 9344
rect 23534 9288 23539 9344
rect 21449 9286 23539 9288
rect 21449 9283 21515 9286
rect 23473 9283 23539 9286
rect 29821 9346 29887 9349
rect 35893 9346 35959 9349
rect 29821 9344 35959 9346
rect 29821 9288 29826 9344
rect 29882 9288 35898 9344
rect 35954 9288 35959 9344
rect 29821 9286 35959 9288
rect 29821 9283 29887 9286
rect 35893 9283 35959 9286
rect 36629 9346 36695 9349
rect 39520 9346 40000 9376
rect 36629 9344 40000 9346
rect 36629 9288 36634 9344
rect 36690 9288 40000 9344
rect 36629 9286 40000 9288
rect 36629 9283 36695 9286
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9286
rect 27610 9215 27930 9216
rect 23933 9210 23999 9213
rect 28257 9212 28323 9213
rect 14736 9208 23999 9210
rect 14736 9152 23938 9208
rect 23994 9152 23999 9208
rect 14736 9150 23999 9152
rect 10961 9147 11027 9150
rect 13261 9147 13327 9150
rect 23933 9147 23999 9150
rect 28206 9148 28212 9212
rect 28276 9210 28323 9212
rect 28276 9208 28368 9210
rect 28318 9152 28368 9208
rect 28276 9150 28368 9152
rect 28276 9148 28323 9150
rect 28942 9148 28948 9212
rect 29012 9210 29018 9212
rect 33685 9210 33751 9213
rect 29012 9208 33751 9210
rect 29012 9152 33690 9208
rect 33746 9152 33751 9208
rect 29012 9150 33751 9152
rect 29012 9148 29018 9150
rect 28257 9147 28323 9148
rect 33685 9147 33751 9150
rect 34053 9210 34119 9213
rect 36353 9210 36419 9213
rect 34053 9208 36419 9210
rect 34053 9152 34058 9208
rect 34114 9152 36358 9208
rect 36414 9152 36419 9208
rect 34053 9150 36419 9152
rect 34053 9147 34119 9150
rect 36353 9147 36419 9150
rect 6545 9074 6611 9077
rect 10041 9074 10107 9077
rect 6545 9072 10107 9074
rect 6545 9016 6550 9072
rect 6606 9016 10046 9072
rect 10102 9016 10107 9072
rect 6545 9014 10107 9016
rect 6545 9011 6611 9014
rect 10041 9011 10107 9014
rect 10685 9074 10751 9077
rect 12525 9074 12591 9077
rect 10685 9072 12591 9074
rect 10685 9016 10690 9072
rect 10746 9016 12530 9072
rect 12586 9016 12591 9072
rect 10685 9014 12591 9016
rect 10685 9011 10751 9014
rect 12525 9011 12591 9014
rect 17953 9074 18019 9077
rect 24025 9074 24091 9077
rect 17953 9072 24091 9074
rect 17953 9016 17958 9072
rect 18014 9016 24030 9072
rect 24086 9016 24091 9072
rect 17953 9014 24091 9016
rect 17953 9011 18019 9014
rect 24025 9011 24091 9014
rect 28901 9074 28967 9077
rect 29085 9074 29151 9077
rect 34881 9074 34947 9077
rect 28901 9072 29151 9074
rect 28901 9016 28906 9072
rect 28962 9016 29090 9072
rect 29146 9016 29151 9072
rect 28901 9014 29151 9016
rect 28901 9011 28967 9014
rect 29085 9011 29151 9014
rect 34102 9072 34947 9074
rect 34102 9016 34886 9072
rect 34942 9016 34947 9072
rect 34102 9014 34947 9016
rect 2129 8938 2195 8941
rect 4429 8938 4495 8941
rect 2129 8936 4495 8938
rect 2129 8880 2134 8936
rect 2190 8880 4434 8936
rect 4490 8880 4495 8936
rect 2129 8878 4495 8880
rect 2129 8875 2195 8878
rect 4429 8875 4495 8878
rect 5717 8938 5783 8941
rect 18045 8938 18111 8941
rect 5717 8936 18111 8938
rect 5717 8880 5722 8936
rect 5778 8880 18050 8936
rect 18106 8880 18111 8936
rect 5717 8878 18111 8880
rect 5717 8875 5783 8878
rect 18045 8875 18111 8878
rect 19977 8938 20043 8941
rect 28625 8938 28691 8941
rect 28942 8938 28948 8940
rect 19977 8936 21466 8938
rect 19977 8880 19982 8936
rect 20038 8880 21466 8936
rect 19977 8878 21466 8880
rect 19977 8875 20043 8878
rect 2313 8802 2379 8805
rect 6545 8802 6611 8805
rect 2313 8800 6611 8802
rect 2313 8744 2318 8800
rect 2374 8744 6550 8800
rect 6606 8744 6611 8800
rect 2313 8742 6611 8744
rect 2313 8739 2379 8742
rect 6545 8739 6611 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 2497 8666 2563 8669
rect 7189 8666 7255 8669
rect 2497 8664 7255 8666
rect 2497 8608 2502 8664
rect 2558 8608 7194 8664
rect 7250 8608 7255 8664
rect 2497 8606 7255 8608
rect 21406 8666 21466 8878
rect 28625 8936 28948 8938
rect 28625 8880 28630 8936
rect 28686 8880 28948 8936
rect 28625 8878 28948 8880
rect 28625 8875 28691 8878
rect 28942 8876 28948 8878
rect 29012 8876 29018 8940
rect 22829 8802 22895 8805
rect 33777 8802 33843 8805
rect 34102 8802 34162 9014
rect 34881 9011 34947 9014
rect 22829 8800 34162 8802
rect 22829 8744 22834 8800
rect 22890 8744 33782 8800
rect 33838 8744 34162 8800
rect 22829 8742 34162 8744
rect 22829 8739 22895 8742
rect 33777 8739 33843 8742
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 33961 8666 34027 8669
rect 21406 8664 34027 8666
rect 21406 8608 33966 8664
rect 34022 8608 34027 8664
rect 21406 8606 34027 8608
rect 2497 8603 2563 8606
rect 7189 8603 7255 8606
rect 33961 8603 34027 8606
rect 0 8530 480 8560
rect 565 8530 631 8533
rect 0 8528 631 8530
rect 0 8472 570 8528
rect 626 8472 631 8528
rect 0 8470 631 8472
rect 0 8440 480 8470
rect 565 8467 631 8470
rect 3049 8530 3115 8533
rect 5533 8530 5599 8533
rect 3049 8528 5599 8530
rect 3049 8472 3054 8528
rect 3110 8472 5538 8528
rect 5594 8472 5599 8528
rect 3049 8470 5599 8472
rect 3049 8467 3115 8470
rect 5533 8467 5599 8470
rect 18045 8530 18111 8533
rect 19333 8530 19399 8533
rect 18045 8528 19399 8530
rect 18045 8472 18050 8528
rect 18106 8472 19338 8528
rect 19394 8472 19399 8528
rect 18045 8470 19399 8472
rect 18045 8467 18111 8470
rect 19333 8467 19399 8470
rect 36629 8530 36695 8533
rect 39520 8530 40000 8560
rect 36629 8528 40000 8530
rect 36629 8472 36634 8528
rect 36690 8472 40000 8528
rect 36629 8470 40000 8472
rect 36629 8467 36695 8470
rect 39520 8440 40000 8470
rect 3785 8394 3851 8397
rect 4705 8394 4771 8397
rect 3785 8392 4771 8394
rect 3785 8336 3790 8392
rect 3846 8336 4710 8392
rect 4766 8336 4771 8392
rect 3785 8334 4771 8336
rect 3785 8331 3851 8334
rect 4705 8331 4771 8334
rect 7005 8394 7071 8397
rect 7373 8394 7439 8397
rect 7005 8392 7439 8394
rect 7005 8336 7010 8392
rect 7066 8336 7378 8392
rect 7434 8336 7439 8392
rect 7005 8334 7439 8336
rect 7005 8331 7071 8334
rect 7373 8331 7439 8334
rect 32673 8394 32739 8397
rect 35065 8394 35131 8397
rect 32673 8392 35131 8394
rect 32673 8336 32678 8392
rect 32734 8336 35070 8392
rect 35126 8336 35131 8392
rect 32673 8334 35131 8336
rect 32673 8331 32739 8334
rect 35065 8331 35131 8334
rect 10685 8258 10751 8261
rect 9446 8256 10751 8258
rect 9446 8200 10690 8256
rect 10746 8200 10751 8256
rect 9446 8198 10751 8200
rect 3601 8122 3667 8125
rect 9446 8122 9506 8198
rect 10685 8195 10751 8198
rect 17174 8198 27538 8258
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 3601 8120 9506 8122
rect 3601 8064 3606 8120
rect 3662 8064 9506 8120
rect 3601 8062 9506 8064
rect 9581 8122 9647 8125
rect 12801 8122 12867 8125
rect 9581 8120 12867 8122
rect 9581 8064 9586 8120
rect 9642 8064 12806 8120
rect 12862 8064 12867 8120
rect 9581 8062 12867 8064
rect 3601 8059 3667 8062
rect 9581 8059 9647 8062
rect 12801 8059 12867 8062
rect 4521 7986 4587 7989
rect 10317 7986 10383 7989
rect 4521 7984 10383 7986
rect 4521 7928 4526 7984
rect 4582 7928 10322 7984
rect 10378 7928 10383 7984
rect 4521 7926 10383 7928
rect 4521 7923 4587 7926
rect 10317 7923 10383 7926
rect 10685 7986 10751 7989
rect 17174 7986 17234 8198
rect 21817 8122 21883 8125
rect 23657 8122 23723 8125
rect 21817 8120 23723 8122
rect 21817 8064 21822 8120
rect 21878 8064 23662 8120
rect 23718 8064 23723 8120
rect 21817 8062 23723 8064
rect 21817 8059 21883 8062
rect 23657 8059 23723 8062
rect 10685 7984 17234 7986
rect 10685 7928 10690 7984
rect 10746 7928 17234 7984
rect 10685 7926 17234 7928
rect 27478 7986 27538 8198
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 30373 7986 30439 7989
rect 33869 7986 33935 7989
rect 27478 7984 33935 7986
rect 27478 7928 30378 7984
rect 30434 7928 33874 7984
rect 33930 7928 33935 7984
rect 27478 7926 33935 7928
rect 10685 7923 10751 7926
rect 30373 7923 30439 7926
rect 33869 7923 33935 7926
rect 6269 7850 6335 7853
rect 13445 7850 13511 7853
rect 6269 7848 13511 7850
rect 6269 7792 6274 7848
rect 6330 7792 13450 7848
rect 13506 7792 13511 7848
rect 6269 7790 13511 7792
rect 6269 7787 6335 7790
rect 13445 7787 13511 7790
rect 13721 7850 13787 7853
rect 16481 7850 16547 7853
rect 13721 7848 16547 7850
rect 13721 7792 13726 7848
rect 13782 7792 16486 7848
rect 16542 7792 16547 7848
rect 13721 7790 16547 7792
rect 13721 7787 13787 7790
rect 16481 7787 16547 7790
rect 25405 7850 25471 7853
rect 30741 7850 30807 7853
rect 25405 7848 30807 7850
rect 25405 7792 25410 7848
rect 25466 7792 30746 7848
rect 30802 7792 30807 7848
rect 25405 7790 30807 7792
rect 25405 7787 25471 7790
rect 30741 7787 30807 7790
rect 5349 7714 5415 7717
rect 6913 7714 6979 7717
rect 5349 7712 6979 7714
rect 5349 7656 5354 7712
rect 5410 7656 6918 7712
rect 6974 7656 6979 7712
rect 5349 7654 6979 7656
rect 5349 7651 5415 7654
rect 6913 7651 6979 7654
rect 13169 7714 13235 7717
rect 16849 7714 16915 7717
rect 13169 7712 16915 7714
rect 13169 7656 13174 7712
rect 13230 7656 16854 7712
rect 16910 7656 16915 7712
rect 13169 7654 16915 7656
rect 13169 7651 13235 7654
rect 16849 7651 16915 7654
rect 27429 7714 27495 7717
rect 29453 7714 29519 7717
rect 27429 7712 29519 7714
rect 27429 7656 27434 7712
rect 27490 7656 29458 7712
rect 29514 7656 29519 7712
rect 27429 7654 29519 7656
rect 27429 7651 27495 7654
rect 29453 7651 29519 7654
rect 7610 7648 7930 7649
rect 0 7578 480 7608
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 4061 7578 4127 7581
rect 15745 7578 15811 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 480 7518
rect 4061 7515 4127 7518
rect 14414 7576 15811 7578
rect 14414 7520 15750 7576
rect 15806 7520 15811 7576
rect 14414 7518 15811 7520
rect 6821 7442 6887 7445
rect 8293 7442 8359 7445
rect 6821 7440 8359 7442
rect 6821 7384 6826 7440
rect 6882 7384 8298 7440
rect 8354 7384 8359 7440
rect 6821 7382 8359 7384
rect 6821 7379 6887 7382
rect 8293 7379 8359 7382
rect 8661 7442 8727 7445
rect 14089 7442 14155 7445
rect 14414 7442 14474 7518
rect 15745 7515 15811 7518
rect 24393 7578 24459 7581
rect 29821 7578 29887 7581
rect 24393 7576 29887 7578
rect 24393 7520 24398 7576
rect 24454 7520 29826 7576
rect 29882 7520 29887 7576
rect 24393 7518 29887 7520
rect 24393 7515 24459 7518
rect 29821 7515 29887 7518
rect 34881 7578 34947 7581
rect 39520 7578 40000 7608
rect 34881 7576 40000 7578
rect 34881 7520 34886 7576
rect 34942 7520 40000 7576
rect 34881 7518 40000 7520
rect 34881 7515 34947 7518
rect 39520 7488 40000 7518
rect 8661 7440 14474 7442
rect 8661 7384 8666 7440
rect 8722 7384 14094 7440
rect 14150 7384 14474 7440
rect 8661 7382 14474 7384
rect 14549 7442 14615 7445
rect 25957 7442 26023 7445
rect 28165 7442 28231 7445
rect 14549 7440 15946 7442
rect 14549 7384 14554 7440
rect 14610 7384 15946 7440
rect 14549 7382 15946 7384
rect 8661 7379 8727 7382
rect 14089 7379 14155 7382
rect 14549 7379 14615 7382
rect 9949 7306 10015 7309
rect 14733 7306 14799 7309
rect 15886 7306 15946 7382
rect 25957 7440 28231 7442
rect 25957 7384 25962 7440
rect 26018 7384 28170 7440
rect 28226 7384 28231 7440
rect 25957 7382 28231 7384
rect 25957 7379 26023 7382
rect 28165 7379 28231 7382
rect 34145 7442 34211 7445
rect 36537 7442 36603 7445
rect 34145 7440 36603 7442
rect 34145 7384 34150 7440
rect 34206 7384 36542 7440
rect 36598 7384 36603 7440
rect 34145 7382 36603 7384
rect 34145 7379 34211 7382
rect 36537 7379 36603 7382
rect 19793 7306 19859 7309
rect 24853 7306 24919 7309
rect 36261 7306 36327 7309
rect 37549 7306 37615 7309
rect 9949 7304 15762 7306
rect 9949 7248 9954 7304
rect 10010 7248 14738 7304
rect 14794 7248 15762 7304
rect 9949 7246 15762 7248
rect 15886 7304 24919 7306
rect 15886 7248 19798 7304
rect 19854 7248 24858 7304
rect 24914 7248 24919 7304
rect 15886 7246 24919 7248
rect 9949 7243 10015 7246
rect 14733 7243 14799 7246
rect 8385 7170 8451 7173
rect 8518 7170 8524 7172
rect 8385 7168 8524 7170
rect 8385 7112 8390 7168
rect 8446 7112 8524 7168
rect 8385 7110 8524 7112
rect 8385 7107 8451 7110
rect 8518 7108 8524 7110
rect 8588 7108 8594 7172
rect 9857 7170 9923 7173
rect 14089 7170 14155 7173
rect 9857 7168 14155 7170
rect 9857 7112 9862 7168
rect 9918 7112 14094 7168
rect 14150 7112 14155 7168
rect 9857 7110 14155 7112
rect 15702 7170 15762 7246
rect 19793 7243 19859 7246
rect 24853 7243 24919 7246
rect 26926 7304 37615 7306
rect 26926 7248 36266 7304
rect 36322 7248 37554 7304
rect 37610 7248 37615 7304
rect 26926 7246 37615 7248
rect 26926 7170 26986 7246
rect 36261 7243 36327 7246
rect 37549 7243 37615 7246
rect 15702 7110 26986 7170
rect 9857 7107 9923 7110
rect 14089 7107 14155 7110
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 6177 7034 6243 7037
rect 5950 7032 6243 7034
rect 5950 6976 6182 7032
rect 6238 6976 6243 7032
rect 5950 6974 6243 6976
rect 3785 6898 3851 6901
rect 5950 6898 6010 6974
rect 6177 6971 6243 6974
rect 3785 6896 6010 6898
rect 3785 6840 3790 6896
rect 3846 6840 6010 6896
rect 3785 6838 6010 6840
rect 6177 6898 6243 6901
rect 7465 6898 7531 6901
rect 6177 6896 7531 6898
rect 6177 6840 6182 6896
rect 6238 6840 7470 6896
rect 7526 6840 7531 6896
rect 6177 6838 7531 6840
rect 3785 6835 3851 6838
rect 6177 6835 6243 6838
rect 7465 6835 7531 6838
rect 8385 6898 8451 6901
rect 9581 6898 9647 6901
rect 22645 6898 22711 6901
rect 8385 6896 22711 6898
rect 8385 6840 8390 6896
rect 8446 6840 9586 6896
rect 9642 6840 22650 6896
rect 22706 6840 22711 6896
rect 8385 6838 22711 6840
rect 8385 6835 8451 6838
rect 9581 6835 9647 6838
rect 22645 6835 22711 6838
rect 22829 6898 22895 6901
rect 24945 6898 25011 6901
rect 22829 6896 25011 6898
rect 22829 6840 22834 6896
rect 22890 6840 24950 6896
rect 25006 6840 25011 6896
rect 22829 6838 25011 6840
rect 22829 6835 22895 6838
rect 24945 6835 25011 6838
rect 7005 6762 7071 6765
rect 9949 6762 10015 6765
rect 7005 6760 10015 6762
rect 7005 6704 7010 6760
rect 7066 6704 9954 6760
rect 10010 6704 10015 6760
rect 7005 6702 10015 6704
rect 7005 6699 7071 6702
rect 9949 6699 10015 6702
rect 10133 6762 10199 6765
rect 14825 6762 14891 6765
rect 10133 6760 14891 6762
rect 10133 6704 10138 6760
rect 10194 6704 14830 6760
rect 14886 6704 14891 6760
rect 10133 6702 14891 6704
rect 10133 6699 10199 6702
rect 14825 6699 14891 6702
rect 26877 6762 26943 6765
rect 26877 6760 35634 6762
rect 26877 6704 26882 6760
rect 26938 6704 35634 6760
rect 26877 6702 35634 6704
rect 26877 6699 26943 6702
rect 0 6626 480 6656
rect 5901 6626 5967 6629
rect 0 6624 5967 6626
rect 0 6568 5906 6624
rect 5962 6568 5967 6624
rect 0 6566 5967 6568
rect 0 6536 480 6566
rect 5901 6563 5967 6566
rect 8845 6626 8911 6629
rect 13353 6626 13419 6629
rect 16849 6626 16915 6629
rect 8845 6624 16915 6626
rect 8845 6568 8850 6624
rect 8906 6568 13358 6624
rect 13414 6568 16854 6624
rect 16910 6568 16915 6624
rect 8845 6566 16915 6568
rect 35574 6626 35634 6702
rect 39520 6626 40000 6656
rect 35574 6566 40000 6626
rect 8845 6563 8911 6566
rect 13353 6563 13419 6566
rect 16849 6563 16915 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6566
rect 34277 6495 34597 6496
rect 24945 6490 25011 6493
rect 30833 6490 30899 6493
rect 24945 6488 30899 6490
rect 24945 6432 24950 6488
rect 25006 6432 30838 6488
rect 30894 6432 30899 6488
rect 24945 6430 30899 6432
rect 24945 6427 25011 6430
rect 30833 6427 30899 6430
rect 11329 6354 11395 6357
rect 13813 6354 13879 6357
rect 20069 6354 20135 6357
rect 11329 6352 20135 6354
rect 11329 6296 11334 6352
rect 11390 6296 13818 6352
rect 13874 6296 20074 6352
rect 20130 6296 20135 6352
rect 11329 6294 20135 6296
rect 11329 6291 11395 6294
rect 13813 6291 13879 6294
rect 20069 6291 20135 6294
rect 21633 6354 21699 6357
rect 28993 6354 29059 6357
rect 32305 6354 32371 6357
rect 21633 6352 32371 6354
rect 21633 6296 21638 6352
rect 21694 6296 28998 6352
rect 29054 6296 32310 6352
rect 32366 6296 32371 6352
rect 21633 6294 32371 6296
rect 21633 6291 21699 6294
rect 28993 6291 29059 6294
rect 32305 6291 32371 6294
rect 6637 6218 6703 6221
rect 10133 6218 10199 6221
rect 6637 6216 10199 6218
rect 6637 6160 6642 6216
rect 6698 6160 10138 6216
rect 10194 6160 10199 6216
rect 6637 6158 10199 6160
rect 6637 6155 6703 6158
rect 10133 6155 10199 6158
rect 11237 6218 11303 6221
rect 21817 6218 21883 6221
rect 11237 6216 21883 6218
rect 11237 6160 11242 6216
rect 11298 6160 21822 6216
rect 21878 6160 21883 6216
rect 11237 6158 21883 6160
rect 11237 6155 11303 6158
rect 21817 6155 21883 6158
rect 24393 6218 24459 6221
rect 29545 6218 29611 6221
rect 24393 6216 29611 6218
rect 24393 6160 24398 6216
rect 24454 6160 29550 6216
rect 29606 6160 29611 6216
rect 24393 6158 29611 6160
rect 24393 6155 24459 6158
rect 29545 6155 29611 6158
rect 35249 6218 35315 6221
rect 36537 6218 36603 6221
rect 35249 6216 36603 6218
rect 35249 6160 35254 6216
rect 35310 6160 36542 6216
rect 36598 6160 36603 6216
rect 35249 6158 36603 6160
rect 35249 6155 35315 6158
rect 36537 6155 36603 6158
rect 15561 6082 15627 6085
rect 21633 6082 21699 6085
rect 15561 6080 21699 6082
rect 15561 6024 15566 6080
rect 15622 6024 21638 6080
rect 21694 6024 21699 6080
rect 15561 6022 21699 6024
rect 15561 6019 15627 6022
rect 21633 6019 21699 6022
rect 31201 6082 31267 6085
rect 33133 6082 33199 6085
rect 31201 6080 33199 6082
rect 31201 6024 31206 6080
rect 31262 6024 33138 6080
rect 33194 6024 33199 6080
rect 31201 6022 33199 6024
rect 31201 6019 31267 6022
rect 33133 6019 33199 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 3141 5946 3207 5949
rect 6269 5946 6335 5949
rect 3141 5944 6335 5946
rect 3141 5888 3146 5944
rect 3202 5888 6274 5944
rect 6330 5888 6335 5944
rect 3141 5886 6335 5888
rect 3141 5883 3207 5886
rect 6269 5883 6335 5886
rect 33041 5946 33107 5949
rect 35801 5946 35867 5949
rect 33041 5944 35867 5946
rect 33041 5888 33046 5944
rect 33102 5888 35806 5944
rect 35862 5888 35867 5944
rect 33041 5886 35867 5888
rect 33041 5883 33107 5886
rect 35801 5883 35867 5886
rect 0 5810 480 5840
rect 9029 5810 9095 5813
rect 0 5808 9095 5810
rect 0 5752 9034 5808
rect 9090 5752 9095 5808
rect 0 5750 9095 5752
rect 0 5720 480 5750
rect 9029 5747 9095 5750
rect 31201 5810 31267 5813
rect 35433 5810 35499 5813
rect 31201 5808 35499 5810
rect 31201 5752 31206 5808
rect 31262 5752 35438 5808
rect 35494 5752 35499 5808
rect 31201 5750 35499 5752
rect 31201 5747 31267 5750
rect 35433 5747 35499 5750
rect 37181 5810 37247 5813
rect 39520 5810 40000 5840
rect 37181 5808 40000 5810
rect 37181 5752 37186 5808
rect 37242 5752 40000 5808
rect 37181 5750 40000 5752
rect 37181 5747 37247 5750
rect 39520 5720 40000 5750
rect 10041 5674 10107 5677
rect 15653 5674 15719 5677
rect 19333 5674 19399 5677
rect 25313 5674 25379 5677
rect 27337 5674 27403 5677
rect 29269 5674 29335 5677
rect 10041 5672 19399 5674
rect 10041 5616 10046 5672
rect 10102 5616 15658 5672
rect 15714 5616 19338 5672
rect 19394 5616 19399 5672
rect 10041 5614 19399 5616
rect 10041 5611 10107 5614
rect 15653 5611 15719 5614
rect 19333 5611 19399 5614
rect 20670 5614 21466 5674
rect 2773 5538 2839 5541
rect 3325 5538 3391 5541
rect 2773 5536 3391 5538
rect 2773 5480 2778 5536
rect 2834 5480 3330 5536
rect 3386 5480 3391 5536
rect 2773 5478 3391 5480
rect 2773 5475 2839 5478
rect 3325 5475 3391 5478
rect 17033 5538 17099 5541
rect 20670 5538 20730 5614
rect 17033 5536 20730 5538
rect 17033 5480 17038 5536
rect 17094 5480 20730 5536
rect 17033 5478 20730 5480
rect 21406 5538 21466 5614
rect 25313 5672 29335 5674
rect 25313 5616 25318 5672
rect 25374 5616 27342 5672
rect 27398 5616 29274 5672
rect 29330 5616 29335 5672
rect 25313 5614 29335 5616
rect 25313 5611 25379 5614
rect 27337 5611 27403 5614
rect 29269 5611 29335 5614
rect 23105 5538 23171 5541
rect 21406 5536 23171 5538
rect 21406 5480 23110 5536
rect 23166 5480 23171 5536
rect 21406 5478 23171 5480
rect 17033 5475 17099 5478
rect 23105 5475 23171 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 1577 5402 1643 5405
rect 2957 5402 3023 5405
rect 1577 5400 3023 5402
rect 1577 5344 1582 5400
rect 1638 5344 2962 5400
rect 3018 5344 3023 5400
rect 1577 5342 3023 5344
rect 1577 5339 1643 5342
rect 2957 5339 3023 5342
rect 3969 5402 4035 5405
rect 5533 5402 5599 5405
rect 3969 5400 5599 5402
rect 3969 5344 3974 5400
rect 4030 5344 5538 5400
rect 5594 5344 5599 5400
rect 3969 5342 5599 5344
rect 3969 5339 4035 5342
rect 5533 5339 5599 5342
rect 9949 5266 10015 5269
rect 18229 5266 18295 5269
rect 9949 5264 18295 5266
rect 9949 5208 9954 5264
rect 10010 5208 18234 5264
rect 18290 5208 18295 5264
rect 9949 5206 18295 5208
rect 9949 5203 10015 5206
rect 18229 5203 18295 5206
rect 19057 5266 19123 5269
rect 22093 5266 22159 5269
rect 19057 5264 22159 5266
rect 19057 5208 19062 5264
rect 19118 5208 22098 5264
rect 22154 5208 22159 5264
rect 19057 5206 22159 5208
rect 19057 5203 19123 5206
rect 22093 5203 22159 5206
rect 26969 5266 27035 5269
rect 28441 5266 28507 5269
rect 26969 5264 28507 5266
rect 26969 5208 26974 5264
rect 27030 5208 28446 5264
rect 28502 5208 28507 5264
rect 26969 5206 28507 5208
rect 26969 5203 27035 5206
rect 28441 5203 28507 5206
rect 33317 5266 33383 5269
rect 37365 5266 37431 5269
rect 33317 5264 37431 5266
rect 33317 5208 33322 5264
rect 33378 5208 37370 5264
rect 37426 5208 37431 5264
rect 33317 5206 37431 5208
rect 33317 5203 33383 5206
rect 37365 5203 37431 5206
rect 10593 5130 10659 5133
rect 12525 5130 12591 5133
rect 10593 5128 12591 5130
rect 10593 5072 10598 5128
rect 10654 5072 12530 5128
rect 12586 5072 12591 5128
rect 10593 5070 12591 5072
rect 10593 5067 10659 5070
rect 12525 5067 12591 5070
rect 13077 5130 13143 5133
rect 14641 5130 14707 5133
rect 13077 5128 14707 5130
rect 13077 5072 13082 5128
rect 13138 5072 14646 5128
rect 14702 5072 14707 5128
rect 13077 5070 14707 5072
rect 13077 5067 13143 5070
rect 14641 5067 14707 5070
rect 15377 5130 15443 5133
rect 25405 5130 25471 5133
rect 15377 5128 25471 5130
rect 15377 5072 15382 5128
rect 15438 5072 25410 5128
rect 25466 5072 25471 5128
rect 15377 5070 25471 5072
rect 15377 5067 15443 5070
rect 25405 5067 25471 5070
rect 11697 4994 11763 4997
rect 13813 4994 13879 4997
rect 11697 4992 13879 4994
rect 11697 4936 11702 4992
rect 11758 4936 13818 4992
rect 13874 4936 13879 4992
rect 11697 4934 13879 4936
rect 11697 4931 11763 4934
rect 13813 4931 13879 4934
rect 16389 4994 16455 4997
rect 18045 4994 18111 4997
rect 16389 4992 18111 4994
rect 16389 4936 16394 4992
rect 16450 4936 18050 4992
rect 18106 4936 18111 4992
rect 16389 4934 18111 4936
rect 16389 4931 16455 4934
rect 18045 4931 18111 4934
rect 24577 4994 24643 4997
rect 26877 4994 26943 4997
rect 24577 4992 26943 4994
rect 24577 4936 24582 4992
rect 24638 4936 26882 4992
rect 26938 4936 26943 4992
rect 24577 4934 26943 4936
rect 24577 4931 24643 4934
rect 26877 4931 26943 4934
rect 14277 4928 14597 4929
rect 0 4858 480 4888
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 565 4858 631 4861
rect 0 4856 631 4858
rect 0 4800 570 4856
rect 626 4800 631 4856
rect 0 4798 631 4800
rect 0 4768 480 4798
rect 565 4795 631 4798
rect 4153 4858 4219 4861
rect 9765 4858 9831 4861
rect 4153 4856 9831 4858
rect 4153 4800 4158 4856
rect 4214 4800 9770 4856
rect 9826 4800 9831 4856
rect 4153 4798 9831 4800
rect 4153 4795 4219 4798
rect 9765 4795 9831 4798
rect 17769 4858 17835 4861
rect 21265 4858 21331 4861
rect 17769 4856 21331 4858
rect 17769 4800 17774 4856
rect 17830 4800 21270 4856
rect 21326 4800 21331 4856
rect 17769 4798 21331 4800
rect 17769 4795 17835 4798
rect 21265 4795 21331 4798
rect 35525 4858 35591 4861
rect 39520 4858 40000 4888
rect 35525 4856 40000 4858
rect 35525 4800 35530 4856
rect 35586 4800 40000 4856
rect 35525 4798 40000 4800
rect 35525 4795 35591 4798
rect 39520 4768 40000 4798
rect 7833 4722 7899 4725
rect 9673 4722 9739 4725
rect 7833 4720 9739 4722
rect 7833 4664 7838 4720
rect 7894 4664 9678 4720
rect 9734 4664 9739 4720
rect 7833 4662 9739 4664
rect 7833 4659 7899 4662
rect 9673 4659 9739 4662
rect 11513 4722 11579 4725
rect 19885 4722 19951 4725
rect 11513 4720 19951 4722
rect 11513 4664 11518 4720
rect 11574 4664 19890 4720
rect 19946 4664 19951 4720
rect 11513 4662 19951 4664
rect 11513 4659 11579 4662
rect 19885 4659 19951 4662
rect 23105 4722 23171 4725
rect 23565 4722 23631 4725
rect 30373 4722 30439 4725
rect 23105 4720 30439 4722
rect 23105 4664 23110 4720
rect 23166 4664 23570 4720
rect 23626 4664 30378 4720
rect 30434 4664 30439 4720
rect 23105 4662 30439 4664
rect 23105 4659 23171 4662
rect 23565 4659 23631 4662
rect 30373 4659 30439 4662
rect 4797 4586 4863 4589
rect 8201 4586 8267 4589
rect 4797 4584 8267 4586
rect 4797 4528 4802 4584
rect 4858 4528 8206 4584
rect 8262 4528 8267 4584
rect 4797 4526 8267 4528
rect 4797 4523 4863 4526
rect 8201 4523 8267 4526
rect 11881 4586 11947 4589
rect 14733 4586 14799 4589
rect 11881 4584 14799 4586
rect 11881 4528 11886 4584
rect 11942 4528 14738 4584
rect 14794 4528 14799 4584
rect 11881 4526 14799 4528
rect 11881 4523 11947 4526
rect 14733 4523 14799 4526
rect 15745 4586 15811 4589
rect 32581 4586 32647 4589
rect 15745 4584 32647 4586
rect 15745 4528 15750 4584
rect 15806 4528 32586 4584
rect 32642 4528 32647 4584
rect 15745 4526 32647 4528
rect 15745 4523 15811 4526
rect 32581 4523 32647 4526
rect 3049 4450 3115 4453
rect 5717 4450 5783 4453
rect 3049 4448 5783 4450
rect 3049 4392 3054 4448
rect 3110 4392 5722 4448
rect 5778 4392 5783 4448
rect 3049 4390 5783 4392
rect 3049 4387 3115 4390
rect 5717 4387 5783 4390
rect 26785 4450 26851 4453
rect 30557 4450 30623 4453
rect 26785 4448 30623 4450
rect 26785 4392 26790 4448
rect 26846 4392 30562 4448
rect 30618 4392 30623 4448
rect 26785 4390 30623 4392
rect 26785 4387 26851 4390
rect 30557 4387 30623 4390
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 28809 4314 28875 4317
rect 28809 4312 34162 4314
rect 28809 4256 28814 4312
rect 28870 4256 34162 4312
rect 28809 4254 34162 4256
rect 28809 4251 28875 4254
rect 4705 4178 4771 4181
rect 9029 4178 9095 4181
rect 9765 4178 9831 4181
rect 4705 4176 9831 4178
rect 4705 4120 4710 4176
rect 4766 4120 9034 4176
rect 9090 4120 9770 4176
rect 9826 4120 9831 4176
rect 4705 4118 9831 4120
rect 4705 4115 4771 4118
rect 9029 4115 9095 4118
rect 9765 4115 9831 4118
rect 11145 4178 11211 4181
rect 18045 4178 18111 4181
rect 11145 4176 18111 4178
rect 11145 4120 11150 4176
rect 11206 4120 18050 4176
rect 18106 4120 18111 4176
rect 11145 4118 18111 4120
rect 11145 4115 11211 4118
rect 18045 4115 18111 4118
rect 29729 4178 29795 4181
rect 32121 4178 32187 4181
rect 29729 4176 32187 4178
rect 29729 4120 29734 4176
rect 29790 4120 32126 4176
rect 32182 4120 32187 4176
rect 29729 4118 32187 4120
rect 34102 4178 34162 4254
rect 36353 4178 36419 4181
rect 34102 4176 36419 4178
rect 34102 4120 36358 4176
rect 36414 4120 36419 4176
rect 34102 4118 36419 4120
rect 29729 4115 29795 4118
rect 32121 4115 32187 4118
rect 36353 4115 36419 4118
rect 0 4042 480 4072
rect 2497 4042 2563 4045
rect 3509 4042 3575 4045
rect 0 3982 1410 4042
rect 0 3952 480 3982
rect 1350 3906 1410 3982
rect 2497 4040 3575 4042
rect 2497 3984 2502 4040
rect 2558 3984 3514 4040
rect 3570 3984 3575 4040
rect 2497 3982 3575 3984
rect 2497 3979 2563 3982
rect 3509 3979 3575 3982
rect 4245 4042 4311 4045
rect 6913 4042 6979 4045
rect 4245 4040 6979 4042
rect 4245 3984 4250 4040
rect 4306 3984 6918 4040
rect 6974 3984 6979 4040
rect 4245 3982 6979 3984
rect 4245 3979 4311 3982
rect 6913 3979 6979 3982
rect 9581 4042 9647 4045
rect 11237 4042 11303 4045
rect 9581 4040 11303 4042
rect 9581 3984 9586 4040
rect 9642 3984 11242 4040
rect 11298 3984 11303 4040
rect 9581 3982 11303 3984
rect 9581 3979 9647 3982
rect 11237 3979 11303 3982
rect 12985 4042 13051 4045
rect 16941 4042 17007 4045
rect 12985 4040 17007 4042
rect 12985 3984 12990 4040
rect 13046 3984 16946 4040
rect 17002 3984 17007 4040
rect 12985 3982 17007 3984
rect 12985 3979 13051 3982
rect 16941 3979 17007 3982
rect 18781 4042 18847 4045
rect 28073 4042 28139 4045
rect 31569 4042 31635 4045
rect 35249 4042 35315 4045
rect 18781 4040 27538 4042
rect 18781 3984 18786 4040
rect 18842 3984 27538 4040
rect 18781 3982 27538 3984
rect 18781 3979 18847 3982
rect 3785 3906 3851 3909
rect 1350 3904 3851 3906
rect 1350 3848 3790 3904
rect 3846 3848 3851 3904
rect 1350 3846 3851 3848
rect 3785 3843 3851 3846
rect 5533 3906 5599 3909
rect 10225 3906 10291 3909
rect 5533 3904 10291 3906
rect 5533 3848 5538 3904
rect 5594 3848 10230 3904
rect 10286 3848 10291 3904
rect 5533 3846 10291 3848
rect 5533 3843 5599 3846
rect 10225 3843 10291 3846
rect 24669 3906 24735 3909
rect 26325 3906 26391 3909
rect 24669 3904 26391 3906
rect 24669 3848 24674 3904
rect 24730 3848 26330 3904
rect 26386 3848 26391 3904
rect 24669 3846 26391 3848
rect 24669 3843 24735 3846
rect 26325 3843 26391 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 1117 3772 1183 3773
rect 1117 3770 1164 3772
rect 1072 3768 1164 3770
rect 1072 3712 1122 3768
rect 1072 3710 1164 3712
rect 1117 3708 1164 3710
rect 1228 3708 1234 3772
rect 7373 3770 7439 3773
rect 13077 3770 13143 3773
rect 7373 3768 13143 3770
rect 7373 3712 7378 3768
rect 7434 3712 13082 3768
rect 13138 3712 13143 3768
rect 7373 3710 13143 3712
rect 1117 3707 1183 3708
rect 7373 3707 7439 3710
rect 13077 3707 13143 3710
rect 17861 3770 17927 3773
rect 24117 3770 24183 3773
rect 17861 3768 24183 3770
rect 17861 3712 17866 3768
rect 17922 3712 24122 3768
rect 24178 3712 24183 3768
rect 17861 3710 24183 3712
rect 17861 3707 17927 3710
rect 24117 3707 24183 3710
rect 5349 3634 5415 3637
rect 12157 3634 12223 3637
rect 5349 3632 12223 3634
rect 5349 3576 5354 3632
rect 5410 3576 12162 3632
rect 12218 3576 12223 3632
rect 5349 3574 12223 3576
rect 5349 3571 5415 3574
rect 12157 3571 12223 3574
rect 13537 3634 13603 3637
rect 15469 3634 15535 3637
rect 19057 3634 19123 3637
rect 13537 3632 19123 3634
rect 13537 3576 13542 3632
rect 13598 3576 15474 3632
rect 15530 3576 19062 3632
rect 19118 3576 19123 3632
rect 13537 3574 19123 3576
rect 27478 3634 27538 3982
rect 28073 4040 35315 4042
rect 28073 3984 28078 4040
rect 28134 3984 31574 4040
rect 31630 3984 35254 4040
rect 35310 3984 35315 4040
rect 28073 3982 35315 3984
rect 28073 3979 28139 3982
rect 31569 3979 31635 3982
rect 35249 3979 35315 3982
rect 38009 4042 38075 4045
rect 39520 4042 40000 4072
rect 38009 4040 40000 4042
rect 38009 3984 38014 4040
rect 38070 3984 40000 4040
rect 38009 3982 40000 3984
rect 38009 3979 38075 3982
rect 39520 3952 40000 3982
rect 28349 3906 28415 3909
rect 36445 3906 36511 3909
rect 28349 3904 36511 3906
rect 28349 3848 28354 3904
rect 28410 3848 36450 3904
rect 36506 3848 36511 3904
rect 28349 3846 36511 3848
rect 28349 3843 28415 3846
rect 36445 3843 36511 3846
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 30189 3634 30255 3637
rect 27478 3632 30255 3634
rect 27478 3576 30194 3632
rect 30250 3576 30255 3632
rect 27478 3574 30255 3576
rect 13537 3571 13603 3574
rect 15469 3571 15535 3574
rect 19057 3571 19123 3574
rect 30189 3571 30255 3574
rect 8753 3498 8819 3501
rect 10501 3498 10567 3501
rect 8753 3496 10567 3498
rect 8753 3440 8758 3496
rect 8814 3440 10506 3496
rect 10562 3440 10567 3496
rect 8753 3438 10567 3440
rect 8753 3435 8819 3438
rect 10501 3435 10567 3438
rect 12801 3498 12867 3501
rect 14917 3498 14983 3501
rect 12801 3496 14983 3498
rect 12801 3440 12806 3496
rect 12862 3440 14922 3496
rect 14978 3440 14983 3496
rect 12801 3438 14983 3440
rect 12801 3435 12867 3438
rect 14917 3435 14983 3438
rect 24025 3498 24091 3501
rect 30833 3498 30899 3501
rect 24025 3496 30899 3498
rect 24025 3440 24030 3496
rect 24086 3440 30838 3496
rect 30894 3440 30899 3496
rect 24025 3438 30899 3440
rect 24025 3435 24091 3438
rect 30833 3435 30899 3438
rect 12617 3362 12683 3365
rect 15745 3362 15811 3365
rect 12617 3360 15811 3362
rect 12617 3304 12622 3360
rect 12678 3304 15750 3360
rect 15806 3304 15811 3360
rect 12617 3302 15811 3304
rect 12617 3299 12683 3302
rect 15745 3299 15811 3302
rect 22737 3362 22803 3365
rect 25497 3362 25563 3365
rect 22737 3360 25563 3362
rect 22737 3304 22742 3360
rect 22798 3304 25502 3360
rect 25558 3304 25563 3360
rect 22737 3302 25563 3304
rect 22737 3299 22803 3302
rect 25497 3299 25563 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 34973 3226 35039 3229
rect 37273 3226 37339 3229
rect 34973 3224 37339 3226
rect 34973 3168 34978 3224
rect 35034 3168 37278 3224
rect 37334 3168 37339 3224
rect 34973 3166 37339 3168
rect 34973 3163 35039 3166
rect 37273 3163 37339 3166
rect 0 3090 480 3120
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 0 3000 480 3030
rect 3417 3027 3483 3030
rect 6085 3090 6151 3093
rect 6085 3088 7114 3090
rect 6085 3032 6090 3088
rect 6146 3032 7114 3088
rect 6085 3030 7114 3032
rect 6085 3027 6151 3030
rect 1669 2954 1735 2957
rect 6913 2954 6979 2957
rect 1669 2952 6979 2954
rect 1669 2896 1674 2952
rect 1730 2896 6918 2952
rect 6974 2896 6979 2952
rect 1669 2894 6979 2896
rect 7054 2954 7114 3030
rect 15142 3028 15148 3092
rect 15212 3090 15218 3092
rect 16021 3090 16087 3093
rect 15212 3088 16087 3090
rect 15212 3032 16026 3088
rect 16082 3032 16087 3088
rect 15212 3030 16087 3032
rect 15212 3028 15218 3030
rect 16021 3027 16087 3030
rect 16573 3090 16639 3093
rect 21265 3090 21331 3093
rect 16573 3088 21331 3090
rect 16573 3032 16578 3088
rect 16634 3032 21270 3088
rect 21326 3032 21331 3088
rect 16573 3030 21331 3032
rect 16573 3027 16639 3030
rect 21265 3027 21331 3030
rect 22001 3090 22067 3093
rect 39389 3090 39455 3093
rect 39520 3090 40000 3120
rect 22001 3088 22202 3090
rect 22001 3032 22006 3088
rect 22062 3032 22202 3088
rect 22001 3030 22202 3032
rect 22001 3027 22067 3030
rect 8109 2954 8175 2957
rect 12525 2954 12591 2957
rect 7054 2952 12591 2954
rect 7054 2896 8114 2952
rect 8170 2896 12530 2952
rect 12586 2896 12591 2952
rect 7054 2894 12591 2896
rect 1669 2891 1735 2894
rect 6913 2891 6979 2894
rect 8109 2891 8175 2894
rect 12525 2891 12591 2894
rect 14089 2954 14155 2957
rect 18321 2954 18387 2957
rect 14089 2952 18387 2954
rect 14089 2896 14094 2952
rect 14150 2896 18326 2952
rect 18382 2896 18387 2952
rect 14089 2894 18387 2896
rect 22142 2954 22202 3030
rect 39389 3088 40000 3090
rect 39389 3032 39394 3088
rect 39450 3032 40000 3088
rect 39389 3030 40000 3032
rect 39389 3027 39455 3030
rect 39520 3000 40000 3030
rect 39389 2954 39455 2957
rect 22142 2952 39455 2954
rect 22142 2896 39394 2952
rect 39450 2896 39455 2952
rect 22142 2894 39455 2896
rect 14089 2891 14155 2894
rect 18321 2891 18387 2894
rect 39389 2891 39455 2894
rect 5901 2818 5967 2821
rect 9489 2818 9555 2821
rect 5901 2816 9555 2818
rect 5901 2760 5906 2816
rect 5962 2760 9494 2816
rect 9550 2760 9555 2816
rect 5901 2758 9555 2760
rect 5901 2755 5967 2758
rect 9489 2755 9555 2758
rect 29453 2818 29519 2821
rect 29821 2818 29887 2821
rect 29453 2816 29887 2818
rect 29453 2760 29458 2816
rect 29514 2760 29826 2816
rect 29882 2760 29887 2816
rect 29453 2758 29887 2760
rect 29453 2755 29519 2758
rect 29821 2755 29887 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 9397 2682 9463 2685
rect 13261 2682 13327 2685
rect 9397 2680 13327 2682
rect 9397 2624 9402 2680
rect 9458 2624 13266 2680
rect 13322 2624 13327 2680
rect 9397 2622 13327 2624
rect 9397 2619 9463 2622
rect 13261 2619 13327 2622
rect 17033 2682 17099 2685
rect 20897 2682 20963 2685
rect 38745 2682 38811 2685
rect 17033 2680 20963 2682
rect 17033 2624 17038 2680
rect 17094 2624 20902 2680
rect 20958 2624 20963 2680
rect 17033 2622 20963 2624
rect 17033 2619 17099 2622
rect 20897 2619 20963 2622
rect 34654 2680 38811 2682
rect 34654 2624 38750 2680
rect 38806 2624 38811 2680
rect 34654 2622 38811 2624
rect 6913 2546 6979 2549
rect 13905 2546 13971 2549
rect 6913 2544 13971 2546
rect 6913 2488 6918 2544
rect 6974 2488 13910 2544
rect 13966 2488 13971 2544
rect 6913 2486 13971 2488
rect 6913 2483 6979 2486
rect 13905 2483 13971 2486
rect 15561 2546 15627 2549
rect 18321 2546 18387 2549
rect 15561 2544 18387 2546
rect 15561 2488 15566 2544
rect 15622 2488 18326 2544
rect 18382 2488 18387 2544
rect 15561 2486 18387 2488
rect 15561 2483 15627 2486
rect 18321 2483 18387 2486
rect 20621 2546 20687 2549
rect 21817 2546 21883 2549
rect 22645 2546 22711 2549
rect 26693 2546 26759 2549
rect 20621 2544 26759 2546
rect 20621 2488 20626 2544
rect 20682 2488 21822 2544
rect 21878 2488 22650 2544
rect 22706 2488 26698 2544
rect 26754 2488 26759 2544
rect 20621 2486 26759 2488
rect 20621 2483 20687 2486
rect 21817 2483 21883 2486
rect 22645 2483 22711 2486
rect 26693 2483 26759 2486
rect 27705 2546 27771 2549
rect 29545 2546 29611 2549
rect 27705 2544 29611 2546
rect 27705 2488 27710 2544
rect 27766 2488 29550 2544
rect 29606 2488 29611 2544
rect 27705 2486 29611 2488
rect 27705 2483 27771 2486
rect 29545 2483 29611 2486
rect 11881 2410 11947 2413
rect 34654 2410 34714 2622
rect 38745 2619 38811 2622
rect 35893 2410 35959 2413
rect 11881 2408 34714 2410
rect 11881 2352 11886 2408
rect 11942 2352 34714 2408
rect 11881 2350 34714 2352
rect 34838 2408 35959 2410
rect 34838 2352 35898 2408
rect 35954 2352 35959 2408
rect 34838 2350 35959 2352
rect 11881 2347 11947 2350
rect 0 2274 480 2304
rect 4889 2274 4955 2277
rect 0 2272 4955 2274
rect 0 2216 4894 2272
rect 4950 2216 4955 2272
rect 0 2214 4955 2216
rect 0 2184 480 2214
rect 4889 2211 4955 2214
rect 12893 2274 12959 2277
rect 20069 2274 20135 2277
rect 12893 2272 20135 2274
rect 12893 2216 12898 2272
rect 12954 2216 20074 2272
rect 20130 2216 20135 2272
rect 12893 2214 20135 2216
rect 12893 2211 12959 2214
rect 20069 2211 20135 2214
rect 25957 2274 26023 2277
rect 34053 2274 34119 2277
rect 25957 2272 34119 2274
rect 25957 2216 25962 2272
rect 26018 2216 34058 2272
rect 34114 2216 34119 2272
rect 25957 2214 34119 2216
rect 25957 2211 26023 2214
rect 34053 2211 34119 2214
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 27061 2138 27127 2141
rect 33133 2138 33199 2141
rect 27061 2136 33199 2138
rect 27061 2080 27066 2136
rect 27122 2080 33138 2136
rect 33194 2080 33199 2136
rect 27061 2078 33199 2080
rect 27061 2075 27127 2078
rect 33133 2075 33199 2078
rect 5257 2002 5323 2005
rect 14825 2002 14891 2005
rect 5257 2000 14891 2002
rect 5257 1944 5262 2000
rect 5318 1944 14830 2000
rect 14886 1944 14891 2000
rect 5257 1942 14891 1944
rect 5257 1939 5323 1942
rect 14825 1939 14891 1942
rect 26969 2002 27035 2005
rect 34838 2002 34898 2350
rect 35893 2347 35959 2350
rect 39520 2274 40000 2304
rect 26969 2000 34898 2002
rect 26969 1944 26974 2000
rect 27030 1944 34898 2000
rect 26969 1942 34898 1944
rect 35574 2214 40000 2274
rect 26969 1939 27035 1942
rect 27429 1458 27495 1461
rect 35574 1458 35634 2214
rect 39520 2184 40000 2214
rect 27429 1456 35634 1458
rect 27429 1400 27434 1456
rect 27490 1400 35634 1456
rect 27429 1398 35634 1400
rect 27429 1395 27495 1398
rect 0 1322 480 1352
rect 7005 1322 7071 1325
rect 0 1320 7071 1322
rect 0 1264 7010 1320
rect 7066 1264 7071 1320
rect 0 1262 7071 1264
rect 0 1232 480 1262
rect 7005 1259 7071 1262
rect 35341 1322 35407 1325
rect 39520 1322 40000 1352
rect 35341 1320 40000 1322
rect 35341 1264 35346 1320
rect 35402 1264 40000 1320
rect 35341 1262 40000 1264
rect 35341 1259 35407 1262
rect 39520 1232 40000 1262
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
rect 36077 506 36143 509
rect 39520 506 40000 536
rect 36077 504 40000 506
rect 36077 448 36082 504
rect 36138 448 40000 504
rect 36077 446 40000 448
rect 36077 443 36143 446
rect 39520 416 40000 446
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 12204 11520 12268 11524
rect 12204 11464 12218 11520
rect 12218 11464 12268 11520
rect 12204 11460 12268 11464
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 11284 11248 11348 11252
rect 11284 11192 11298 11248
rect 11298 11192 11348 11248
rect 11284 11188 11348 11192
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 28212 10568 28276 10572
rect 28212 10512 28226 10568
rect 28226 10512 28276 10568
rect 28212 10508 28276 10512
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 11652 9888 11716 9892
rect 11652 9832 11702 9888
rect 11702 9832 11716 9888
rect 11652 9828 11716 9832
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 28212 9208 28276 9212
rect 28212 9152 28262 9208
rect 28262 9152 28276 9208
rect 28212 9148 28276 9152
rect 28948 9148 29012 9212
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 28948 8876 29012 8940
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 8524 7108 8588 7172
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 1164 3768 1228 3772
rect 1164 3712 1178 3768
rect 1178 3712 1228 3768
rect 1164 3708 1228 3712
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 15148 3028 15212 3092
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 12203 11524 12269 11525
rect 12203 11460 12204 11524
rect 12268 11460 12269 11524
rect 12203 11459 12269 11460
rect 11283 11252 11349 11253
rect 11283 11188 11284 11252
rect 11348 11188 11349 11252
rect 11283 11187 11349 11188
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 11286 9298 11346 11187
rect 12206 10658 12266 11459
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 11651 9892 11717 9893
rect 11651 9828 11652 9892
rect 11716 9828 11717 9892
rect 11651 9827 11717 9828
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 8523 7172 8589 7173
rect 8523 7108 8524 7172
rect 8588 7108 8589 7172
rect 8523 7107 8589 7108
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 8526 3178 8586 7107
rect 11654 3858 11714 9827
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 2752 14597 3776
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 28947 9212 29013 9213
rect 28947 9148 28948 9212
rect 29012 9148 29013 9212
rect 28947 9147 29013 9148
rect 28950 8941 29010 9147
rect 28947 8940 29013 8941
rect 28947 8876 28948 8940
rect 29012 8876 29013 8940
rect 28947 8875 29013 8876
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
<< via4 >>
rect 12118 10422 12354 10658
rect 11198 9062 11434 9298
rect 1078 3772 1314 3858
rect 1078 3708 1164 3772
rect 1164 3708 1228 3772
rect 1228 3708 1314 3772
rect 1078 3622 1314 3708
rect 11566 3622 11802 3858
rect 8438 2942 8674 3178
rect 15062 3092 15298 3178
rect 15062 3028 15148 3092
rect 15148 3028 15212 3092
rect 15212 3028 15298 3092
rect 15062 2942 15298 3028
rect 28126 10572 28362 10658
rect 28126 10508 28212 10572
rect 28212 10508 28276 10572
rect 28276 10508 28362 10572
rect 28126 10422 28362 10508
rect 28126 9212 28362 9298
rect 28126 9148 28212 9212
rect 28212 9148 28276 9212
rect 28276 9148 28362 9212
rect 28126 9062 28362 9148
<< metal5 >>
rect 12076 10658 28404 10700
rect 12076 10422 12118 10658
rect 12354 10422 28126 10658
rect 28362 10422 28404 10658
rect 12076 10380 28404 10422
rect 11156 9298 28404 9340
rect 11156 9062 11198 9298
rect 11434 9062 28126 9298
rect 28362 9062 28404 9298
rect 11156 9020 28404 9062
rect 1036 3858 11844 3900
rect 1036 3622 1078 3858
rect 1314 3622 11566 3858
rect 11802 3622 11844 3858
rect 1036 3580 11844 3622
rect 8396 3178 15340 3220
rect 8396 2942 8438 3178
rect 8674 2942 15062 3178
rect 15298 2942 15340 3178
rect 8396 2900 15340 2942
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_7
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_20
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_24 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_20
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_24
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _093_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__C
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_or3_4  _092_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _079_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_50
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_66 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _162_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_100
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_or3_4  _089_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_or4_4  _167_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use scs8hd_buf_1  _095_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__D
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_177
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _097_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _112_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _140_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_229
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_conb_1  _188_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23736 0 1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_272
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 27416 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_285
timestamp 1586364061
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_289
timestamp 1586364061
transform 1 0 27692 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_295
timestamp 1586364061
transform 1 0 28244 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27968 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_299
timestamp 1586364061
transform 1 0 28612 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28704 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_315
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 30636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_320
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_325
timestamp 1586364061
transform 1 0 31004 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_331
timestamp 1586364061
transform 1 0 31556 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_319
timestamp 1586364061
transform 1 0 30452 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_332
timestamp 1586364061
transform 1 0 31648 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_336
timestamp 1586364061
transform 1 0 32016 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_339
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 31832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 32200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_345
timestamp 1586364061
transform 1 0 32844 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 32384 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_349
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_349
timestamp 1586364061
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 33028 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_353
timestamp 1586364061
transform 1 0 33580 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33580 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_356
timestamp 1586364061
transform 1 0 33856 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_356
timestamp 1586364061
transform 1 0 33856 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34040 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_360
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_360
timestamp 1586364061
transform 1 0 34224 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_369
timestamp 1586364061
transform 1 0 35052 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_380
timestamp 1586364061
transform 1 0 36064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_376
timestamp 1586364061
transform 1 0 35696 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_380
timestamp 1586364061
transform 1 0 36064 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_376
timestamp 1586364061
transform 1 0 35696 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_387
timestamp 1586364061
transform 1 0 36708 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 36432 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_387 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36708 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_391 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 37076 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_398
timestamp 1586364061
transform 1 0 37720 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_402
timestamp 1586364061
transform 1 0 38088 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_406
timestamp 1586364061
transform 1 0 38456 0 1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_16
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_20
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_28
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_58
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _080_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 406 592
use scs8hd_nor3_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_103
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _076_
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_136
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _155_
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__D
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_188
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _147_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_222
timestamp 1586364061
transform 1 0 21528 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_226
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_242
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_259
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25484 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26588 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_6  FILLER_2_286
timestamp 1586364061
transform 1 0 27416 0 -1 3808
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28152 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 30176 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 29348 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_305
timestamp 1586364061
transform 1 0 29164 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_309
timestamp 1586364061
transform 1 0 29532 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_313
timestamp 1586364061
transform 1 0 29900 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_327
timestamp 1586364061
transform 1 0 31188 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_331
timestamp 1586364061
transform 1 0 31556 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_335
timestamp 1586364061
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_2_346
timestamp 1586364061
transform 1 0 32936 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35144 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_365
timestamp 1586364061
transform 1 0 34684 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_369
timestamp 1586364061
transform 1 0 35052 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_372
timestamp 1586364061
transform 1 0 35328 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_382
timestamp 1586364061
transform 1 0 36248 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_394
timestamp 1586364061
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_8
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_25
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_65
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _164_
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_128
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _138_
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_145
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 314 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_or4_4  _122_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 406 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_248
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_252
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_255
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26680 0 1 3808
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_3_289
timestamp 1586364061
transform 1 0 27692 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_295
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_299
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 29348 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_316
timestamp 1586364061
transform 1 0 30176 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31004 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_321
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 32384 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_334
timestamp 1586364061
transform 1 0 31832 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_351
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_355
timestamp 1586364061
transform 1 0 33764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_363
timestamp 1586364061
transform 1 0 34500 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  _206_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36432 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_376
timestamp 1586364061
transform 1 0 35696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_380
timestamp 1586364061
transform 1 0 36064 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 36984 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_388
timestamp 1586364061
transform 1 0 36800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_392
timestamp 1586364061
transform 1 0 37168 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_399
timestamp 1586364061
transform 1 0 37812 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_52
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 130 592
use scs8hd_nand2_4  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__122__C
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_240
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_250
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_254
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_267
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_302
timestamp 1586364061
transform 1 0 28888 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_308
timestamp 1586364061
transform 1 0 29440 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_316
timestamp 1586364061
transform 1 0 30176 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 30452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_328
timestamp 1586364061
transform 1 0 31280 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_332
timestamp 1586364061
transform 1 0 31648 0 -1 4896
box -38 -48 406 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 32568 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_340
timestamp 1586364061
transform 1 0 32384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_344
timestamp 1586364061
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33396 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_348
timestamp 1586364061
transform 1 0 33120 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35144 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_362
timestamp 1586364061
transform 1 0 34408 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_366
timestamp 1586364061
transform 1 0 34776 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_369
timestamp 1586364061
transform 1 0 35052 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_381
timestamp 1586364061
transform 1 0 36156 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_386
timestamp 1586364061
transform 1 0 36616 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_394
timestamp 1586364061
transform 1 0 37352 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_28
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_45
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _074_
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_103
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_256
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_260
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 406 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_267
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_272
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_289
timestamp 1586364061
transform 1 0 27692 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_299
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 31280 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_326
timestamp 1586364061
transform 1 0 31096 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 31740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_335
timestamp 1586364061
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 33856 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_350
timestamp 1586364061
transform 1 0 33304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_358
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_362
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_376
timestamp 1586364061
transform 1 0 35696 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_380
timestamp 1586364061
transform 1 0 36064 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_63
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_85
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_109
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_124
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _166_
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 15364 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_177
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_185
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_207
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_238
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_264
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_273
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_285
timestamp 1586364061
transform 1 0 27324 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_277
timestamp 1586364061
transform 1 0 26588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_290
timestamp 1586364061
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_302
timestamp 1586364061
transform 1 0 28888 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_294
timestamp 1586364061
transform 1 0 28152 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_298
timestamp 1586364061
transform 1 0 28520 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_302
timestamp 1586364061
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_308
timestamp 1586364061
transform 1 0 29440 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29624 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 29256 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_315
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_316
timestamp 1586364061
transform 1 0 30176 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 30268 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 31096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 30912 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_328
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_319
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_323
timestamp 1586364061
transform 1 0 30820 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 32476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_335
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_339
timestamp 1586364061
transform 1 0 32292 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_343
timestamp 1586364061
transform 1 0 32660 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33856 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_348
timestamp 1586364061
transform 1 0 33120 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35052 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_367
timestamp 1586364061
transform 1 0 34868 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_371
timestamp 1586364061
transform 1 0 35236 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36616 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_384
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_380
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_388
timestamp 1586364061
transform 1 0 36800 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_396
timestamp 1586364061
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_393
timestamp 1586364061
transform 1 0 37260 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_405
timestamp 1586364061
transform 1 0 38364 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_47
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_96
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_100
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use scs8hd_or2_4  _114_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 21804 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_222
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_268
timestamp 1586364061
transform 1 0 25760 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 27784 0 -1 7072
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26772 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_282
timestamp 1586364061
transform 1 0 27048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_286
timestamp 1586364061
transform 1 0 27416 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_301
timestamp 1586364061
transform 1 0 28796 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_305
timestamp 1586364061
transform 1 0 29164 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_308
timestamp 1586364061
transform 1 0 29440 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 31096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 30728 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_320
timestamp 1586364061
transform 1 0 30544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_332
timestamp 1586364061
transform 1 0 31648 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 33764 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_346
timestamp 1586364061
transform 1 0 32936 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_351
timestamp 1586364061
transform 1 0 33396 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34960 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35328 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_366
timestamp 1586364061
transform 1 0 34776 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_370
timestamp 1586364061
transform 1 0 35144 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35512 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36708 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_389
timestamp 1586364061
transform 1 0 36892 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_8
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _165_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_195
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_237
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_264
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_268
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27784 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_282
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_286
timestamp 1586364061
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 30268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_315
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 30820 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 30636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_319
timestamp 1586364061
transform 1 0 30452 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_332
timestamp 1586364061
transform 1 0 31648 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_336
timestamp 1586364061
transform 1 0 32016 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_339
timestamp 1586364061
transform 1 0 32292 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_343
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 36248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_393
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_118
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_287
timestamp 1586364061
transform 1 0 27508 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28428 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_291
timestamp 1586364061
transform 1 0 27876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_295
timestamp 1586364061
transform 1 0 28244 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_306
timestamp 1586364061
transform 1 0 29256 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_310
timestamp 1586364061
transform 1 0 29624 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_318
timestamp 1586364061
transform 1 0 30360 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_328
timestamp 1586364061
transform 1 0 31280 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33856 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_348
timestamp 1586364061
transform 1 0 33120 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_352
timestamp 1586364061
transform 1 0 33488 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_359
timestamp 1586364061
transform 1 0 34132 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_363
timestamp 1586364061
transform 1 0 34500 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_376
timestamp 1586364061
transform 1 0 35696 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_380
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_388
timestamp 1586364061
transform 1 0 36800 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_396
timestamp 1586364061
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_76
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_212
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 24288 0 1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_280
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_286
timestamp 1586364061
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_315
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 31188 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_320
timestamp 1586364061
transform 1 0 30544 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_324
timestamp 1586364061
transform 1 0 30912 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 32384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_338
timestamp 1586364061
transform 1 0 32200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  FILLER_11_346
timestamp 1586364061
transform 1 0 32936 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_388
timestamp 1586364061
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_392
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_399
timestamp 1586364061
transform 1 0 37812 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_123
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_231
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_12_249
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_255
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_6  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28796 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_293
timestamp 1586364061
transform 1 0 28060 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_297
timestamp 1586364061
transform 1 0 28428 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30360 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_310
timestamp 1586364061
transform 1 0 29624 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_321
timestamp 1586364061
transform 1 0 30636 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_12_329
timestamp 1586364061
transform 1 0 31372 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_335
timestamp 1586364061
transform 1 0 31924 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33580 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_346
timestamp 1586364061
transform 1 0 32936 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_351
timestamp 1586364061
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_355
timestamp 1586364061
transform 1 0 33764 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_365
timestamp 1586364061
transform 1 0 34684 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_382
timestamp 1586364061
transform 1 0 36248 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_394
timestamp 1586364061
transform 1 0 37352 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_33
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _181_
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _182_
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _175_
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_218
timestamp 1586364061
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_233
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_222
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_229
timestamp 1586364061
transform 1 0 22172 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_240
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _131_
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_256
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_277
timestamp 1586364061
transform 1 0 26588 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28796 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_294
timestamp 1586364061
transform 1 0 28152 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_298
timestamp 1586364061
transform 1 0 28520 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_303
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_293
timestamp 1586364061
transform 1 0 28060 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_304
timestamp 1586364061
transform 1 0 29072 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _123_
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_309
timestamp 1586364061
transform 1 0 29532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_313
timestamp 1586364061
transform 1 0 29900 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_316
timestamp 1586364061
transform 1 0 30176 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 30728 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_320
timestamp 1586364061
transform 1 0 30544 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_324
timestamp 1586364061
transform 1 0 30912 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_332
timestamp 1586364061
transform 1 0 31648 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_328
timestamp 1586364061
transform 1 0 31280 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31740 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32752 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32200 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_336
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_340
timestamp 1586364061
transform 1 0 32384 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33396 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_347
timestamp 1586364061
transform 1 0 33028 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_353
timestamp 1586364061
transform 1 0 33580 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_354
timestamp 1586364061
transform 1 0 33672 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34408 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 35144 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 35328 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_365
timestamp 1586364061
transform 1 0 34684 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 35880 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_380
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_377
timestamp 1586364061
transform 1 0 35788 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 36984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37352 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_388
timestamp 1586364061
transform 1 0 36800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_392
timestamp 1586364061
transform 1 0 37168 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_396
timestamp 1586364061
transform 1 0 37536 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_388
timestamp 1586364061
transform 1 0 36800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_396
timestamp 1586364061
transform 1 0 37536 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_404
timestamp 1586364061
transform 1 0 38272 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _168_
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_78
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _073_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_187
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_228
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_274
timestamp 1586364061
transform 1 0 26312 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26680 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27692 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_285
timestamp 1586364061
transform 1 0 27324 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_292
timestamp 1586364061
transform 1 0 27968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_296
timestamp 1586364061
transform 1 0 28336 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_304
timestamp 1586364061
transform 1 0 29072 0 1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_348
timestamp 1586364061
transform 1 0 33120 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_352
timestamp 1586364061
transform 1 0 33488 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_356
timestamp 1586364061
transform 1 0 33856 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 35420 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 35236 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_360
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_363
timestamp 1586364061
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_377
timestamp 1586364061
transform 1 0 35788 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_381
timestamp 1586364061
transform 1 0 36156 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_393
timestamp 1586364061
transform 1 0 37260 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_405
timestamp 1586364061
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_17
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_39
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_161
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_280
timestamp 1586364061
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_292
timestamp 1586364061
transform 1 0 27968 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_304
timestamp 1586364061
transform 1 0 29072 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_316
timestamp 1586364061
transform 1 0 30176 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_328
timestamp 1586364061
transform 1 0 31280 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_364
timestamp 1586364061
transform 1 0 34592 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_372
timestamp 1586364061
transform 1 0 35328 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_17
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_21
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_17_54
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_65
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 590 592
use scs8hd_buf_1  _108_
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_233
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_35
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_55
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _176_
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_48
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_381
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_405
timestamp 1586364061
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 3422 0 3478 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 5814 0 5870 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 8114 0 8170 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 10506 0 10562 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 12806 0 12862 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 15198 0 15254 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 17590 0 17646 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 22282 0 22338 480 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 34058 0 34114 480 6 bottom_grid_pin_10_
port 8 nsew default tristate
rlabel metal2 s 36358 0 36414 480 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal2 s 38750 0 38806 480 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 bottom_grid_pin_2_
port 11 nsew default tristate
rlabel metal2 s 26974 0 27030 480 6 bottom_grid_pin_4_
port 12 nsew default tristate
rlabel metal2 s 29366 0 29422 480 6 bottom_grid_pin_6_
port 13 nsew default tristate
rlabel metal2 s 31666 0 31722 480 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[0]
port 33 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[1]
port 34 nsew default input
rlabel metal3 s 39520 2184 40000 2304 6 chanx_right_in[2]
port 35 nsew default input
rlabel metal3 s 39520 3000 40000 3120 6 chanx_right_in[3]
port 36 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[4]
port 37 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[5]
port 38 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[6]
port 39 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[7]
port 40 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[8]
port 41 nsew default input
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[0]
port 42 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[1]
port 43 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[2]
port 44 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[3]
port 45 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[4]
port 46 nsew default tristate
rlabel metal3 s 39520 12792 40000 12912 6 chanx_right_out[5]
port 47 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[6]
port 48 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[7]
port 49 nsew default tristate
rlabel metal3 s 39520 15512 40000 15632 6 chanx_right_out[8]
port 50 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 data_in
port 51 nsew default input
rlabel metal2 s 1122 0 1178 480 6 enable
port 52 nsew default input
rlabel metal2 s 33322 15520 33378 16000 6 top_grid_pin_14_
port 53 nsew default tristate
rlabel metal2 s 6642 15520 6698 16000 6 top_grid_pin_2_
port 54 nsew default tristate
rlabel metal2 s 19982 15520 20038 16000 6 top_grid_pin_6_
port 55 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 56 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 57 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
