magic
tech EFS8A
magscale 1 2
timestamp 1602874310
<< locali >>
rect 19803 9367 19837 9435
rect 19803 9333 19809 9367
<< viali >>
rect 12909 10217 12943 10251
rect 26709 10217 26743 10251
rect 39405 10217 39439 10251
rect 66361 10217 66395 10251
rect 79885 10217 79919 10251
rect 49617 10149 49651 10183
rect 10425 10081 10459 10115
rect 11069 10081 11103 10115
rect 12725 10081 12759 10115
rect 21833 10081 21867 10115
rect 26525 10081 26559 10115
rect 35633 10081 35667 10115
rect 39221 10081 39255 10115
rect 48973 10081 49007 10115
rect 52745 10081 52779 10115
rect 61485 10081 61519 10115
rect 62129 10081 62163 10115
rect 66177 10081 66211 10115
rect 79701 10081 79735 10115
rect 88441 10081 88475 10115
rect 1409 10013 1443 10047
rect 1593 10013 1627 10047
rect 10609 10013 10643 10047
rect 22017 10013 22051 10047
rect 34989 10013 35023 10047
rect 35173 10013 35207 10047
rect 49157 10013 49191 10047
rect 61669 10013 61703 10047
rect 75101 10013 75135 10047
rect 75285 10013 75319 10047
rect 88257 10013 88291 10047
rect 2053 9877 2087 9911
rect 22477 9877 22511 9911
rect 36185 9877 36219 9911
rect 52929 9877 52963 9911
rect 75745 9877 75779 9911
rect 88717 9877 88751 9911
rect 2697 9673 2731 9707
rect 10425 9673 10459 9707
rect 21833 9673 21867 9707
rect 49065 9673 49099 9707
rect 52745 9673 52779 9707
rect 61577 9673 61611 9707
rect 89085 9673 89119 9707
rect 2421 9605 2455 9639
rect 20361 9605 20395 9639
rect 22201 9605 22235 9639
rect 35173 9605 35207 9639
rect 75193 9605 75227 9639
rect 61853 9537 61887 9571
rect 1409 9469 1443 9503
rect 19441 9469 19475 9503
rect 36185 9469 36219 9503
rect 37105 9469 37139 9503
rect 88073 9469 88107 9503
rect 2053 9401 2087 9435
rect 36506 9401 36540 9435
rect 1593 9333 1627 9367
rect 10885 9333 10919 9367
rect 12725 9333 12759 9367
rect 19349 9333 19383 9367
rect 19809 9333 19843 9367
rect 26617 9333 26651 9367
rect 35449 9333 35483 9367
rect 36093 9333 36127 9367
rect 39313 9333 39347 9367
rect 49341 9333 49375 9367
rect 66269 9333 66303 9367
rect 75469 9333 75503 9367
rect 79977 9333 80011 9367
rect 87889 9333 87923 9367
rect 88257 9333 88291 9367
rect 88717 9333 88751 9367
rect 2329 9129 2363 9163
rect 11805 9129 11839 9163
rect 21833 9129 21867 9163
rect 33057 9129 33091 9163
rect 38669 9129 38703 9163
rect 1730 9061 1764 9095
rect 11247 9061 11281 9095
rect 21925 9061 21959 9095
rect 22017 9061 22051 9095
rect 22385 9061 22419 9095
rect 32458 9061 32492 9095
rect 36230 9061 36264 9095
rect 38070 9061 38104 9095
rect 36829 8993 36863 9027
rect 1409 8925 1443 8959
rect 10885 8925 10919 8959
rect 21649 8925 21683 8959
rect 32137 8925 32171 8959
rect 35909 8925 35943 8959
rect 37749 8925 37783 8959
rect 9965 8789 9999 8823
rect 13093 8789 13127 8823
rect 19533 8789 19567 8823
rect 19809 8789 19843 8823
rect 1593 8585 1627 8619
rect 11437 8585 11471 8619
rect 32505 8585 32539 8619
rect 22017 8517 22051 8551
rect 12173 8449 12207 8483
rect 19625 8449 19659 8483
rect 35449 8449 35483 8483
rect 9689 8381 9723 8415
rect 10149 8381 10183 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 12817 8381 12851 8415
rect 13277 8381 13311 8415
rect 13461 8381 13495 8415
rect 13829 8381 13863 8415
rect 14197 8381 14231 8415
rect 15301 8381 15335 8415
rect 15761 8381 15795 8415
rect 19809 8381 19843 8415
rect 20269 8381 20303 8415
rect 20821 8381 20855 8415
rect 21005 8381 21039 8415
rect 21281 8381 21315 8415
rect 36369 8381 36403 8415
rect 37289 8381 37323 8415
rect 36690 8313 36724 8347
rect 38117 8313 38151 8347
rect 2053 8245 2087 8279
rect 9137 8245 9171 8279
rect 9505 8245 9539 8279
rect 9781 8245 9815 8279
rect 13093 8245 13127 8279
rect 15485 8245 15519 8279
rect 19349 8245 19383 8279
rect 21649 8245 21683 8279
rect 22385 8245 22419 8279
rect 22845 8245 22879 8279
rect 32137 8245 32171 8279
rect 35817 8245 35851 8279
rect 36185 8245 36219 8279
rect 37749 8245 37783 8279
rect 10977 8041 11011 8075
rect 19533 8041 19567 8075
rect 23213 8041 23247 8075
rect 36369 8041 36403 8075
rect 9965 7973 9999 8007
rect 13001 7973 13035 8007
rect 21741 7973 21775 8007
rect 22109 7973 22143 8007
rect 23305 7973 23339 8007
rect 23673 7973 23707 8007
rect 18337 7905 18371 7939
rect 18797 7905 18831 7939
rect 19165 7905 19199 7939
rect 19625 7905 19659 7939
rect 21557 7905 21591 7939
rect 21649 7905 21683 7939
rect 23121 7905 23155 7939
rect 21373 7837 21407 7871
rect 22937 7837 22971 7871
rect 20085 7701 20119 7735
rect 21281 7701 21315 7735
rect 17417 7497 17451 7531
rect 19809 7497 19843 7531
rect 20637 7497 20671 7531
rect 21005 7497 21039 7531
rect 22201 7497 22235 7531
rect 22937 7497 22971 7531
rect 23305 7497 23339 7531
rect 17785 7429 17819 7463
rect 18245 7429 18279 7463
rect 19533 7429 19567 7463
rect 22569 7429 22603 7463
rect 21925 7361 21959 7395
rect 18521 7293 18555 7327
rect 21373 7293 21407 7327
rect 21541 7293 21575 7327
rect 18429 7225 18463 7259
rect 20361 7225 20395 7259
rect 21189 7225 21223 7259
rect 21465 7157 21499 7191
rect 18797 6953 18831 6987
rect 20637 6953 20671 6987
rect 23305 6953 23339 6987
rect 21649 6885 21683 6919
rect 18429 6817 18463 6851
rect 21005 6817 21039 6851
rect 22937 6817 22971 6851
rect 21925 6749 21959 6783
rect 21005 6409 21039 6443
rect 18337 6069 18371 6103
<< metal1 >>
rect 1104 11450 106812 11472
rect 1104 11398 36982 11450
rect 37034 11398 37046 11450
rect 37098 11398 37110 11450
rect 37162 11398 37174 11450
rect 37226 11398 72982 11450
rect 73034 11398 73046 11450
rect 73098 11398 73110 11450
rect 73162 11398 73174 11450
rect 73226 11398 106812 11450
rect 1104 11376 106812 11398
rect 1104 10906 106812 10928
rect 1104 10854 18982 10906
rect 19034 10854 19046 10906
rect 19098 10854 19110 10906
rect 19162 10854 19174 10906
rect 19226 10854 54982 10906
rect 55034 10854 55046 10906
rect 55098 10854 55110 10906
rect 55162 10854 55174 10906
rect 55226 10854 90982 10906
rect 91034 10854 91046 10906
rect 91098 10854 91110 10906
rect 91162 10854 91174 10906
rect 91226 10854 106812 10906
rect 1104 10832 106812 10854
rect 1104 10362 106812 10384
rect 1104 10310 36982 10362
rect 37034 10310 37046 10362
rect 37098 10310 37110 10362
rect 37162 10310 37174 10362
rect 37226 10310 72982 10362
rect 73034 10310 73046 10362
rect 73098 10310 73110 10362
rect 73162 10310 73174 10362
rect 73226 10310 106812 10362
rect 1104 10288 106812 10310
rect 12894 10248 12900 10260
rect 12855 10220 12900 10248
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 26694 10248 26700 10260
rect 26655 10220 26700 10248
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 39390 10248 39396 10260
rect 39351 10220 39396 10248
rect 39390 10208 39396 10220
rect 39448 10208 39454 10260
rect 66346 10248 66352 10260
rect 66307 10220 66352 10248
rect 66346 10208 66352 10220
rect 66404 10208 66410 10260
rect 79870 10248 79876 10260
rect 79831 10220 79876 10248
rect 79870 10208 79876 10220
rect 79928 10208 79934 10260
rect 16758 10180 16764 10192
rect 10428 10152 16764 10180
rect 10428 10124 10456 10152
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 49605 10183 49663 10189
rect 49605 10149 49617 10183
rect 49651 10180 49663 10183
rect 49651 10152 52408 10180
rect 49651 10149 49663 10152
rect 49605 10143 49663 10149
rect 52380 10124 52408 10152
rect 10410 10112 10416 10124
rect 10323 10084 10416 10112
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 12710 10112 12716 10124
rect 11103 10084 12716 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 21818 10112 21824 10124
rect 21779 10084 21824 10112
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 26513 10115 26571 10121
rect 26513 10081 26525 10115
rect 26559 10112 26571 10115
rect 26602 10112 26608 10124
rect 26559 10084 26608 10112
rect 26559 10081 26571 10084
rect 26513 10075 26571 10081
rect 26602 10072 26608 10084
rect 26660 10072 26666 10124
rect 35621 10115 35679 10121
rect 35621 10081 35633 10115
rect 35667 10112 35679 10115
rect 39209 10115 39267 10121
rect 39209 10112 39221 10115
rect 35667 10084 39221 10112
rect 35667 10081 35679 10084
rect 35621 10075 35679 10081
rect 39209 10081 39221 10084
rect 39255 10112 39267 10115
rect 39298 10112 39304 10124
rect 39255 10084 39304 10112
rect 39255 10081 39267 10084
rect 39209 10075 39267 10081
rect 39298 10072 39304 10084
rect 39356 10072 39362 10124
rect 48961 10115 49019 10121
rect 48961 10081 48973 10115
rect 49007 10112 49019 10115
rect 49050 10112 49056 10124
rect 49007 10084 49056 10112
rect 49007 10081 49019 10084
rect 48961 10075 49019 10081
rect 49050 10072 49056 10084
rect 49108 10112 49114 10124
rect 49108 10084 50108 10112
rect 49108 10072 49114 10084
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10044 10655 10047
rect 10870 10044 10876 10056
rect 10643 10016 10876 10044
rect 10643 10013 10655 10016
rect 10597 10007 10655 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 22002 10044 22008 10056
rect 21963 10016 22008 10044
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 34977 10047 35035 10053
rect 34977 10013 34989 10047
rect 35023 10044 35035 10047
rect 35066 10044 35072 10056
rect 35023 10016 35072 10044
rect 35023 10013 35035 10016
rect 34977 10007 35035 10013
rect 35066 10004 35072 10016
rect 35124 10004 35130 10056
rect 35161 10047 35219 10053
rect 35161 10013 35173 10047
rect 35207 10044 35219 10047
rect 35434 10044 35440 10056
rect 35207 10016 35440 10044
rect 35207 10013 35219 10016
rect 35161 10007 35219 10013
rect 35434 10004 35440 10016
rect 35492 10004 35498 10056
rect 49145 10047 49203 10053
rect 49145 10013 49157 10047
rect 49191 10044 49203 10047
rect 49326 10044 49332 10056
rect 49191 10016 49332 10044
rect 49191 10013 49203 10016
rect 49145 10007 49203 10013
rect 49326 10004 49332 10016
rect 49384 10004 49390 10056
rect 50080 10044 50108 10084
rect 52362 10072 52368 10124
rect 52420 10112 52426 10124
rect 52730 10112 52736 10124
rect 52420 10084 52736 10112
rect 52420 10072 52426 10084
rect 52730 10072 52736 10084
rect 52788 10072 52794 10124
rect 61473 10115 61531 10121
rect 61473 10081 61485 10115
rect 61519 10112 61531 10115
rect 61562 10112 61568 10124
rect 61519 10084 61568 10112
rect 61519 10081 61531 10084
rect 61473 10075 61531 10081
rect 61562 10072 61568 10084
rect 61620 10112 61626 10124
rect 62117 10115 62175 10121
rect 61620 10084 61792 10112
rect 61620 10072 61626 10084
rect 57330 10044 57336 10056
rect 50080 10016 57336 10044
rect 57330 10004 57336 10016
rect 57388 10004 57394 10056
rect 61657 10047 61715 10053
rect 61657 10013 61669 10047
rect 61703 10013 61715 10047
rect 61764 10044 61792 10084
rect 62117 10081 62129 10115
rect 62163 10112 62175 10115
rect 66165 10115 66223 10121
rect 66165 10112 66177 10115
rect 62163 10084 66177 10112
rect 62163 10081 62175 10084
rect 62117 10075 62175 10081
rect 66165 10081 66177 10084
rect 66211 10112 66223 10115
rect 66254 10112 66260 10124
rect 66211 10084 66260 10112
rect 66211 10081 66223 10084
rect 66165 10075 66223 10081
rect 66254 10072 66260 10084
rect 66312 10072 66318 10124
rect 79686 10112 79692 10124
rect 79647 10084 79692 10112
rect 79686 10072 79692 10084
rect 79744 10072 79750 10124
rect 87874 10072 87880 10124
rect 87932 10112 87938 10124
rect 88429 10115 88487 10121
rect 88429 10112 88441 10115
rect 87932 10084 88441 10112
rect 87932 10072 87938 10084
rect 88429 10081 88441 10084
rect 88475 10081 88487 10115
rect 88429 10075 88487 10081
rect 70762 10044 70768 10056
rect 61764 10016 70768 10044
rect 61657 10007 61715 10013
rect 61672 9976 61700 10007
rect 70762 10004 70768 10016
rect 70820 10004 70826 10056
rect 75089 10047 75147 10053
rect 75089 10013 75101 10047
rect 75135 10044 75147 10047
rect 75178 10044 75184 10056
rect 75135 10016 75184 10044
rect 75135 10013 75147 10016
rect 75089 10007 75147 10013
rect 75178 10004 75184 10016
rect 75236 10004 75242 10056
rect 75273 10047 75331 10053
rect 75273 10013 75285 10047
rect 75319 10044 75331 10047
rect 75454 10044 75460 10056
rect 75319 10016 75460 10044
rect 75319 10013 75331 10016
rect 75273 10007 75331 10013
rect 75454 10004 75460 10016
rect 75512 10004 75518 10056
rect 88245 10047 88303 10053
rect 88245 10013 88257 10047
rect 88291 10044 88303 10047
rect 89070 10044 89076 10056
rect 88291 10016 89076 10044
rect 88291 10013 88303 10016
rect 88245 10007 88303 10013
rect 89070 10004 89076 10016
rect 89128 10004 89134 10056
rect 61838 9976 61844 9988
rect 61672 9948 61844 9976
rect 61838 9936 61844 9948
rect 61896 9936 61902 9988
rect 2038 9908 2044 9920
rect 1999 9880 2044 9908
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 22465 9911 22523 9917
rect 22465 9877 22477 9911
rect 22511 9908 22523 9911
rect 23382 9908 23388 9920
rect 22511 9880 23388 9908
rect 22511 9877 22523 9880
rect 22465 9871 22523 9877
rect 23382 9868 23388 9880
rect 23440 9868 23446 9920
rect 36170 9908 36176 9920
rect 36131 9880 36176 9908
rect 36170 9868 36176 9880
rect 36228 9868 36234 9920
rect 52917 9911 52975 9917
rect 52917 9877 52929 9911
rect 52963 9908 52975 9911
rect 61470 9908 61476 9920
rect 52963 9880 61476 9908
rect 52963 9877 52975 9880
rect 52917 9871 52975 9877
rect 61470 9868 61476 9880
rect 61528 9868 61534 9920
rect 75733 9911 75791 9917
rect 75733 9877 75745 9911
rect 75779 9908 75791 9911
rect 78582 9908 78588 9920
rect 75779 9880 78588 9908
rect 75779 9877 75791 9880
rect 75733 9871 75791 9877
rect 78582 9868 78588 9880
rect 78640 9868 78646 9920
rect 88702 9908 88708 9920
rect 88663 9880 88708 9908
rect 88702 9868 88708 9880
rect 88760 9868 88766 9920
rect 1104 9818 106812 9840
rect 1104 9766 18982 9818
rect 19034 9766 19046 9818
rect 19098 9766 19110 9818
rect 19162 9766 19174 9818
rect 19226 9766 54982 9818
rect 55034 9766 55046 9818
rect 55098 9766 55110 9818
rect 55162 9766 55174 9818
rect 55226 9766 90982 9818
rect 91034 9766 91046 9818
rect 91098 9766 91110 9818
rect 91162 9766 91174 9818
rect 91226 9766 106812 9818
rect 1104 9744 106812 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 2314 9704 2320 9716
rect 1636 9676 2320 9704
rect 1636 9664 1642 9676
rect 2314 9664 2320 9676
rect 2372 9704 2378 9716
rect 2685 9707 2743 9713
rect 2685 9704 2697 9707
rect 2372 9676 2697 9704
rect 2372 9664 2378 9676
rect 2685 9673 2697 9676
rect 2731 9673 2743 9707
rect 10410 9704 10416 9716
rect 10371 9676 10416 9704
rect 2685 9667 2743 9673
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 21818 9704 21824 9716
rect 21779 9676 21824 9704
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 49050 9704 49056 9716
rect 49011 9676 49056 9704
rect 49050 9664 49056 9676
rect 49108 9664 49114 9716
rect 52730 9704 52736 9716
rect 52691 9676 52736 9704
rect 52730 9664 52736 9676
rect 52788 9664 52794 9716
rect 61562 9704 61568 9716
rect 61523 9676 61568 9704
rect 61562 9664 61568 9676
rect 61620 9664 61626 9716
rect 89070 9704 89076 9716
rect 89031 9676 89076 9704
rect 89070 9664 89076 9676
rect 89128 9664 89134 9716
rect 1394 9596 1400 9648
rect 1452 9636 1458 9648
rect 2409 9639 2467 9645
rect 2409 9636 2421 9639
rect 1452 9608 2421 9636
rect 1452 9596 1458 9608
rect 2409 9605 2421 9608
rect 2455 9636 2467 9639
rect 3326 9636 3332 9648
rect 2455 9608 3332 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 20349 9639 20407 9645
rect 20349 9605 20361 9639
rect 20395 9636 20407 9639
rect 22002 9636 22008 9648
rect 20395 9608 22008 9636
rect 20395 9605 20407 9608
rect 20349 9599 20407 9605
rect 22002 9596 22008 9608
rect 22060 9636 22066 9648
rect 22189 9639 22247 9645
rect 22189 9636 22201 9639
rect 22060 9608 22201 9636
rect 22060 9596 22066 9608
rect 22189 9605 22201 9608
rect 22235 9605 22247 9639
rect 22189 9599 22247 9605
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 26602 9636 26608 9648
rect 23440 9608 26608 9636
rect 23440 9596 23446 9608
rect 26602 9596 26608 9608
rect 26660 9596 26666 9648
rect 35158 9636 35164 9648
rect 35119 9608 35164 9636
rect 35158 9596 35164 9608
rect 35216 9596 35222 9648
rect 75178 9636 75184 9648
rect 75139 9608 75184 9636
rect 75178 9596 75184 9608
rect 75236 9596 75242 9648
rect 61838 9568 61844 9580
rect 61799 9540 61844 9568
rect 61838 9528 61844 9540
rect 61896 9528 61902 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19518 9500 19524 9512
rect 19475 9472 19524 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 1412 9432 1440 9463
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 36170 9500 36176 9512
rect 36131 9472 36176 9500
rect 36170 9460 36176 9472
rect 36228 9460 36234 9512
rect 37093 9503 37151 9509
rect 37093 9469 37105 9503
rect 37139 9500 37151 9503
rect 39942 9500 39948 9512
rect 37139 9472 39948 9500
rect 37139 9469 37151 9472
rect 37093 9463 37151 9469
rect 39942 9460 39948 9472
rect 40000 9460 40006 9512
rect 88061 9503 88119 9509
rect 88061 9469 88073 9503
rect 88107 9500 88119 9503
rect 88702 9500 88708 9512
rect 88107 9472 88708 9500
rect 88107 9469 88119 9472
rect 88061 9463 88119 9469
rect 88702 9460 88708 9472
rect 88760 9460 88766 9512
rect 2038 9432 2044 9444
rect 1412 9404 2044 9432
rect 2038 9392 2044 9404
rect 2096 9432 2102 9444
rect 6454 9432 6460 9444
rect 2096 9404 6460 9432
rect 2096 9392 2102 9404
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 36494 9435 36552 9441
rect 36494 9432 36506 9435
rect 36096 9404 36506 9432
rect 36096 9376 36124 9404
rect 36494 9401 36506 9404
rect 36540 9401 36552 9435
rect 36494 9395 36552 9401
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 1670 9364 1676 9376
rect 1627 9336 1676 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 10870 9364 10876 9376
rect 10831 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 12710 9364 12716 9376
rect 12671 9336 12716 9364
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 19337 9367 19395 9373
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 19794 9364 19800 9376
rect 19383 9336 19800 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 26602 9364 26608 9376
rect 26563 9336 26608 9364
rect 26602 9324 26608 9336
rect 26660 9324 26666 9376
rect 35434 9364 35440 9376
rect 35395 9336 35440 9364
rect 35434 9324 35440 9336
rect 35492 9324 35498 9376
rect 36078 9364 36084 9376
rect 36039 9336 36084 9364
rect 36078 9324 36084 9336
rect 36136 9324 36142 9376
rect 39298 9364 39304 9376
rect 39259 9336 39304 9364
rect 39298 9324 39304 9336
rect 39356 9324 39362 9376
rect 49326 9364 49332 9376
rect 49287 9336 49332 9364
rect 49326 9324 49332 9336
rect 49384 9324 49390 9376
rect 66254 9364 66260 9376
rect 66215 9336 66260 9364
rect 66254 9324 66260 9336
rect 66312 9324 66318 9376
rect 75454 9364 75460 9376
rect 75415 9336 75460 9364
rect 75454 9324 75460 9336
rect 75512 9324 75518 9376
rect 78582 9324 78588 9376
rect 78640 9364 78646 9376
rect 79686 9364 79692 9376
rect 78640 9336 79692 9364
rect 78640 9324 78646 9336
rect 79686 9324 79692 9336
rect 79744 9364 79750 9376
rect 79965 9367 80023 9373
rect 79965 9364 79977 9367
rect 79744 9336 79977 9364
rect 79744 9324 79750 9336
rect 79965 9333 79977 9336
rect 80011 9333 80023 9367
rect 87874 9364 87880 9376
rect 87835 9336 87880 9364
rect 79965 9327 80023 9333
rect 87874 9324 87880 9336
rect 87932 9324 87938 9376
rect 88242 9364 88248 9376
rect 88203 9336 88248 9364
rect 88242 9324 88248 9336
rect 88300 9324 88306 9376
rect 88702 9364 88708 9376
rect 88663 9336 88708 9364
rect 88702 9324 88708 9336
rect 88760 9324 88766 9376
rect 1104 9274 106812 9296
rect 1104 9222 36982 9274
rect 37034 9222 37046 9274
rect 37098 9222 37110 9274
rect 37162 9222 37174 9274
rect 37226 9222 72982 9274
rect 73034 9222 73046 9274
rect 73098 9222 73110 9274
rect 73162 9222 73174 9274
rect 73226 9222 106812 9274
rect 1104 9200 106812 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 10928 9132 11805 9160
rect 10928 9120 10934 9132
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 21818 9160 21824 9172
rect 21779 9132 21824 9160
rect 11793 9123 11851 9129
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 33045 9163 33103 9169
rect 33045 9129 33057 9163
rect 33091 9160 33103 9163
rect 35434 9160 35440 9172
rect 33091 9132 35440 9160
rect 33091 9129 33103 9132
rect 33045 9123 33103 9129
rect 35434 9120 35440 9132
rect 35492 9120 35498 9172
rect 38657 9163 38715 9169
rect 38657 9129 38669 9163
rect 38703 9160 38715 9163
rect 49326 9160 49332 9172
rect 38703 9132 49332 9160
rect 38703 9129 38715 9132
rect 38657 9123 38715 9129
rect 49326 9120 49332 9132
rect 49384 9120 49390 9172
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 1718 9095 1776 9101
rect 1718 9092 1730 9095
rect 1544 9064 1730 9092
rect 1544 9052 1550 9064
rect 1718 9061 1730 9064
rect 1764 9061 1776 9095
rect 1718 9055 1776 9061
rect 11235 9095 11293 9101
rect 11235 9061 11247 9095
rect 11281 9092 11293 9095
rect 11422 9092 11428 9104
rect 11281 9064 11428 9092
rect 11281 9061 11293 9064
rect 11235 9055 11293 9061
rect 11422 9052 11428 9064
rect 11480 9052 11486 9104
rect 21910 9092 21916 9104
rect 21871 9064 21916 9092
rect 21910 9052 21916 9064
rect 21968 9052 21974 9104
rect 22005 9095 22063 9101
rect 22005 9061 22017 9095
rect 22051 9092 22063 9095
rect 22094 9092 22100 9104
rect 22051 9064 22100 9092
rect 22051 9061 22063 9064
rect 22005 9055 22063 9061
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 22373 9095 22431 9101
rect 22373 9061 22385 9095
rect 22419 9092 22431 9095
rect 23290 9092 23296 9104
rect 22419 9064 23296 9092
rect 22419 9061 22431 9064
rect 22373 9055 22431 9061
rect 23290 9052 23296 9064
rect 23348 9052 23354 9104
rect 32122 9052 32128 9104
rect 32180 9092 32186 9104
rect 32446 9095 32504 9101
rect 32446 9092 32458 9095
rect 32180 9064 32458 9092
rect 32180 9052 32186 9064
rect 32446 9061 32458 9064
rect 32492 9061 32504 9095
rect 32446 9055 32504 9061
rect 36078 9052 36084 9104
rect 36136 9092 36142 9104
rect 36218 9095 36276 9101
rect 36218 9092 36230 9095
rect 36136 9064 36230 9092
rect 36136 9052 36142 9064
rect 36218 9061 36230 9064
rect 36264 9092 36276 9095
rect 38058 9095 38116 9101
rect 38058 9092 38070 9095
rect 36264 9064 38070 9092
rect 36264 9061 36276 9064
rect 36218 9055 36276 9061
rect 38058 9061 38070 9064
rect 38104 9061 38116 9095
rect 38058 9055 38116 9061
rect 36817 9027 36875 9033
rect 36817 8993 36829 9027
rect 36863 9024 36875 9027
rect 39758 9024 39764 9036
rect 36863 8996 39764 9024
rect 36863 8993 36875 8996
rect 36817 8987 36875 8993
rect 39758 8984 39764 8996
rect 39816 8984 39822 9036
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2038 8956 2044 8968
rect 1443 8928 2044 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 10870 8956 10876 8968
rect 10831 8928 10876 8956
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 21634 8956 21640 8968
rect 21595 8928 21640 8956
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 32125 8959 32183 8965
rect 32125 8925 32137 8959
rect 32171 8956 32183 8959
rect 32490 8956 32496 8968
rect 32171 8928 32496 8956
rect 32171 8925 32183 8928
rect 32125 8919 32183 8925
rect 32490 8916 32496 8928
rect 32548 8916 32554 8968
rect 35434 8916 35440 8968
rect 35492 8956 35498 8968
rect 35897 8959 35955 8965
rect 35897 8956 35909 8959
rect 35492 8928 35909 8956
rect 35492 8916 35498 8928
rect 35897 8925 35909 8928
rect 35943 8925 35955 8959
rect 35897 8919 35955 8925
rect 37642 8916 37648 8968
rect 37700 8956 37706 8968
rect 37737 8959 37795 8965
rect 37737 8956 37749 8959
rect 37700 8928 37749 8956
rect 37700 8916 37706 8928
rect 37737 8925 37749 8928
rect 37783 8925 37795 8959
rect 37737 8919 37795 8925
rect 9950 8820 9956 8832
rect 9911 8792 9956 8820
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 13081 8823 13139 8829
rect 13081 8789 13093 8823
rect 13127 8820 13139 8823
rect 13262 8820 13268 8832
rect 13127 8792 13268 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 19518 8820 19524 8832
rect 19479 8792 19524 8820
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 19760 8792 19809 8820
rect 19760 8780 19766 8792
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 19797 8783 19855 8789
rect 1104 8730 106812 8752
rect 1104 8678 18982 8730
rect 19034 8678 19046 8730
rect 19098 8678 19110 8730
rect 19162 8678 19174 8730
rect 19226 8678 54982 8730
rect 55034 8678 55046 8730
rect 55098 8678 55110 8730
rect 55162 8678 55174 8730
rect 55226 8678 90982 8730
rect 91034 8678 91046 8730
rect 91098 8678 91110 8730
rect 91162 8678 91174 8730
rect 91226 8678 106812 8730
rect 1104 8656 106812 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 11422 8616 11428 8628
rect 11383 8588 11428 8616
rect 1581 8579 1639 8585
rect 11422 8576 11428 8588
rect 11480 8616 11486 8628
rect 19794 8616 19800 8628
rect 11480 8588 19800 8616
rect 11480 8576 11486 8588
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 21910 8576 21916 8628
rect 21968 8576 21974 8628
rect 32490 8616 32496 8628
rect 32451 8588 32496 8616
rect 32490 8576 32496 8588
rect 32548 8576 32554 8628
rect 21928 8548 21956 8576
rect 22005 8551 22063 8557
rect 22005 8548 22017 8551
rect 19306 8520 22017 8548
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 12161 8483 12219 8489
rect 12161 8480 12173 8483
rect 9548 8452 9720 8480
rect 9548 8440 9554 8452
rect 9692 8421 9720 8452
rect 10152 8452 12173 8480
rect 9677 8415 9735 8421
rect 4126 8384 9628 8412
rect 2038 8276 2044 8288
rect 1951 8248 2044 8276
rect 2038 8236 2044 8248
rect 2096 8276 2102 8288
rect 4126 8276 4154 8384
rect 9122 8276 9128 8288
rect 2096 8248 4154 8276
rect 9083 8248 9128 8276
rect 2096 8236 2102 8248
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9490 8276 9496 8288
rect 9451 8248 9496 8276
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9600 8276 9628 8384
rect 9677 8381 9689 8415
rect 9723 8381 9735 8415
rect 9677 8375 9735 8381
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10152 8421 10180 8452
rect 12161 8449 12173 8452
rect 12207 8480 12219 8483
rect 18782 8480 18788 8492
rect 12207 8452 18788 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 10008 8384 10149 8412
rect 10008 8372 10014 8384
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10686 8412 10692 8424
rect 10647 8384 10692 8412
rect 10137 8375 10195 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 10836 8384 10885 8412
rect 10836 8372 10842 8384
rect 10873 8381 10885 8384
rect 10919 8412 10931 8415
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 10919 8384 12817 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 13262 8412 13268 8424
rect 13223 8384 13268 8412
rect 12805 8375 12863 8381
rect 12820 8344 12848 8375
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13464 8421 13492 8452
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8381 13507 8415
rect 13449 8375 13507 8381
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 14185 8415 14243 8421
rect 13872 8384 13917 8412
rect 13872 8372 13878 8384
rect 14185 8381 14197 8415
rect 14231 8381 14243 8415
rect 15286 8412 15292 8424
rect 15247 8384 15292 8412
rect 14185 8375 14243 8381
rect 14200 8344 14228 8375
rect 15286 8372 15292 8384
rect 15344 8412 15350 8424
rect 15749 8415 15807 8421
rect 15749 8412 15761 8415
rect 15344 8384 15761 8412
rect 15344 8372 15350 8384
rect 15749 8381 15761 8384
rect 15795 8412 15807 8415
rect 19306 8412 19334 8520
rect 22005 8517 22017 8520
rect 22051 8548 22063 8551
rect 23198 8548 23204 8560
rect 22051 8520 23204 8548
rect 22051 8517 22063 8520
rect 22005 8511 22063 8517
rect 23198 8508 23204 8520
rect 23256 8508 23262 8560
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 19484 8452 19625 8480
rect 19484 8440 19490 8452
rect 19613 8449 19625 8452
rect 19659 8480 19671 8483
rect 22094 8480 22100 8492
rect 19659 8452 20852 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 20824 8424 20852 8452
rect 21008 8452 22100 8480
rect 15795 8384 19334 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 19702 8372 19708 8424
rect 19760 8412 19766 8424
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 19760 8384 19809 8412
rect 19760 8372 19766 8384
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 19797 8375 19855 8381
rect 20070 8372 20076 8424
rect 20128 8412 20134 8424
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 20128 8384 20269 8412
rect 20128 8372 20134 8384
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 20806 8412 20812 8424
rect 20767 8384 20812 8412
rect 20257 8375 20315 8381
rect 20806 8372 20812 8384
rect 20864 8372 20870 8424
rect 21008 8421 21036 8452
rect 22094 8440 22100 8452
rect 22152 8480 22158 8492
rect 35434 8480 35440 8492
rect 22152 8452 22876 8480
rect 35395 8452 35440 8480
rect 22152 8440 22158 8452
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8381 21051 8415
rect 21266 8412 21272 8424
rect 21227 8384 21272 8412
rect 20993 8375 21051 8381
rect 20530 8344 20536 8356
rect 12820 8316 20536 8344
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 9769 8279 9827 8285
rect 9769 8276 9781 8279
rect 9600 8248 9781 8276
rect 9769 8245 9781 8248
rect 9815 8245 9827 8279
rect 13078 8276 13084 8288
rect 13039 8248 13084 8276
rect 9769 8239 9827 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 15470 8276 15476 8288
rect 13872 8248 15476 8276
rect 13872 8236 13878 8248
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 19337 8279 19395 8285
rect 19337 8245 19349 8279
rect 19383 8276 19395 8279
rect 19610 8276 19616 8288
rect 19383 8248 19616 8276
rect 19383 8245 19395 8248
rect 19337 8239 19395 8245
rect 19610 8236 19616 8248
rect 19668 8276 19674 8288
rect 21008 8276 21036 8375
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21634 8276 21640 8288
rect 19668 8248 21036 8276
rect 21595 8248 21640 8276
rect 19668 8236 19674 8248
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 21818 8236 21824 8288
rect 21876 8276 21882 8288
rect 22848 8285 22876 8452
rect 35434 8440 35440 8452
rect 35492 8440 35498 8492
rect 36354 8412 36360 8424
rect 36315 8384 36360 8412
rect 36354 8372 36360 8384
rect 36412 8372 36418 8424
rect 37277 8415 37335 8421
rect 37277 8381 37289 8415
rect 37323 8412 37335 8415
rect 40034 8412 40040 8424
rect 37323 8384 40040 8412
rect 37323 8381 37335 8384
rect 37277 8375 37335 8381
rect 40034 8372 40040 8384
rect 40092 8372 40098 8424
rect 36678 8347 36736 8353
rect 36678 8344 36690 8347
rect 36188 8316 36690 8344
rect 22373 8279 22431 8285
rect 22373 8276 22385 8279
rect 21876 8248 22385 8276
rect 21876 8236 21882 8248
rect 22373 8245 22385 8248
rect 22419 8245 22431 8279
rect 22373 8239 22431 8245
rect 22833 8279 22891 8285
rect 22833 8245 22845 8279
rect 22879 8276 22891 8279
rect 23290 8276 23296 8288
rect 22879 8248 23296 8276
rect 22879 8245 22891 8248
rect 22833 8239 22891 8245
rect 23290 8236 23296 8248
rect 23348 8236 23354 8288
rect 32122 8276 32128 8288
rect 32083 8248 32128 8276
rect 32122 8236 32128 8248
rect 32180 8276 32186 8288
rect 35805 8279 35863 8285
rect 35805 8276 35817 8279
rect 32180 8248 35817 8276
rect 32180 8236 32186 8248
rect 35805 8245 35817 8248
rect 35851 8276 35863 8279
rect 36078 8276 36084 8288
rect 35851 8248 36084 8276
rect 35851 8245 35863 8248
rect 35805 8239 35863 8245
rect 36078 8236 36084 8248
rect 36136 8276 36142 8288
rect 36188 8285 36216 8316
rect 36678 8313 36690 8316
rect 36724 8313 36736 8347
rect 36678 8307 36736 8313
rect 36173 8279 36231 8285
rect 36173 8276 36185 8279
rect 36136 8248 36185 8276
rect 36136 8236 36142 8248
rect 36173 8245 36185 8248
rect 36219 8245 36231 8279
rect 36693 8276 36721 8307
rect 36814 8304 36820 8356
rect 36872 8344 36878 8356
rect 37642 8344 37648 8356
rect 36872 8316 37648 8344
rect 36872 8304 36878 8316
rect 37642 8304 37648 8316
rect 37700 8344 37706 8356
rect 38105 8347 38163 8353
rect 38105 8344 38117 8347
rect 37700 8316 38117 8344
rect 37700 8304 37706 8316
rect 38105 8313 38117 8316
rect 38151 8313 38163 8347
rect 38105 8307 38163 8313
rect 37737 8279 37795 8285
rect 37737 8276 37749 8279
rect 36693 8248 37749 8276
rect 36173 8239 36231 8245
rect 37737 8245 37749 8248
rect 37783 8245 37795 8279
rect 37737 8239 37795 8245
rect 1104 8186 106812 8208
rect 1104 8134 36982 8186
rect 37034 8134 37046 8186
rect 37098 8134 37110 8186
rect 37162 8134 37174 8186
rect 37226 8134 72982 8186
rect 73034 8134 73046 8186
rect 73098 8134 73110 8186
rect 73162 8134 73174 8186
rect 73226 8134 106812 8186
rect 1104 8112 106812 8134
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10928 8044 10977 8072
rect 10928 8032 10934 8044
rect 10965 8041 10977 8044
rect 11011 8072 11023 8075
rect 13078 8072 13084 8084
rect 11011 8044 13084 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 19518 8072 19524 8084
rect 19479 8044 19524 8072
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 23198 8072 23204 8084
rect 22888 8044 23204 8072
rect 22888 8032 22894 8044
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 36354 8072 36360 8084
rect 36315 8044 36360 8072
rect 36354 8032 36360 8044
rect 36412 8032 36418 8084
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 8004 10011 8007
rect 10686 8004 10692 8016
rect 9999 7976 10692 8004
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 10686 7964 10692 7976
rect 10744 8004 10750 8016
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 10744 7976 13001 8004
rect 10744 7964 10750 7976
rect 12989 7973 13001 7976
rect 13035 8004 13047 8007
rect 13814 8004 13820 8016
rect 13035 7976 13820 8004
rect 13035 7973 13047 7976
rect 12989 7967 13047 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 21266 7964 21272 8016
rect 21324 8004 21330 8016
rect 21729 8007 21787 8013
rect 21729 8004 21741 8007
rect 21324 7976 21741 8004
rect 21324 7964 21330 7976
rect 21729 7973 21741 7976
rect 21775 8004 21787 8007
rect 21818 8004 21824 8016
rect 21775 7976 21824 8004
rect 21775 7973 21787 7976
rect 21729 7967 21787 7973
rect 21818 7964 21824 7976
rect 21876 7964 21882 8016
rect 22097 8007 22155 8013
rect 22097 7973 22109 8007
rect 22143 8004 22155 8007
rect 23014 8004 23020 8016
rect 22143 7976 23020 8004
rect 22143 7973 22155 7976
rect 22097 7967 22155 7973
rect 23014 7964 23020 7976
rect 23072 7964 23078 8016
rect 23290 8004 23296 8016
rect 23251 7976 23296 8004
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 23658 8004 23664 8016
rect 23619 7976 23664 8004
rect 23658 7964 23664 7976
rect 23716 7964 23722 8016
rect 18322 7936 18328 7948
rect 18283 7908 18328 7936
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 18782 7936 18788 7948
rect 18743 7908 18788 7936
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7936 19211 7939
rect 19426 7936 19432 7948
rect 19199 7908 19432 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 19168 7868 19196 7899
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 19610 7936 19616 7948
rect 19571 7908 19616 7936
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 20530 7896 20536 7948
rect 20588 7936 20594 7948
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 20588 7908 21557 7936
rect 20588 7896 20594 7908
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 21836 7936 21864 7964
rect 23109 7939 23167 7945
rect 23109 7936 23121 7939
rect 21692 7908 21785 7936
rect 21836 7908 23121 7936
rect 21692 7896 21698 7908
rect 23109 7905 23121 7908
rect 23155 7936 23167 7939
rect 23198 7936 23204 7948
rect 23155 7908 23204 7936
rect 23155 7905 23167 7908
rect 23109 7899 23167 7905
rect 23198 7896 23204 7908
rect 23256 7896 23262 7948
rect 18656 7840 19196 7868
rect 18656 7828 18662 7840
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21174 7868 21180 7880
rect 20864 7840 21180 7868
rect 20864 7828 20870 7840
rect 21174 7828 21180 7840
rect 21232 7868 21238 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21232 7840 21373 7868
rect 21232 7828 21238 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 18322 7760 18328 7812
rect 18380 7800 18386 7812
rect 21652 7800 21680 7896
rect 22922 7868 22928 7880
rect 22883 7840 22928 7868
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 18380 7772 21680 7800
rect 18380 7760 18386 7772
rect 20070 7732 20076 7744
rect 20031 7704 20076 7732
rect 20070 7692 20076 7704
rect 20128 7692 20134 7744
rect 21266 7732 21272 7744
rect 21227 7704 21272 7732
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 1104 7642 106812 7664
rect 1104 7590 18982 7642
rect 19034 7590 19046 7642
rect 19098 7590 19110 7642
rect 19162 7590 19174 7642
rect 19226 7590 54982 7642
rect 55034 7590 55046 7642
rect 55098 7590 55110 7642
rect 55162 7590 55174 7642
rect 55226 7590 90982 7642
rect 91034 7590 91046 7642
rect 91098 7590 91110 7642
rect 91162 7590 91174 7642
rect 91226 7590 106812 7642
rect 1104 7568 106812 7590
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 15528 7500 17417 7528
rect 15528 7488 15534 7500
rect 17405 7497 17417 7500
rect 17451 7528 17463 7531
rect 18598 7528 18604 7540
rect 17451 7500 18604 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 19797 7531 19855 7537
rect 19797 7528 19809 7531
rect 18840 7500 19809 7528
rect 18840 7488 18846 7500
rect 19797 7497 19809 7500
rect 19843 7528 19855 7531
rect 20070 7528 20076 7540
rect 19843 7500 20076 7528
rect 19843 7497 19855 7500
rect 19797 7491 19855 7497
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 20625 7531 20683 7537
rect 20625 7528 20637 7531
rect 20588 7500 20637 7528
rect 20588 7488 20594 7500
rect 20625 7497 20637 7500
rect 20671 7528 20683 7531
rect 20993 7531 21051 7537
rect 20993 7528 21005 7531
rect 20671 7500 21005 7528
rect 20671 7497 20683 7500
rect 20625 7491 20683 7497
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 17773 7463 17831 7469
rect 17773 7460 17785 7463
rect 9548 7432 17785 7460
rect 9548 7420 9554 7432
rect 17773 7429 17785 7432
rect 17819 7460 17831 7463
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 17819 7432 18245 7460
rect 17819 7429 17831 7432
rect 17773 7423 17831 7429
rect 18233 7429 18245 7432
rect 18279 7460 18291 7463
rect 18322 7460 18328 7472
rect 18279 7432 18328 7460
rect 18279 7429 18291 7432
rect 18233 7423 18291 7429
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13320 7364 13814 7392
rect 13320 7352 13326 7364
rect 13786 7256 13814 7364
rect 18248 7324 18276 7423
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 19521 7463 19579 7469
rect 19521 7429 19533 7463
rect 19567 7460 19579 7463
rect 19610 7460 19616 7472
rect 19567 7432 19616 7460
rect 19567 7429 19579 7432
rect 19521 7423 19579 7429
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18248 7296 18521 7324
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 20916 7324 20944 7500
rect 20993 7497 21005 7500
rect 21039 7497 21051 7531
rect 20993 7491 21051 7497
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 22189 7531 22247 7537
rect 22189 7528 22201 7531
rect 21692 7500 22201 7528
rect 21692 7488 21698 7500
rect 22189 7497 22201 7500
rect 22235 7497 22247 7531
rect 22189 7491 22247 7497
rect 22830 7488 22836 7540
rect 22888 7528 22894 7540
rect 22925 7531 22983 7537
rect 22925 7528 22937 7531
rect 22888 7500 22937 7528
rect 22888 7488 22894 7500
rect 22925 7497 22937 7500
rect 22971 7497 22983 7531
rect 22925 7491 22983 7497
rect 23198 7488 23204 7540
rect 23256 7528 23262 7540
rect 23293 7531 23351 7537
rect 23293 7528 23305 7531
rect 23256 7500 23305 7528
rect 23256 7488 23262 7500
rect 23293 7497 23305 7500
rect 23339 7497 23351 7531
rect 23293 7491 23351 7497
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 22557 7463 22615 7469
rect 22557 7460 22569 7463
rect 21232 7432 22569 7460
rect 21232 7420 21238 7432
rect 22557 7429 22569 7432
rect 22603 7429 22615 7463
rect 22557 7423 22615 7429
rect 21266 7352 21272 7404
rect 21324 7392 21330 7404
rect 21910 7392 21916 7404
rect 21324 7364 21588 7392
rect 21871 7364 21916 7392
rect 21324 7352 21330 7364
rect 20990 7324 20996 7336
rect 20903 7296 20996 7324
rect 18509 7287 18567 7293
rect 20990 7284 20996 7296
rect 21048 7324 21054 7336
rect 21560 7333 21588 7364
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 21361 7327 21419 7333
rect 21361 7324 21373 7327
rect 21048 7296 21373 7324
rect 21048 7284 21054 7296
rect 21361 7293 21373 7296
rect 21407 7293 21419 7327
rect 21361 7287 21419 7293
rect 21529 7327 21588 7333
rect 21529 7293 21541 7327
rect 21575 7296 21588 7327
rect 21575 7293 21587 7296
rect 21529 7287 21587 7293
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 13786 7228 18429 7256
rect 18417 7225 18429 7228
rect 18463 7256 18475 7259
rect 19702 7256 19708 7268
rect 18463 7228 19708 7256
rect 18463 7225 18475 7228
rect 18417 7219 18475 7225
rect 19702 7216 19708 7228
rect 19760 7216 19766 7268
rect 20349 7259 20407 7265
rect 20349 7225 20361 7259
rect 20395 7256 20407 7259
rect 21174 7256 21180 7268
rect 20395 7228 21180 7256
rect 20395 7225 20407 7228
rect 20349 7219 20407 7225
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 21450 7188 21456 7200
rect 21411 7160 21456 7188
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 1104 7098 106812 7120
rect 1104 7046 36982 7098
rect 37034 7046 37046 7098
rect 37098 7046 37110 7098
rect 37162 7046 37174 7098
rect 37226 7046 72982 7098
rect 73034 7046 73046 7098
rect 73098 7046 73110 7098
rect 73162 7046 73174 7098
rect 73226 7046 106812 7098
rect 1104 7024 106812 7046
rect 18782 6984 18788 6996
rect 18743 6956 18788 6984
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 19702 6944 19708 6996
rect 19760 6984 19766 6996
rect 20625 6987 20683 6993
rect 20625 6984 20637 6987
rect 19760 6956 20637 6984
rect 19760 6944 19766 6956
rect 20625 6953 20637 6956
rect 20671 6984 20683 6987
rect 21450 6984 21456 6996
rect 20671 6956 21456 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 23290 6984 23296 6996
rect 21652 6956 23296 6984
rect 18322 6808 18328 6860
rect 18380 6848 18386 6860
rect 18417 6851 18475 6857
rect 18417 6848 18429 6851
rect 18380 6820 18429 6848
rect 18380 6808 18386 6820
rect 18417 6817 18429 6820
rect 18463 6817 18475 6851
rect 20990 6848 20996 6860
rect 20951 6820 20996 6848
rect 18417 6811 18475 6817
rect 18432 6780 18460 6811
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 21468 6848 21496 6944
rect 21652 6925 21680 6956
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 21637 6919 21695 6925
rect 21637 6885 21649 6919
rect 21683 6885 21695 6919
rect 21637 6879 21695 6885
rect 22922 6848 22928 6860
rect 21468 6820 22928 6848
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 21266 6780 21272 6792
rect 18432 6752 21272 6780
rect 21266 6740 21272 6752
rect 21324 6780 21330 6792
rect 21913 6783 21971 6789
rect 21913 6780 21925 6783
rect 21324 6752 21925 6780
rect 21324 6740 21330 6752
rect 21913 6749 21925 6752
rect 21959 6749 21971 6783
rect 21913 6743 21971 6749
rect 1104 6554 106812 6576
rect 1104 6502 18982 6554
rect 19034 6502 19046 6554
rect 19098 6502 19110 6554
rect 19162 6502 19174 6554
rect 19226 6502 54982 6554
rect 55034 6502 55046 6554
rect 55098 6502 55110 6554
rect 55162 6502 55174 6554
rect 55226 6502 90982 6554
rect 91034 6502 91046 6554
rect 91098 6502 91110 6554
rect 91162 6502 91174 6554
rect 91226 6502 106812 6554
rect 1104 6480 106812 6502
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 18322 6100 18328 6112
rect 18283 6072 18328 6100
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 1104 6010 106812 6032
rect 1104 5958 36982 6010
rect 37034 5958 37046 6010
rect 37098 5958 37110 6010
rect 37162 5958 37174 6010
rect 37226 5958 72982 6010
rect 73034 5958 73046 6010
rect 73098 5958 73110 6010
rect 73162 5958 73174 6010
rect 73226 5958 106812 6010
rect 1104 5936 106812 5958
rect 1104 5466 106812 5488
rect 1104 5414 18982 5466
rect 19034 5414 19046 5466
rect 19098 5414 19110 5466
rect 19162 5414 19174 5466
rect 19226 5414 54982 5466
rect 55034 5414 55046 5466
rect 55098 5414 55110 5466
rect 55162 5414 55174 5466
rect 55226 5414 90982 5466
rect 91034 5414 91046 5466
rect 91098 5414 91110 5466
rect 91162 5414 91174 5466
rect 91226 5414 106812 5466
rect 1104 5392 106812 5414
rect 1104 4922 106812 4944
rect 1104 4870 36982 4922
rect 37034 4870 37046 4922
rect 37098 4870 37110 4922
rect 37162 4870 37174 4922
rect 37226 4870 72982 4922
rect 73034 4870 73046 4922
rect 73098 4870 73110 4922
rect 73162 4870 73174 4922
rect 73226 4870 106812 4922
rect 1104 4848 106812 4870
rect 1104 4378 106812 4400
rect 1104 4326 18982 4378
rect 19034 4326 19046 4378
rect 19098 4326 19110 4378
rect 19162 4326 19174 4378
rect 19226 4326 54982 4378
rect 55034 4326 55046 4378
rect 55098 4326 55110 4378
rect 55162 4326 55174 4378
rect 55226 4326 90982 4378
rect 91034 4326 91046 4378
rect 91098 4326 91110 4378
rect 91162 4326 91174 4378
rect 91226 4326 106812 4378
rect 1104 4304 106812 4326
rect 1104 3834 106812 3856
rect 1104 3782 36982 3834
rect 37034 3782 37046 3834
rect 37098 3782 37110 3834
rect 37162 3782 37174 3834
rect 37226 3782 72982 3834
rect 73034 3782 73046 3834
rect 73098 3782 73110 3834
rect 73162 3782 73174 3834
rect 73226 3782 106812 3834
rect 1104 3760 106812 3782
rect 1104 3290 106812 3312
rect 1104 3238 18982 3290
rect 19034 3238 19046 3290
rect 19098 3238 19110 3290
rect 19162 3238 19174 3290
rect 19226 3238 54982 3290
rect 55034 3238 55046 3290
rect 55098 3238 55110 3290
rect 55162 3238 55174 3290
rect 55226 3238 90982 3290
rect 91034 3238 91046 3290
rect 91098 3238 91110 3290
rect 91162 3238 91174 3290
rect 91226 3238 106812 3290
rect 1104 3216 106812 3238
rect 1104 2746 106812 2768
rect 1104 2694 36982 2746
rect 37034 2694 37046 2746
rect 37098 2694 37110 2746
rect 37162 2694 37174 2746
rect 37226 2694 72982 2746
rect 73034 2694 73046 2746
rect 73098 2694 73110 2746
rect 73162 2694 73174 2746
rect 73226 2694 106812 2746
rect 1104 2672 106812 2694
rect 1104 2202 106812 2224
rect 1104 2150 18982 2202
rect 19034 2150 19046 2202
rect 19098 2150 19110 2202
rect 19162 2150 19174 2202
rect 19226 2150 54982 2202
rect 55034 2150 55046 2202
rect 55098 2150 55110 2202
rect 55162 2150 55174 2202
rect 55226 2150 90982 2202
rect 91034 2150 91046 2202
rect 91098 2150 91110 2202
rect 91162 2150 91174 2202
rect 91226 2150 106812 2202
rect 1104 2128 106812 2150
rect 71866 76 71872 128
rect 71924 116 71930 128
rect 74166 116 74172 128
rect 71924 88 74172 116
rect 71924 76 71930 88
rect 74166 76 74172 88
rect 74224 76 74230 128
<< via1 >>
rect 36982 11398 37034 11450
rect 37046 11398 37098 11450
rect 37110 11398 37162 11450
rect 37174 11398 37226 11450
rect 72982 11398 73034 11450
rect 73046 11398 73098 11450
rect 73110 11398 73162 11450
rect 73174 11398 73226 11450
rect 18982 10854 19034 10906
rect 19046 10854 19098 10906
rect 19110 10854 19162 10906
rect 19174 10854 19226 10906
rect 54982 10854 55034 10906
rect 55046 10854 55098 10906
rect 55110 10854 55162 10906
rect 55174 10854 55226 10906
rect 90982 10854 91034 10906
rect 91046 10854 91098 10906
rect 91110 10854 91162 10906
rect 91174 10854 91226 10906
rect 36982 10310 37034 10362
rect 37046 10310 37098 10362
rect 37110 10310 37162 10362
rect 37174 10310 37226 10362
rect 72982 10310 73034 10362
rect 73046 10310 73098 10362
rect 73110 10310 73162 10362
rect 73174 10310 73226 10362
rect 12900 10251 12952 10260
rect 12900 10217 12909 10251
rect 12909 10217 12943 10251
rect 12943 10217 12952 10251
rect 12900 10208 12952 10217
rect 26700 10251 26752 10260
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 39396 10251 39448 10260
rect 39396 10217 39405 10251
rect 39405 10217 39439 10251
rect 39439 10217 39448 10251
rect 39396 10208 39448 10217
rect 66352 10251 66404 10260
rect 66352 10217 66361 10251
rect 66361 10217 66395 10251
rect 66395 10217 66404 10251
rect 66352 10208 66404 10217
rect 79876 10251 79928 10260
rect 79876 10217 79885 10251
rect 79885 10217 79919 10251
rect 79919 10217 79928 10251
rect 79876 10208 79928 10217
rect 16764 10140 16816 10192
rect 10416 10115 10468 10124
rect 10416 10081 10425 10115
rect 10425 10081 10459 10115
rect 10459 10081 10468 10115
rect 10416 10072 10468 10081
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 21824 10115 21876 10124
rect 21824 10081 21833 10115
rect 21833 10081 21867 10115
rect 21867 10081 21876 10115
rect 21824 10072 21876 10081
rect 26608 10072 26660 10124
rect 39304 10072 39356 10124
rect 49056 10072 49108 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 10876 10004 10928 10056
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 35072 10004 35124 10056
rect 35440 10004 35492 10056
rect 49332 10004 49384 10056
rect 52368 10072 52420 10124
rect 52736 10115 52788 10124
rect 52736 10081 52745 10115
rect 52745 10081 52779 10115
rect 52779 10081 52788 10115
rect 52736 10072 52788 10081
rect 61568 10072 61620 10124
rect 57336 10004 57388 10056
rect 66260 10072 66312 10124
rect 79692 10115 79744 10124
rect 79692 10081 79701 10115
rect 79701 10081 79735 10115
rect 79735 10081 79744 10115
rect 79692 10072 79744 10081
rect 87880 10072 87932 10124
rect 70768 10004 70820 10056
rect 75184 10004 75236 10056
rect 75460 10004 75512 10056
rect 89076 10004 89128 10056
rect 61844 9936 61896 9988
rect 2044 9911 2096 9920
rect 2044 9877 2053 9911
rect 2053 9877 2087 9911
rect 2087 9877 2096 9911
rect 2044 9868 2096 9877
rect 23388 9868 23440 9920
rect 36176 9911 36228 9920
rect 36176 9877 36185 9911
rect 36185 9877 36219 9911
rect 36219 9877 36228 9911
rect 36176 9868 36228 9877
rect 61476 9868 61528 9920
rect 78588 9868 78640 9920
rect 88708 9911 88760 9920
rect 88708 9877 88717 9911
rect 88717 9877 88751 9911
rect 88751 9877 88760 9911
rect 88708 9868 88760 9877
rect 18982 9766 19034 9818
rect 19046 9766 19098 9818
rect 19110 9766 19162 9818
rect 19174 9766 19226 9818
rect 54982 9766 55034 9818
rect 55046 9766 55098 9818
rect 55110 9766 55162 9818
rect 55174 9766 55226 9818
rect 90982 9766 91034 9818
rect 91046 9766 91098 9818
rect 91110 9766 91162 9818
rect 91174 9766 91226 9818
rect 1584 9664 1636 9716
rect 2320 9664 2372 9716
rect 10416 9707 10468 9716
rect 10416 9673 10425 9707
rect 10425 9673 10459 9707
rect 10459 9673 10468 9707
rect 10416 9664 10468 9673
rect 21824 9707 21876 9716
rect 21824 9673 21833 9707
rect 21833 9673 21867 9707
rect 21867 9673 21876 9707
rect 21824 9664 21876 9673
rect 49056 9707 49108 9716
rect 49056 9673 49065 9707
rect 49065 9673 49099 9707
rect 49099 9673 49108 9707
rect 49056 9664 49108 9673
rect 52736 9707 52788 9716
rect 52736 9673 52745 9707
rect 52745 9673 52779 9707
rect 52779 9673 52788 9707
rect 52736 9664 52788 9673
rect 61568 9707 61620 9716
rect 61568 9673 61577 9707
rect 61577 9673 61611 9707
rect 61611 9673 61620 9707
rect 61568 9664 61620 9673
rect 89076 9707 89128 9716
rect 89076 9673 89085 9707
rect 89085 9673 89119 9707
rect 89119 9673 89128 9707
rect 89076 9664 89128 9673
rect 1400 9596 1452 9648
rect 3332 9596 3384 9648
rect 22008 9596 22060 9648
rect 23388 9596 23440 9648
rect 26608 9596 26660 9648
rect 35164 9639 35216 9648
rect 35164 9605 35173 9639
rect 35173 9605 35207 9639
rect 35207 9605 35216 9639
rect 35164 9596 35216 9605
rect 75184 9639 75236 9648
rect 75184 9605 75193 9639
rect 75193 9605 75227 9639
rect 75227 9605 75236 9639
rect 75184 9596 75236 9605
rect 61844 9571 61896 9580
rect 61844 9537 61853 9571
rect 61853 9537 61887 9571
rect 61887 9537 61896 9571
rect 61844 9528 61896 9537
rect 19524 9460 19576 9512
rect 36176 9503 36228 9512
rect 36176 9469 36185 9503
rect 36185 9469 36219 9503
rect 36219 9469 36228 9503
rect 36176 9460 36228 9469
rect 39948 9460 40000 9512
rect 88708 9460 88760 9512
rect 2044 9435 2096 9444
rect 2044 9401 2053 9435
rect 2053 9401 2087 9435
rect 2087 9401 2096 9435
rect 2044 9392 2096 9401
rect 6460 9392 6512 9444
rect 1676 9324 1728 9376
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 19800 9367 19852 9376
rect 19800 9333 19809 9367
rect 19809 9333 19843 9367
rect 19843 9333 19852 9367
rect 19800 9324 19852 9333
rect 26608 9367 26660 9376
rect 26608 9333 26617 9367
rect 26617 9333 26651 9367
rect 26651 9333 26660 9367
rect 26608 9324 26660 9333
rect 35440 9367 35492 9376
rect 35440 9333 35449 9367
rect 35449 9333 35483 9367
rect 35483 9333 35492 9367
rect 35440 9324 35492 9333
rect 36084 9367 36136 9376
rect 36084 9333 36093 9367
rect 36093 9333 36127 9367
rect 36127 9333 36136 9367
rect 36084 9324 36136 9333
rect 39304 9367 39356 9376
rect 39304 9333 39313 9367
rect 39313 9333 39347 9367
rect 39347 9333 39356 9367
rect 39304 9324 39356 9333
rect 49332 9367 49384 9376
rect 49332 9333 49341 9367
rect 49341 9333 49375 9367
rect 49375 9333 49384 9367
rect 49332 9324 49384 9333
rect 66260 9367 66312 9376
rect 66260 9333 66269 9367
rect 66269 9333 66303 9367
rect 66303 9333 66312 9367
rect 66260 9324 66312 9333
rect 75460 9367 75512 9376
rect 75460 9333 75469 9367
rect 75469 9333 75503 9367
rect 75503 9333 75512 9367
rect 75460 9324 75512 9333
rect 78588 9324 78640 9376
rect 79692 9324 79744 9376
rect 87880 9367 87932 9376
rect 87880 9333 87889 9367
rect 87889 9333 87923 9367
rect 87923 9333 87932 9367
rect 87880 9324 87932 9333
rect 88248 9367 88300 9376
rect 88248 9333 88257 9367
rect 88257 9333 88291 9367
rect 88291 9333 88300 9367
rect 88248 9324 88300 9333
rect 88708 9367 88760 9376
rect 88708 9333 88717 9367
rect 88717 9333 88751 9367
rect 88751 9333 88760 9367
rect 88708 9324 88760 9333
rect 36982 9222 37034 9274
rect 37046 9222 37098 9274
rect 37110 9222 37162 9274
rect 37174 9222 37226 9274
rect 72982 9222 73034 9274
rect 73046 9222 73098 9274
rect 73110 9222 73162 9274
rect 73174 9222 73226 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 10876 9120 10928 9172
rect 21824 9163 21876 9172
rect 21824 9129 21833 9163
rect 21833 9129 21867 9163
rect 21867 9129 21876 9163
rect 21824 9120 21876 9129
rect 35440 9120 35492 9172
rect 49332 9120 49384 9172
rect 1492 9052 1544 9104
rect 11428 9052 11480 9104
rect 21916 9095 21968 9104
rect 21916 9061 21925 9095
rect 21925 9061 21959 9095
rect 21959 9061 21968 9095
rect 21916 9052 21968 9061
rect 22100 9052 22152 9104
rect 23296 9052 23348 9104
rect 32128 9052 32180 9104
rect 36084 9052 36136 9104
rect 39764 8984 39816 9036
rect 2044 8916 2096 8968
rect 10876 8959 10928 8968
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 32496 8916 32548 8968
rect 35440 8916 35492 8968
rect 37648 8916 37700 8968
rect 9956 8823 10008 8832
rect 9956 8789 9965 8823
rect 9965 8789 9999 8823
rect 9999 8789 10008 8823
rect 9956 8780 10008 8789
rect 13268 8780 13320 8832
rect 19524 8823 19576 8832
rect 19524 8789 19533 8823
rect 19533 8789 19567 8823
rect 19567 8789 19576 8823
rect 19524 8780 19576 8789
rect 19708 8780 19760 8832
rect 18982 8678 19034 8730
rect 19046 8678 19098 8730
rect 19110 8678 19162 8730
rect 19174 8678 19226 8730
rect 54982 8678 55034 8730
rect 55046 8678 55098 8730
rect 55110 8678 55162 8730
rect 55174 8678 55226 8730
rect 90982 8678 91034 8730
rect 91046 8678 91098 8730
rect 91110 8678 91162 8730
rect 91174 8678 91226 8730
rect 1492 8576 1544 8628
rect 11428 8619 11480 8628
rect 11428 8585 11437 8619
rect 11437 8585 11471 8619
rect 11471 8585 11480 8619
rect 11428 8576 11480 8585
rect 19800 8576 19852 8628
rect 21916 8576 21968 8628
rect 32496 8619 32548 8628
rect 32496 8585 32505 8619
rect 32505 8585 32539 8619
rect 32539 8585 32548 8619
rect 32496 8576 32548 8585
rect 9496 8440 9548 8492
rect 2044 8279 2096 8288
rect 2044 8245 2053 8279
rect 2053 8245 2087 8279
rect 2087 8245 2096 8279
rect 9128 8279 9180 8288
rect 2044 8236 2096 8245
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 9496 8279 9548 8288
rect 9496 8245 9505 8279
rect 9505 8245 9539 8279
rect 9539 8245 9548 8279
rect 9496 8236 9548 8245
rect 9956 8372 10008 8424
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 10784 8372 10836 8424
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 18788 8440 18840 8492
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 23204 8508 23256 8560
rect 19432 8440 19484 8492
rect 19708 8372 19760 8424
rect 20076 8372 20128 8424
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 22100 8440 22152 8492
rect 35440 8483 35492 8492
rect 21272 8415 21324 8424
rect 20536 8304 20588 8356
rect 13084 8279 13136 8288
rect 13084 8245 13093 8279
rect 13093 8245 13127 8279
rect 13127 8245 13136 8279
rect 13084 8236 13136 8245
rect 13820 8236 13872 8288
rect 15476 8279 15528 8288
rect 15476 8245 15485 8279
rect 15485 8245 15519 8279
rect 15519 8245 15528 8279
rect 15476 8236 15528 8245
rect 19616 8236 19668 8288
rect 21272 8381 21281 8415
rect 21281 8381 21315 8415
rect 21315 8381 21324 8415
rect 21272 8372 21324 8381
rect 21640 8279 21692 8288
rect 21640 8245 21649 8279
rect 21649 8245 21683 8279
rect 21683 8245 21692 8279
rect 21640 8236 21692 8245
rect 21824 8236 21876 8288
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 36360 8415 36412 8424
rect 36360 8381 36369 8415
rect 36369 8381 36403 8415
rect 36403 8381 36412 8415
rect 36360 8372 36412 8381
rect 40040 8372 40092 8424
rect 23296 8236 23348 8288
rect 32128 8279 32180 8288
rect 32128 8245 32137 8279
rect 32137 8245 32171 8279
rect 32171 8245 32180 8279
rect 32128 8236 32180 8245
rect 36084 8236 36136 8288
rect 36820 8304 36872 8356
rect 37648 8304 37700 8356
rect 36982 8134 37034 8186
rect 37046 8134 37098 8186
rect 37110 8134 37162 8186
rect 37174 8134 37226 8186
rect 72982 8134 73034 8186
rect 73046 8134 73098 8186
rect 73110 8134 73162 8186
rect 73174 8134 73226 8186
rect 10876 8032 10928 8084
rect 13084 8032 13136 8084
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 22836 8032 22888 8084
rect 23204 8075 23256 8084
rect 23204 8041 23213 8075
rect 23213 8041 23247 8075
rect 23247 8041 23256 8075
rect 23204 8032 23256 8041
rect 36360 8075 36412 8084
rect 36360 8041 36369 8075
rect 36369 8041 36403 8075
rect 36403 8041 36412 8075
rect 36360 8032 36412 8041
rect 10692 7964 10744 8016
rect 13820 7964 13872 8016
rect 21272 7964 21324 8016
rect 21824 7964 21876 8016
rect 23020 7964 23072 8016
rect 23296 8007 23348 8016
rect 23296 7973 23305 8007
rect 23305 7973 23339 8007
rect 23339 7973 23348 8007
rect 23296 7964 23348 7973
rect 23664 8007 23716 8016
rect 23664 7973 23673 8007
rect 23673 7973 23707 8007
rect 23707 7973 23716 8007
rect 23664 7964 23716 7973
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 18788 7939 18840 7948
rect 18788 7905 18797 7939
rect 18797 7905 18831 7939
rect 18831 7905 18840 7939
rect 18788 7896 18840 7905
rect 18604 7828 18656 7880
rect 19432 7896 19484 7948
rect 19616 7939 19668 7948
rect 19616 7905 19625 7939
rect 19625 7905 19659 7939
rect 19659 7905 19668 7939
rect 19616 7896 19668 7905
rect 20536 7896 20588 7948
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 23204 7896 23256 7948
rect 20812 7828 20864 7880
rect 21180 7828 21232 7880
rect 18328 7760 18380 7812
rect 22928 7871 22980 7880
rect 22928 7837 22937 7871
rect 22937 7837 22971 7871
rect 22971 7837 22980 7871
rect 22928 7828 22980 7837
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 18982 7590 19034 7642
rect 19046 7590 19098 7642
rect 19110 7590 19162 7642
rect 19174 7590 19226 7642
rect 54982 7590 55034 7642
rect 55046 7590 55098 7642
rect 55110 7590 55162 7642
rect 55174 7590 55226 7642
rect 90982 7590 91034 7642
rect 91046 7590 91098 7642
rect 91110 7590 91162 7642
rect 91174 7590 91226 7642
rect 15476 7488 15528 7540
rect 18604 7488 18656 7540
rect 18788 7488 18840 7540
rect 20076 7488 20128 7540
rect 20536 7488 20588 7540
rect 9496 7420 9548 7472
rect 13268 7352 13320 7404
rect 18328 7420 18380 7472
rect 19616 7420 19668 7472
rect 21640 7488 21692 7540
rect 22836 7488 22888 7540
rect 23204 7488 23256 7540
rect 21180 7420 21232 7472
rect 21272 7352 21324 7404
rect 21916 7395 21968 7404
rect 20996 7284 21048 7336
rect 21916 7361 21925 7395
rect 21925 7361 21959 7395
rect 21959 7361 21968 7395
rect 21916 7352 21968 7361
rect 19708 7216 19760 7268
rect 21180 7259 21232 7268
rect 21180 7225 21189 7259
rect 21189 7225 21223 7259
rect 21223 7225 21232 7259
rect 21180 7216 21232 7225
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 36982 7046 37034 7098
rect 37046 7046 37098 7098
rect 37110 7046 37162 7098
rect 37174 7046 37226 7098
rect 72982 7046 73034 7098
rect 73046 7046 73098 7098
rect 73110 7046 73162 7098
rect 73174 7046 73226 7098
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 19708 6944 19760 6996
rect 21456 6944 21508 6996
rect 23296 6987 23348 6996
rect 18328 6808 18380 6860
rect 20996 6851 21048 6860
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 23296 6953 23305 6987
rect 23305 6953 23339 6987
rect 23339 6953 23348 6987
rect 23296 6944 23348 6953
rect 22928 6851 22980 6860
rect 22928 6817 22937 6851
rect 22937 6817 22971 6851
rect 22971 6817 22980 6851
rect 22928 6808 22980 6817
rect 21272 6740 21324 6792
rect 18982 6502 19034 6554
rect 19046 6502 19098 6554
rect 19110 6502 19162 6554
rect 19174 6502 19226 6554
rect 54982 6502 55034 6554
rect 55046 6502 55098 6554
rect 55110 6502 55162 6554
rect 55174 6502 55226 6554
rect 90982 6502 91034 6554
rect 91046 6502 91098 6554
rect 91110 6502 91162 6554
rect 91174 6502 91226 6554
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 18328 6103 18380 6112
rect 18328 6069 18337 6103
rect 18337 6069 18371 6103
rect 18371 6069 18380 6103
rect 18328 6060 18380 6069
rect 36982 5958 37034 6010
rect 37046 5958 37098 6010
rect 37110 5958 37162 6010
rect 37174 5958 37226 6010
rect 72982 5958 73034 6010
rect 73046 5958 73098 6010
rect 73110 5958 73162 6010
rect 73174 5958 73226 6010
rect 18982 5414 19034 5466
rect 19046 5414 19098 5466
rect 19110 5414 19162 5466
rect 19174 5414 19226 5466
rect 54982 5414 55034 5466
rect 55046 5414 55098 5466
rect 55110 5414 55162 5466
rect 55174 5414 55226 5466
rect 90982 5414 91034 5466
rect 91046 5414 91098 5466
rect 91110 5414 91162 5466
rect 91174 5414 91226 5466
rect 36982 4870 37034 4922
rect 37046 4870 37098 4922
rect 37110 4870 37162 4922
rect 37174 4870 37226 4922
rect 72982 4870 73034 4922
rect 73046 4870 73098 4922
rect 73110 4870 73162 4922
rect 73174 4870 73226 4922
rect 18982 4326 19034 4378
rect 19046 4326 19098 4378
rect 19110 4326 19162 4378
rect 19174 4326 19226 4378
rect 54982 4326 55034 4378
rect 55046 4326 55098 4378
rect 55110 4326 55162 4378
rect 55174 4326 55226 4378
rect 90982 4326 91034 4378
rect 91046 4326 91098 4378
rect 91110 4326 91162 4378
rect 91174 4326 91226 4378
rect 36982 3782 37034 3834
rect 37046 3782 37098 3834
rect 37110 3782 37162 3834
rect 37174 3782 37226 3834
rect 72982 3782 73034 3834
rect 73046 3782 73098 3834
rect 73110 3782 73162 3834
rect 73174 3782 73226 3834
rect 18982 3238 19034 3290
rect 19046 3238 19098 3290
rect 19110 3238 19162 3290
rect 19174 3238 19226 3290
rect 54982 3238 55034 3290
rect 55046 3238 55098 3290
rect 55110 3238 55162 3290
rect 55174 3238 55226 3290
rect 90982 3238 91034 3290
rect 91046 3238 91098 3290
rect 91110 3238 91162 3290
rect 91174 3238 91226 3290
rect 36982 2694 37034 2746
rect 37046 2694 37098 2746
rect 37110 2694 37162 2746
rect 37174 2694 37226 2746
rect 72982 2694 73034 2746
rect 73046 2694 73098 2746
rect 73110 2694 73162 2746
rect 73174 2694 73226 2746
rect 18982 2150 19034 2202
rect 19046 2150 19098 2202
rect 19110 2150 19162 2202
rect 19174 2150 19226 2202
rect 54982 2150 55034 2202
rect 55046 2150 55098 2202
rect 55110 2150 55162 2202
rect 55174 2150 55226 2202
rect 90982 2150 91034 2202
rect 91046 2150 91098 2202
rect 91110 2150 91162 2202
rect 91174 2150 91226 2202
rect 71872 76 71924 128
rect 74172 76 74224 128
<< metal2 >>
rect 3330 13520 3386 14000
rect 10046 13520 10102 14000
rect 16762 13520 16818 14000
rect 23570 13520 23626 14000
rect 30286 13520 30342 14000
rect 37002 13520 37058 14000
rect 43810 13520 43866 14000
rect 50526 13520 50582 14000
rect 57334 13520 57390 14000
rect 64050 13520 64106 14000
rect 70766 13520 70822 14000
rect 77574 13520 77630 14000
rect 84290 13520 84346 14000
rect 91006 13546 91062 14000
rect 90744 13520 91062 13546
rect 97814 13520 97870 14000
rect 104530 13520 104586 14000
rect 1490 12200 1546 12209
rect 1490 12135 1546 12144
rect 110 10432 166 10441
rect 110 10367 166 10376
rect 124 8945 152 10367
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9654 1440 9998
rect 1400 9648 1452 9654
rect 1400 9590 1452 9596
rect 1504 9217 1532 12135
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9722 1624 9998
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1688 9382 1716 10911
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9450 2084 9862
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1490 9208 1546 9217
rect 2332 9178 2360 9658
rect 3344 9654 3372 13520
rect 10060 10985 10088 13520
rect 10046 10976 10102 10985
rect 10046 10911 10102 10920
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12912 10169 12940 10202
rect 16776 10198 16804 13520
rect 21822 10976 21878 10985
rect 18956 10908 19252 10928
rect 21822 10911 21878 10920
rect 19012 10906 19036 10908
rect 19092 10906 19116 10908
rect 19172 10906 19196 10908
rect 19034 10854 19036 10906
rect 19098 10854 19110 10906
rect 19172 10854 19174 10906
rect 19012 10852 19036 10854
rect 19092 10852 19116 10854
rect 19172 10852 19196 10854
rect 18956 10832 19252 10852
rect 16764 10192 16816 10198
rect 12898 10160 12954 10169
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 12716 10124 12768 10130
rect 16764 10134 16816 10140
rect 21836 10130 21864 10911
rect 12898 10095 12954 10104
rect 21824 10124 21876 10130
rect 12716 10066 12768 10072
rect 21824 10066 21876 10072
rect 10428 9722 10456 10066
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 1490 9143 1546 9152
rect 2320 9172 2372 9178
rect 1504 9110 1532 9143
rect 2320 9114 2372 9120
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 110 8936 166 8945
rect 110 8871 166 8880
rect 1504 8634 1532 9046
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 110 8392 166 8401
rect 110 8327 166 8336
rect 124 8129 152 8327
rect 2056 8294 2084 8910
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 110 8120 166 8129
rect 110 8055 166 8064
rect 6472 82 6500 9386
rect 10888 9382 10916 9998
rect 12728 9382 12756 10066
rect 18956 9820 19252 9840
rect 19012 9818 19036 9820
rect 19092 9818 19116 9820
rect 19172 9818 19196 9820
rect 19034 9766 19036 9818
rect 19098 9766 19110 9818
rect 19172 9766 19174 9818
rect 19012 9764 19036 9766
rect 19092 9764 19116 9766
rect 19172 9764 19196 9766
rect 18956 9744 19252 9764
rect 21836 9722 21864 10066
rect 22008 10056 22060 10062
rect 23584 10033 23612 13520
rect 30300 10985 30328 13520
rect 37016 11914 37044 13520
rect 36832 11886 37044 11914
rect 30286 10976 30342 10985
rect 30286 10911 30342 10920
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26712 10169 26740 10202
rect 36832 10169 36860 11886
rect 36956 11452 37252 11472
rect 37012 11450 37036 11452
rect 37092 11450 37116 11452
rect 37172 11450 37196 11452
rect 37034 11398 37036 11450
rect 37098 11398 37110 11450
rect 37172 11398 37174 11450
rect 37012 11396 37036 11398
rect 37092 11396 37116 11398
rect 37172 11396 37196 11398
rect 36956 11376 37252 11396
rect 36956 10364 37252 10384
rect 37012 10362 37036 10364
rect 37092 10362 37116 10364
rect 37172 10362 37196 10364
rect 37034 10310 37036 10362
rect 37098 10310 37110 10362
rect 37172 10310 37174 10362
rect 37012 10308 37036 10310
rect 37092 10308 37116 10310
rect 37172 10308 37196 10310
rect 36956 10288 37252 10308
rect 39396 10260 39448 10266
rect 39396 10202 39448 10208
rect 39408 10169 39436 10202
rect 26698 10160 26754 10169
rect 26608 10124 26660 10130
rect 26698 10095 26754 10104
rect 36818 10160 36874 10169
rect 39394 10160 39450 10169
rect 36818 10095 36874 10104
rect 39304 10124 39356 10130
rect 26608 10066 26660 10072
rect 39394 10095 39450 10104
rect 39304 10066 39356 10072
rect 22008 9998 22060 10004
rect 23570 10024 23626 10033
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 22020 9654 22048 9998
rect 23570 9959 23626 9968
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23400 9654 23428 9862
rect 26620 9654 26648 10066
rect 35072 10056 35124 10062
rect 35440 10056 35492 10062
rect 35124 10016 35204 10044
rect 35072 9998 35124 10004
rect 35176 9761 35204 10016
rect 35440 9998 35492 10004
rect 35162 9752 35218 9761
rect 35162 9687 35218 9696
rect 35176 9654 35204 9687
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 35164 9648 35216 9654
rect 35164 9590 35216 9596
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 10888 9178 10916 9318
rect 11426 9208 11482 9217
rect 10876 9172 10928 9178
rect 11426 9143 11482 9152
rect 10876 9114 10928 9120
rect 11440 9110 11468 9143
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9126 8392 9182 8401
rect 9126 8327 9182 8336
rect 9140 8294 9168 8327
rect 9508 8294 9536 8434
rect 9968 8430 9996 8774
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9508 7478 9536 8230
rect 10704 8022 10732 8366
rect 10796 8265 10824 8366
rect 10782 8256 10838 8265
rect 10782 8191 10838 8200
rect 10888 8090 10916 8910
rect 11440 8634 11468 9046
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9508 6361 9536 7414
rect 9494 6352 9550 6361
rect 9494 6287 9550 6296
rect 12728 2825 12756 9318
rect 15290 8936 15346 8945
rect 15290 8871 15346 8880
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8430 13308 8774
rect 15304 8430 15332 8871
rect 19536 8838 19564 9454
rect 26620 9382 26648 9590
rect 35452 9382 35480 9998
rect 36176 9920 36228 9926
rect 36176 9862 36228 9868
rect 36188 9518 36216 9862
rect 36176 9512 36228 9518
rect 36176 9454 36228 9460
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 26608 9376 26660 9382
rect 26608 9318 26660 9324
rect 35440 9376 35492 9382
rect 35440 9318 35492 9324
rect 36084 9376 36136 9382
rect 36084 9318 36136 9324
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 18956 8732 19252 8752
rect 19012 8730 19036 8732
rect 19092 8730 19116 8732
rect 19172 8730 19196 8732
rect 19034 8678 19036 8730
rect 19098 8678 19110 8730
rect 19172 8678 19174 8730
rect 19012 8676 19036 8678
rect 19092 8676 19116 8678
rect 19172 8676 19196 8678
rect 18956 8656 19252 8676
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 8090 13124 8230
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13280 7410 13308 8366
rect 13832 8294 13860 8366
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 13832 8022 13860 8230
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 15488 7546 15516 8230
rect 18800 7954 18828 8434
rect 19444 7954 19472 8434
rect 19536 8090 19564 8774
rect 19720 8430 19748 8774
rect 19812 8634 19840 9318
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19628 7954 19656 8230
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 18340 7818 18368 7890
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 18340 7478 18368 7754
rect 18616 7546 18644 7822
rect 18800 7546 18828 7890
rect 18956 7644 19252 7664
rect 19012 7642 19036 7644
rect 19092 7642 19116 7644
rect 19172 7642 19196 7644
rect 19034 7590 19036 7642
rect 19098 7590 19110 7642
rect 19172 7590 19174 7642
rect 19012 7588 19036 7590
rect 19092 7588 19116 7590
rect 19172 7588 19196 7590
rect 18956 7568 19252 7588
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 18800 7002 18828 7482
rect 19628 7478 19656 7890
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19720 7274 19748 8366
rect 19812 8129 19840 8570
rect 21270 8528 21326 8537
rect 21270 8463 21326 8472
rect 21284 8430 21312 8463
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 19798 8120 19854 8129
rect 19798 8055 19854 8064
rect 20088 7750 20116 8366
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20548 7954 20576 8298
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 20088 7546 20116 7686
rect 20548 7546 20576 7890
rect 20824 7886 20852 8366
rect 21652 8294 21680 8910
rect 21836 8294 21864 9114
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 22100 9104 22152 9110
rect 23296 9104 23348 9110
rect 22100 9046 22152 9052
rect 23202 9072 23258 9081
rect 21928 8634 21956 9046
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 22112 8498 22140 9046
rect 23258 9052 23296 9058
rect 23258 9046 23348 9052
rect 23258 9030 23336 9046
rect 23202 9007 23258 9016
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21914 8392 21970 8401
rect 21914 8327 21970 8336
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 21192 7478 21220 7822
rect 21284 7750 21312 7958
rect 21652 7954 21680 8230
rect 21836 8022 21864 8230
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19720 7002 19748 7210
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 21008 6866 21036 7278
rect 21192 7274 21220 7414
rect 21284 7410 21312 7686
rect 21652 7546 21680 7890
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21928 7410 21956 8327
rect 23216 8090 23244 8502
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23662 8256 23718 8265
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 22848 7546 22876 8026
rect 23308 8022 23336 8230
rect 23662 8191 23718 8200
rect 23676 8022 23704 8191
rect 23020 8016 23072 8022
rect 23296 8016 23348 8022
rect 23072 7993 23152 8004
rect 23072 7984 23166 7993
rect 23072 7976 23110 7984
rect 23020 7958 23072 7964
rect 23296 7958 23348 7964
rect 23664 8016 23716 8022
rect 23664 7958 23716 7964
rect 23110 7919 23166 7928
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 18340 6118 18368 6802
rect 18956 6556 19252 6576
rect 19012 6554 19036 6556
rect 19092 6554 19116 6556
rect 19172 6554 19196 6556
rect 19034 6502 19036 6554
rect 19098 6502 19110 6554
rect 19172 6502 19174 6554
rect 19012 6500 19036 6502
rect 19092 6500 19116 6502
rect 19172 6500 19196 6502
rect 18956 6480 19252 6500
rect 21008 6458 21036 6802
rect 21284 6798 21312 7346
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 7002 21496 7142
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 22940 6866 22968 7822
rect 23216 7546 23244 7890
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23308 7002 23336 7958
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 12714 2816 12770 2825
rect 12714 2751 12770 2760
rect 18340 1329 18368 6054
rect 18956 5468 19252 5488
rect 19012 5466 19036 5468
rect 19092 5466 19116 5468
rect 19172 5466 19196 5468
rect 19034 5414 19036 5466
rect 19098 5414 19110 5466
rect 19172 5414 19174 5466
rect 19012 5412 19036 5414
rect 19092 5412 19116 5414
rect 19172 5412 19196 5414
rect 18956 5392 19252 5412
rect 26620 4865 26648 9318
rect 35452 9178 35480 9318
rect 35440 9172 35492 9178
rect 35440 9114 35492 9120
rect 36096 9110 36124 9318
rect 32128 9104 32180 9110
rect 32128 9046 32180 9052
rect 36084 9104 36136 9110
rect 36188 9081 36216 9454
rect 39316 9382 39344 10066
rect 43824 9761 43852 13520
rect 50540 10169 50568 13520
rect 54956 10908 55252 10928
rect 55012 10906 55036 10908
rect 55092 10906 55116 10908
rect 55172 10906 55196 10908
rect 55034 10854 55036 10906
rect 55098 10854 55110 10906
rect 55172 10854 55174 10906
rect 55012 10852 55036 10854
rect 55092 10852 55116 10854
rect 55172 10852 55196 10854
rect 54956 10832 55252 10852
rect 50526 10160 50582 10169
rect 49056 10124 49108 10130
rect 50526 10095 50582 10104
rect 52368 10124 52420 10130
rect 49056 10066 49108 10072
rect 52368 10066 52420 10072
rect 52736 10124 52788 10130
rect 52736 10066 52788 10072
rect 43810 9752 43866 9761
rect 49068 9722 49096 10066
rect 49332 10056 49384 10062
rect 49332 9998 49384 10004
rect 43810 9687 43866 9696
rect 49056 9716 49108 9722
rect 49056 9658 49108 9664
rect 39948 9512 40000 9518
rect 39948 9454 40000 9460
rect 39304 9376 39356 9382
rect 39960 9353 39988 9454
rect 49344 9382 49372 9998
rect 49332 9376 49384 9382
rect 39304 9318 39356 9324
rect 39946 9344 40002 9353
rect 36956 9276 37252 9296
rect 37012 9274 37036 9276
rect 37092 9274 37116 9276
rect 37172 9274 37196 9276
rect 37034 9222 37036 9274
rect 37098 9222 37110 9274
rect 37172 9222 37174 9274
rect 37012 9220 37036 9222
rect 37092 9220 37116 9222
rect 37172 9220 37196 9222
rect 36956 9200 37252 9220
rect 36084 9046 36136 9052
rect 36174 9072 36230 9081
rect 32140 8294 32168 9046
rect 32496 8968 32548 8974
rect 32496 8910 32548 8916
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 32508 8634 32536 8910
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32508 8537 32536 8570
rect 32494 8528 32550 8537
rect 35452 8498 35480 8910
rect 32494 8463 32550 8472
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35452 8401 35480 8434
rect 35438 8392 35494 8401
rect 35438 8327 35494 8336
rect 36096 8294 36124 9046
rect 36174 9007 36230 9016
rect 37648 8968 37700 8974
rect 37648 8910 37700 8916
rect 36360 8424 36412 8430
rect 36360 8366 36412 8372
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 36084 8288 36136 8294
rect 36084 8230 36136 8236
rect 32140 8129 32168 8230
rect 32126 8120 32182 8129
rect 36372 8090 36400 8366
rect 37660 8362 37688 8910
rect 36820 8356 36872 8362
rect 36820 8298 36872 8304
rect 37648 8356 37700 8362
rect 37648 8298 37700 8304
rect 36832 8265 36860 8298
rect 36818 8256 36874 8265
rect 36818 8191 36874 8200
rect 36956 8188 37252 8208
rect 37012 8186 37036 8188
rect 37092 8186 37116 8188
rect 37172 8186 37196 8188
rect 37034 8134 37036 8186
rect 37098 8134 37110 8186
rect 37172 8134 37174 8186
rect 37012 8132 37036 8134
rect 37092 8132 37116 8134
rect 37172 8132 37196 8134
rect 36956 8112 37252 8132
rect 32126 8055 32182 8064
rect 36360 8084 36412 8090
rect 36360 8026 36412 8032
rect 36372 7993 36400 8026
rect 36358 7984 36414 7993
rect 36358 7919 36414 7928
rect 36956 7100 37252 7120
rect 37012 7098 37036 7100
rect 37092 7098 37116 7100
rect 37172 7098 37196 7100
rect 37034 7046 37036 7098
rect 37098 7046 37110 7098
rect 37172 7046 37174 7098
rect 37012 7044 37036 7046
rect 37092 7044 37116 7046
rect 37172 7044 37196 7046
rect 36956 7024 37252 7044
rect 39316 6905 39344 9318
rect 49332 9318 49384 9324
rect 39946 9279 40002 9288
rect 49344 9178 49372 9318
rect 49332 9172 49384 9178
rect 49332 9114 49384 9120
rect 39764 9036 39816 9042
rect 39764 8978 39816 8984
rect 39776 8945 39804 8978
rect 39762 8936 39818 8945
rect 39762 8871 39818 8880
rect 40040 8424 40092 8430
rect 40040 8366 40092 8372
rect 40052 8265 40080 8366
rect 40038 8256 40094 8265
rect 40038 8191 40094 8200
rect 39302 6896 39358 6905
rect 39302 6831 39358 6840
rect 46938 6896 46994 6905
rect 46938 6831 46994 6840
rect 36956 6012 37252 6032
rect 37012 6010 37036 6012
rect 37092 6010 37116 6012
rect 37172 6010 37196 6012
rect 37034 5958 37036 6010
rect 37098 5958 37110 6010
rect 37172 5958 37174 6010
rect 37012 5956 37036 5958
rect 37092 5956 37116 5958
rect 37172 5956 37196 5958
rect 36956 5936 37252 5956
rect 36956 4924 37252 4944
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37034 4870 37036 4922
rect 37098 4870 37110 4922
rect 37172 4870 37174 4922
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 26606 4856 26662 4865
rect 26606 4791 26662 4800
rect 33782 4856 33838 4865
rect 36956 4848 37252 4868
rect 33782 4791 33838 4800
rect 18956 4380 19252 4400
rect 19012 4378 19036 4380
rect 19092 4378 19116 4380
rect 19172 4378 19196 4380
rect 19034 4326 19036 4378
rect 19098 4326 19110 4378
rect 19172 4326 19174 4378
rect 19012 4324 19036 4326
rect 19092 4324 19116 4326
rect 19172 4324 19196 4326
rect 18956 4304 19252 4324
rect 18956 3292 19252 3312
rect 19012 3290 19036 3292
rect 19092 3290 19116 3292
rect 19172 3290 19196 3292
rect 19034 3238 19036 3290
rect 19098 3238 19110 3290
rect 19172 3238 19174 3290
rect 19012 3236 19036 3238
rect 19092 3236 19116 3238
rect 19172 3236 19196 3238
rect 18956 3216 19252 3236
rect 19890 2816 19946 2825
rect 19890 2751 19946 2760
rect 18956 2204 19252 2224
rect 19012 2202 19036 2204
rect 19092 2202 19116 2204
rect 19172 2202 19196 2204
rect 19034 2150 19036 2202
rect 19098 2150 19110 2202
rect 19172 2150 19174 2202
rect 19012 2148 19036 2150
rect 19092 2148 19116 2150
rect 19172 2148 19196 2150
rect 18956 2128 19252 2148
rect 18326 1320 18382 1329
rect 18326 1255 18382 1264
rect 6734 82 6790 480
rect 6472 54 6790 82
rect 19904 82 19932 2751
rect 20166 82 20222 480
rect 19904 54 20222 82
rect 6734 0 6790 54
rect 20166 0 20222 54
rect 33690 82 33746 480
rect 33796 82 33824 4791
rect 36956 3836 37252 3856
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37034 3782 37036 3834
rect 37098 3782 37110 3834
rect 37172 3782 37174 3834
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 36956 3760 37252 3780
rect 36956 2748 37252 2768
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37034 2694 37036 2746
rect 37098 2694 37110 2746
rect 37172 2694 37174 2746
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 36956 2672 37252 2692
rect 33690 54 33824 82
rect 46952 82 46980 6831
rect 52380 6225 52408 10066
rect 52748 9722 52776 10066
rect 57348 10062 57376 13520
rect 61568 10124 61620 10130
rect 61568 10066 61620 10072
rect 57336 10056 57388 10062
rect 57336 9998 57388 10004
rect 61474 10024 61530 10033
rect 61474 9959 61530 9968
rect 61488 9926 61516 9959
rect 61476 9920 61528 9926
rect 61476 9862 61528 9868
rect 54956 9820 55252 9840
rect 55012 9818 55036 9820
rect 55092 9818 55116 9820
rect 55172 9818 55196 9820
rect 55034 9766 55036 9818
rect 55098 9766 55110 9818
rect 55172 9766 55174 9818
rect 55012 9764 55036 9766
rect 55092 9764 55116 9766
rect 55172 9764 55196 9766
rect 54956 9744 55252 9764
rect 61580 9722 61608 10066
rect 64064 10033 64092 13520
rect 66350 10976 66406 10985
rect 66350 10911 66406 10920
rect 66364 10266 66392 10911
rect 66352 10260 66404 10266
rect 66352 10202 66404 10208
rect 66260 10124 66312 10130
rect 66260 10066 66312 10072
rect 64050 10024 64106 10033
rect 61844 9988 61896 9994
rect 64050 9959 64106 9968
rect 61844 9930 61896 9936
rect 52736 9716 52788 9722
rect 52736 9658 52788 9664
rect 61568 9716 61620 9722
rect 61568 9658 61620 9664
rect 61856 9586 61884 9930
rect 61844 9580 61896 9586
rect 61844 9522 61896 9528
rect 61856 9489 61884 9522
rect 61842 9480 61898 9489
rect 61842 9415 61898 9424
rect 66272 9382 66300 10066
rect 70780 10062 70808 13520
rect 72956 11452 73252 11472
rect 73012 11450 73036 11452
rect 73092 11450 73116 11452
rect 73172 11450 73196 11452
rect 73034 11398 73036 11450
rect 73098 11398 73110 11450
rect 73172 11398 73174 11450
rect 73012 11396 73036 11398
rect 73092 11396 73116 11398
rect 73172 11396 73196 11398
rect 72956 11376 73252 11396
rect 77588 10985 77616 13520
rect 77574 10976 77630 10985
rect 77574 10911 77630 10920
rect 72956 10364 73252 10384
rect 73012 10362 73036 10364
rect 73092 10362 73116 10364
rect 73172 10362 73196 10364
rect 73034 10310 73036 10362
rect 73098 10310 73110 10362
rect 73172 10310 73174 10362
rect 73012 10308 73036 10310
rect 73092 10308 73116 10310
rect 73172 10308 73196 10310
rect 72956 10288 73252 10308
rect 79876 10260 79928 10266
rect 79876 10202 79928 10208
rect 79888 10169 79916 10202
rect 79874 10160 79930 10169
rect 79692 10124 79744 10130
rect 79874 10095 79930 10104
rect 79692 10066 79744 10072
rect 70768 10056 70820 10062
rect 70768 9998 70820 10004
rect 75184 10056 75236 10062
rect 75184 9998 75236 10004
rect 75460 10056 75512 10062
rect 75460 9998 75512 10004
rect 75196 9761 75224 9998
rect 75182 9752 75238 9761
rect 75182 9687 75238 9696
rect 75196 9654 75224 9687
rect 75184 9648 75236 9654
rect 75184 9590 75236 9596
rect 75472 9382 75500 9998
rect 78588 9920 78640 9926
rect 78588 9862 78640 9868
rect 78600 9382 78628 9862
rect 79704 9382 79732 10066
rect 84304 9761 84332 13520
rect 90744 13518 91048 13520
rect 89074 10704 89130 10713
rect 89074 10639 89130 10648
rect 87880 10124 87932 10130
rect 87880 10066 87932 10072
rect 84290 9752 84346 9761
rect 84290 9687 84346 9696
rect 87892 9382 87920 10066
rect 89088 10062 89116 10639
rect 90744 10169 90772 13518
rect 90956 10908 91252 10928
rect 91012 10906 91036 10908
rect 91092 10906 91116 10908
rect 91172 10906 91196 10908
rect 91034 10854 91036 10906
rect 91098 10854 91110 10906
rect 91172 10854 91174 10906
rect 91012 10852 91036 10854
rect 91092 10852 91116 10854
rect 91172 10852 91196 10854
rect 90956 10832 91252 10852
rect 97828 10713 97856 13520
rect 97814 10704 97870 10713
rect 97814 10639 97870 10648
rect 90730 10160 90786 10169
rect 90730 10095 90786 10104
rect 89076 10056 89128 10062
rect 89076 9998 89128 10004
rect 88708 9920 88760 9926
rect 88708 9862 88760 9868
rect 88720 9518 88748 9862
rect 89088 9722 89116 9998
rect 90956 9820 91252 9840
rect 91012 9818 91036 9820
rect 91092 9818 91116 9820
rect 91172 9818 91196 9820
rect 91034 9766 91036 9818
rect 91098 9766 91110 9818
rect 91172 9766 91174 9818
rect 91012 9764 91036 9766
rect 91092 9764 91116 9766
rect 91172 9764 91196 9766
rect 90956 9744 91252 9764
rect 89076 9716 89128 9722
rect 89076 9658 89128 9664
rect 88708 9512 88760 9518
rect 88246 9480 88302 9489
rect 104544 9489 104572 13520
rect 88708 9454 88760 9460
rect 104530 9480 104586 9489
rect 88246 9415 88302 9424
rect 88260 9382 88288 9415
rect 88720 9382 88748 9454
rect 104530 9415 104586 9424
rect 66260 9376 66312 9382
rect 66260 9318 66312 9324
rect 75460 9376 75512 9382
rect 75460 9318 75512 9324
rect 78588 9376 78640 9382
rect 78588 9318 78640 9324
rect 79692 9376 79744 9382
rect 79692 9318 79744 9324
rect 87880 9376 87932 9382
rect 87880 9318 87932 9324
rect 88248 9376 88300 9382
rect 88248 9318 88300 9324
rect 88708 9376 88760 9382
rect 88708 9318 88760 9324
rect 54956 8732 55252 8752
rect 55012 8730 55036 8732
rect 55092 8730 55116 8732
rect 55172 8730 55196 8732
rect 55034 8678 55036 8730
rect 55098 8678 55110 8730
rect 55172 8678 55174 8730
rect 55012 8676 55036 8678
rect 55092 8676 55116 8678
rect 55172 8676 55196 8678
rect 54956 8656 55252 8676
rect 66272 8265 66300 9318
rect 72956 9276 73252 9296
rect 73012 9274 73036 9276
rect 73092 9274 73116 9276
rect 73172 9274 73196 9276
rect 73034 9222 73036 9274
rect 73098 9222 73110 9274
rect 73172 9222 73174 9274
rect 73012 9220 73036 9222
rect 73092 9220 73116 9222
rect 73172 9220 73196 9222
rect 72956 9200 73252 9220
rect 75472 8945 75500 9318
rect 75458 8936 75514 8945
rect 75458 8871 75514 8880
rect 66258 8256 66314 8265
rect 66258 8191 66314 8200
rect 71870 8256 71926 8265
rect 71870 8191 71926 8200
rect 54956 7644 55252 7664
rect 55012 7642 55036 7644
rect 55092 7642 55116 7644
rect 55172 7642 55196 7644
rect 55034 7590 55036 7642
rect 55098 7590 55110 7642
rect 55172 7590 55174 7642
rect 55012 7588 55036 7590
rect 55092 7588 55116 7590
rect 55172 7588 55196 7590
rect 54956 7568 55252 7588
rect 54956 6556 55252 6576
rect 55012 6554 55036 6556
rect 55092 6554 55116 6556
rect 55172 6554 55196 6556
rect 55034 6502 55036 6554
rect 55098 6502 55110 6554
rect 55172 6502 55174 6554
rect 55012 6500 55036 6502
rect 55092 6500 55116 6502
rect 55172 6500 55196 6502
rect 54956 6480 55252 6500
rect 52366 6216 52422 6225
rect 52366 6151 52422 6160
rect 60830 6216 60886 6225
rect 60830 6151 60886 6160
rect 54956 5468 55252 5488
rect 55012 5466 55036 5468
rect 55092 5466 55116 5468
rect 55172 5466 55196 5468
rect 55034 5414 55036 5466
rect 55098 5414 55110 5466
rect 55172 5414 55174 5466
rect 55012 5412 55036 5414
rect 55092 5412 55116 5414
rect 55172 5412 55196 5414
rect 54956 5392 55252 5412
rect 54956 4380 55252 4400
rect 55012 4378 55036 4380
rect 55092 4378 55116 4380
rect 55172 4378 55196 4380
rect 55034 4326 55036 4378
rect 55098 4326 55110 4378
rect 55172 4326 55174 4378
rect 55012 4324 55036 4326
rect 55092 4324 55116 4326
rect 55172 4324 55196 4326
rect 54956 4304 55252 4324
rect 54956 3292 55252 3312
rect 55012 3290 55036 3292
rect 55092 3290 55116 3292
rect 55172 3290 55196 3292
rect 55034 3238 55036 3290
rect 55098 3238 55110 3290
rect 55172 3238 55174 3290
rect 55012 3236 55036 3238
rect 55092 3236 55116 3238
rect 55172 3236 55196 3238
rect 54956 3216 55252 3236
rect 54956 2204 55252 2224
rect 55012 2202 55036 2204
rect 55092 2202 55116 2204
rect 55172 2202 55196 2204
rect 55034 2150 55036 2202
rect 55098 2150 55110 2202
rect 55172 2150 55174 2202
rect 55012 2148 55036 2150
rect 55092 2148 55116 2150
rect 55172 2148 55196 2150
rect 54956 2128 55252 2148
rect 47214 82 47270 480
rect 46952 54 47270 82
rect 33690 0 33746 54
rect 47214 0 47270 54
rect 60738 82 60794 480
rect 60844 82 60872 6151
rect 71884 134 71912 8191
rect 72956 8188 73252 8208
rect 73012 8186 73036 8188
rect 73092 8186 73116 8188
rect 73172 8186 73196 8188
rect 73034 8134 73036 8186
rect 73098 8134 73110 8186
rect 73172 8134 73174 8186
rect 73012 8132 73036 8134
rect 73092 8132 73116 8134
rect 73172 8132 73196 8134
rect 72956 8112 73252 8132
rect 72956 7100 73252 7120
rect 73012 7098 73036 7100
rect 73092 7098 73116 7100
rect 73172 7098 73196 7100
rect 73034 7046 73036 7098
rect 73098 7046 73110 7098
rect 73172 7046 73174 7098
rect 73012 7044 73036 7046
rect 73092 7044 73116 7046
rect 73172 7044 73196 7046
rect 72956 7024 73252 7044
rect 72956 6012 73252 6032
rect 73012 6010 73036 6012
rect 73092 6010 73116 6012
rect 73172 6010 73196 6012
rect 73034 5958 73036 6010
rect 73098 5958 73110 6010
rect 73172 5958 73174 6010
rect 73012 5956 73036 5958
rect 73092 5956 73116 5958
rect 73172 5956 73196 5958
rect 72956 5936 73252 5956
rect 72956 4924 73252 4944
rect 73012 4922 73036 4924
rect 73092 4922 73116 4924
rect 73172 4922 73196 4924
rect 73034 4870 73036 4922
rect 73098 4870 73110 4922
rect 73172 4870 73174 4922
rect 73012 4868 73036 4870
rect 73092 4868 73116 4870
rect 73172 4868 73196 4870
rect 72956 4848 73252 4868
rect 72956 3836 73252 3856
rect 73012 3834 73036 3836
rect 73092 3834 73116 3836
rect 73172 3834 73196 3836
rect 73034 3782 73036 3834
rect 73098 3782 73110 3834
rect 73172 3782 73174 3834
rect 73012 3780 73036 3782
rect 73092 3780 73116 3782
rect 73172 3780 73196 3782
rect 72956 3760 73252 3780
rect 78600 2825 78628 9318
rect 87892 8401 87920 9318
rect 87878 8392 87934 8401
rect 87878 8327 87934 8336
rect 88720 8265 88748 9318
rect 90956 8732 91252 8752
rect 91012 8730 91036 8732
rect 91092 8730 91116 8732
rect 91172 8730 91196 8732
rect 91034 8678 91036 8730
rect 91098 8678 91110 8730
rect 91172 8678 91174 8730
rect 91012 8676 91036 8678
rect 91092 8676 91116 8678
rect 91172 8676 91196 8678
rect 90956 8656 91252 8676
rect 88706 8256 88762 8265
rect 88706 8191 88762 8200
rect 101310 8256 101366 8265
rect 101310 8191 101366 8200
rect 90956 7644 91252 7664
rect 91012 7642 91036 7644
rect 91092 7642 91116 7644
rect 91172 7642 91196 7644
rect 91034 7590 91036 7642
rect 91098 7590 91110 7642
rect 91172 7590 91174 7642
rect 91012 7588 91036 7590
rect 91092 7588 91116 7590
rect 91172 7588 91196 7590
rect 90956 7568 91252 7588
rect 90956 6556 91252 6576
rect 91012 6554 91036 6556
rect 91092 6554 91116 6556
rect 91172 6554 91196 6556
rect 91034 6502 91036 6554
rect 91098 6502 91110 6554
rect 91172 6502 91174 6554
rect 91012 6500 91036 6502
rect 91092 6500 91116 6502
rect 91172 6500 91196 6502
rect 90956 6480 91252 6500
rect 90956 5468 91252 5488
rect 91012 5466 91036 5468
rect 91092 5466 91116 5468
rect 91172 5466 91196 5468
rect 91034 5414 91036 5466
rect 91098 5414 91110 5466
rect 91172 5414 91174 5466
rect 91012 5412 91036 5414
rect 91092 5412 91116 5414
rect 91172 5412 91196 5414
rect 90956 5392 91252 5412
rect 90956 4380 91252 4400
rect 91012 4378 91036 4380
rect 91092 4378 91116 4380
rect 91172 4378 91196 4380
rect 91034 4326 91036 4378
rect 91098 4326 91110 4378
rect 91172 4326 91174 4378
rect 91012 4324 91036 4326
rect 91092 4324 91116 4326
rect 91172 4324 91196 4326
rect 90956 4304 91252 4324
rect 90956 3292 91252 3312
rect 91012 3290 91036 3292
rect 91092 3290 91116 3292
rect 91172 3290 91196 3292
rect 91034 3238 91036 3290
rect 91098 3238 91110 3290
rect 91172 3238 91174 3290
rect 91012 3236 91036 3238
rect 91092 3236 91116 3238
rect 91172 3236 91196 3238
rect 90956 3216 91252 3236
rect 78586 2816 78642 2825
rect 72956 2748 73252 2768
rect 78586 2751 78642 2760
rect 87418 2816 87474 2825
rect 87418 2751 87474 2760
rect 73012 2746 73036 2748
rect 73092 2746 73116 2748
rect 73172 2746 73196 2748
rect 73034 2694 73036 2746
rect 73098 2694 73110 2746
rect 73172 2694 73174 2746
rect 73012 2692 73036 2694
rect 73092 2692 73116 2694
rect 73172 2692 73196 2694
rect 72956 2672 73252 2692
rect 60738 54 60872 82
rect 71872 128 71924 134
rect 71872 70 71924 76
rect 74170 128 74226 480
rect 74170 76 74172 128
rect 74224 76 74226 128
rect 60738 0 60794 54
rect 74170 0 74226 76
rect 87432 82 87460 2751
rect 90956 2204 91252 2224
rect 91012 2202 91036 2204
rect 91092 2202 91116 2204
rect 91172 2202 91196 2204
rect 91034 2150 91036 2202
rect 91098 2150 91110 2202
rect 91172 2150 91174 2202
rect 91012 2148 91036 2150
rect 91092 2148 91116 2150
rect 91172 2148 91196 2150
rect 90956 2128 91252 2148
rect 87694 82 87750 480
rect 87432 54 87750 82
rect 87694 0 87750 54
rect 101218 82 101274 480
rect 101324 82 101352 8191
rect 101218 54 101352 82
rect 101218 0 101274 54
<< via2 >>
rect 1490 12144 1546 12200
rect 110 10376 166 10432
rect 1674 10920 1730 10976
rect 1490 9152 1546 9208
rect 10046 10920 10102 10976
rect 21822 10920 21878 10976
rect 18956 10906 19012 10908
rect 19036 10906 19092 10908
rect 19116 10906 19172 10908
rect 19196 10906 19252 10908
rect 18956 10854 18982 10906
rect 18982 10854 19012 10906
rect 19036 10854 19046 10906
rect 19046 10854 19092 10906
rect 19116 10854 19162 10906
rect 19162 10854 19172 10906
rect 19196 10854 19226 10906
rect 19226 10854 19252 10906
rect 18956 10852 19012 10854
rect 19036 10852 19092 10854
rect 19116 10852 19172 10854
rect 19196 10852 19252 10854
rect 12898 10104 12954 10160
rect 110 8880 166 8936
rect 110 8336 166 8392
rect 110 8064 166 8120
rect 18956 9818 19012 9820
rect 19036 9818 19092 9820
rect 19116 9818 19172 9820
rect 19196 9818 19252 9820
rect 18956 9766 18982 9818
rect 18982 9766 19012 9818
rect 19036 9766 19046 9818
rect 19046 9766 19092 9818
rect 19116 9766 19162 9818
rect 19162 9766 19172 9818
rect 19196 9766 19226 9818
rect 19226 9766 19252 9818
rect 18956 9764 19012 9766
rect 19036 9764 19092 9766
rect 19116 9764 19172 9766
rect 19196 9764 19252 9766
rect 30286 10920 30342 10976
rect 36956 11450 37012 11452
rect 37036 11450 37092 11452
rect 37116 11450 37172 11452
rect 37196 11450 37252 11452
rect 36956 11398 36982 11450
rect 36982 11398 37012 11450
rect 37036 11398 37046 11450
rect 37046 11398 37092 11450
rect 37116 11398 37162 11450
rect 37162 11398 37172 11450
rect 37196 11398 37226 11450
rect 37226 11398 37252 11450
rect 36956 11396 37012 11398
rect 37036 11396 37092 11398
rect 37116 11396 37172 11398
rect 37196 11396 37252 11398
rect 36956 10362 37012 10364
rect 37036 10362 37092 10364
rect 37116 10362 37172 10364
rect 37196 10362 37252 10364
rect 36956 10310 36982 10362
rect 36982 10310 37012 10362
rect 37036 10310 37046 10362
rect 37046 10310 37092 10362
rect 37116 10310 37162 10362
rect 37162 10310 37172 10362
rect 37196 10310 37226 10362
rect 37226 10310 37252 10362
rect 36956 10308 37012 10310
rect 37036 10308 37092 10310
rect 37116 10308 37172 10310
rect 37196 10308 37252 10310
rect 26698 10104 26754 10160
rect 36818 10104 36874 10160
rect 39394 10104 39450 10160
rect 23570 9968 23626 10024
rect 35162 9696 35218 9752
rect 11426 9152 11482 9208
rect 9126 8336 9182 8392
rect 10782 8200 10838 8256
rect 9494 6296 9550 6352
rect 15290 8880 15346 8936
rect 18956 8730 19012 8732
rect 19036 8730 19092 8732
rect 19116 8730 19172 8732
rect 19196 8730 19252 8732
rect 18956 8678 18982 8730
rect 18982 8678 19012 8730
rect 19036 8678 19046 8730
rect 19046 8678 19092 8730
rect 19116 8678 19162 8730
rect 19162 8678 19172 8730
rect 19196 8678 19226 8730
rect 19226 8678 19252 8730
rect 18956 8676 19012 8678
rect 19036 8676 19092 8678
rect 19116 8676 19172 8678
rect 19196 8676 19252 8678
rect 18956 7642 19012 7644
rect 19036 7642 19092 7644
rect 19116 7642 19172 7644
rect 19196 7642 19252 7644
rect 18956 7590 18982 7642
rect 18982 7590 19012 7642
rect 19036 7590 19046 7642
rect 19046 7590 19092 7642
rect 19116 7590 19162 7642
rect 19162 7590 19172 7642
rect 19196 7590 19226 7642
rect 19226 7590 19252 7642
rect 18956 7588 19012 7590
rect 19036 7588 19092 7590
rect 19116 7588 19172 7590
rect 19196 7588 19252 7590
rect 21270 8472 21326 8528
rect 19798 8064 19854 8120
rect 23202 9016 23258 9072
rect 21914 8336 21970 8392
rect 23662 8200 23718 8256
rect 23110 7928 23166 7984
rect 18956 6554 19012 6556
rect 19036 6554 19092 6556
rect 19116 6554 19172 6556
rect 19196 6554 19252 6556
rect 18956 6502 18982 6554
rect 18982 6502 19012 6554
rect 19036 6502 19046 6554
rect 19046 6502 19092 6554
rect 19116 6502 19162 6554
rect 19162 6502 19172 6554
rect 19196 6502 19226 6554
rect 19226 6502 19252 6554
rect 18956 6500 19012 6502
rect 19036 6500 19092 6502
rect 19116 6500 19172 6502
rect 19196 6500 19252 6502
rect 12714 2760 12770 2816
rect 18956 5466 19012 5468
rect 19036 5466 19092 5468
rect 19116 5466 19172 5468
rect 19196 5466 19252 5468
rect 18956 5414 18982 5466
rect 18982 5414 19012 5466
rect 19036 5414 19046 5466
rect 19046 5414 19092 5466
rect 19116 5414 19162 5466
rect 19162 5414 19172 5466
rect 19196 5414 19226 5466
rect 19226 5414 19252 5466
rect 18956 5412 19012 5414
rect 19036 5412 19092 5414
rect 19116 5412 19172 5414
rect 19196 5412 19252 5414
rect 54956 10906 55012 10908
rect 55036 10906 55092 10908
rect 55116 10906 55172 10908
rect 55196 10906 55252 10908
rect 54956 10854 54982 10906
rect 54982 10854 55012 10906
rect 55036 10854 55046 10906
rect 55046 10854 55092 10906
rect 55116 10854 55162 10906
rect 55162 10854 55172 10906
rect 55196 10854 55226 10906
rect 55226 10854 55252 10906
rect 54956 10852 55012 10854
rect 55036 10852 55092 10854
rect 55116 10852 55172 10854
rect 55196 10852 55252 10854
rect 50526 10104 50582 10160
rect 43810 9696 43866 9752
rect 36956 9274 37012 9276
rect 37036 9274 37092 9276
rect 37116 9274 37172 9276
rect 37196 9274 37252 9276
rect 36956 9222 36982 9274
rect 36982 9222 37012 9274
rect 37036 9222 37046 9274
rect 37046 9222 37092 9274
rect 37116 9222 37162 9274
rect 37162 9222 37172 9274
rect 37196 9222 37226 9274
rect 37226 9222 37252 9274
rect 36956 9220 37012 9222
rect 37036 9220 37092 9222
rect 37116 9220 37172 9222
rect 37196 9220 37252 9222
rect 32494 8472 32550 8528
rect 35438 8336 35494 8392
rect 36174 9016 36230 9072
rect 32126 8064 32182 8120
rect 36818 8200 36874 8256
rect 36956 8186 37012 8188
rect 37036 8186 37092 8188
rect 37116 8186 37172 8188
rect 37196 8186 37252 8188
rect 36956 8134 36982 8186
rect 36982 8134 37012 8186
rect 37036 8134 37046 8186
rect 37046 8134 37092 8186
rect 37116 8134 37162 8186
rect 37162 8134 37172 8186
rect 37196 8134 37226 8186
rect 37226 8134 37252 8186
rect 36956 8132 37012 8134
rect 37036 8132 37092 8134
rect 37116 8132 37172 8134
rect 37196 8132 37252 8134
rect 36358 7928 36414 7984
rect 36956 7098 37012 7100
rect 37036 7098 37092 7100
rect 37116 7098 37172 7100
rect 37196 7098 37252 7100
rect 36956 7046 36982 7098
rect 36982 7046 37012 7098
rect 37036 7046 37046 7098
rect 37046 7046 37092 7098
rect 37116 7046 37162 7098
rect 37162 7046 37172 7098
rect 37196 7046 37226 7098
rect 37226 7046 37252 7098
rect 36956 7044 37012 7046
rect 37036 7044 37092 7046
rect 37116 7044 37172 7046
rect 37196 7044 37252 7046
rect 39946 9288 40002 9344
rect 39762 8880 39818 8936
rect 40038 8200 40094 8256
rect 39302 6840 39358 6896
rect 46938 6840 46994 6896
rect 36956 6010 37012 6012
rect 37036 6010 37092 6012
rect 37116 6010 37172 6012
rect 37196 6010 37252 6012
rect 36956 5958 36982 6010
rect 36982 5958 37012 6010
rect 37036 5958 37046 6010
rect 37046 5958 37092 6010
rect 37116 5958 37162 6010
rect 37162 5958 37172 6010
rect 37196 5958 37226 6010
rect 37226 5958 37252 6010
rect 36956 5956 37012 5958
rect 37036 5956 37092 5958
rect 37116 5956 37172 5958
rect 37196 5956 37252 5958
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 36982 4922
rect 36982 4870 37012 4922
rect 37036 4870 37046 4922
rect 37046 4870 37092 4922
rect 37116 4870 37162 4922
rect 37162 4870 37172 4922
rect 37196 4870 37226 4922
rect 37226 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 26606 4800 26662 4856
rect 33782 4800 33838 4856
rect 18956 4378 19012 4380
rect 19036 4378 19092 4380
rect 19116 4378 19172 4380
rect 19196 4378 19252 4380
rect 18956 4326 18982 4378
rect 18982 4326 19012 4378
rect 19036 4326 19046 4378
rect 19046 4326 19092 4378
rect 19116 4326 19162 4378
rect 19162 4326 19172 4378
rect 19196 4326 19226 4378
rect 19226 4326 19252 4378
rect 18956 4324 19012 4326
rect 19036 4324 19092 4326
rect 19116 4324 19172 4326
rect 19196 4324 19252 4326
rect 18956 3290 19012 3292
rect 19036 3290 19092 3292
rect 19116 3290 19172 3292
rect 19196 3290 19252 3292
rect 18956 3238 18982 3290
rect 18982 3238 19012 3290
rect 19036 3238 19046 3290
rect 19046 3238 19092 3290
rect 19116 3238 19162 3290
rect 19162 3238 19172 3290
rect 19196 3238 19226 3290
rect 19226 3238 19252 3290
rect 18956 3236 19012 3238
rect 19036 3236 19092 3238
rect 19116 3236 19172 3238
rect 19196 3236 19252 3238
rect 19890 2760 19946 2816
rect 18956 2202 19012 2204
rect 19036 2202 19092 2204
rect 19116 2202 19172 2204
rect 19196 2202 19252 2204
rect 18956 2150 18982 2202
rect 18982 2150 19012 2202
rect 19036 2150 19046 2202
rect 19046 2150 19092 2202
rect 19116 2150 19162 2202
rect 19162 2150 19172 2202
rect 19196 2150 19226 2202
rect 19226 2150 19252 2202
rect 18956 2148 19012 2150
rect 19036 2148 19092 2150
rect 19116 2148 19172 2150
rect 19196 2148 19252 2150
rect 18326 1264 18382 1320
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 36982 3834
rect 36982 3782 37012 3834
rect 37036 3782 37046 3834
rect 37046 3782 37092 3834
rect 37116 3782 37162 3834
rect 37162 3782 37172 3834
rect 37196 3782 37226 3834
rect 37226 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 36982 2746
rect 36982 2694 37012 2746
rect 37036 2694 37046 2746
rect 37046 2694 37092 2746
rect 37116 2694 37162 2746
rect 37162 2694 37172 2746
rect 37196 2694 37226 2746
rect 37226 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 61474 9968 61530 10024
rect 54956 9818 55012 9820
rect 55036 9818 55092 9820
rect 55116 9818 55172 9820
rect 55196 9818 55252 9820
rect 54956 9766 54982 9818
rect 54982 9766 55012 9818
rect 55036 9766 55046 9818
rect 55046 9766 55092 9818
rect 55116 9766 55162 9818
rect 55162 9766 55172 9818
rect 55196 9766 55226 9818
rect 55226 9766 55252 9818
rect 54956 9764 55012 9766
rect 55036 9764 55092 9766
rect 55116 9764 55172 9766
rect 55196 9764 55252 9766
rect 66350 10920 66406 10976
rect 64050 9968 64106 10024
rect 61842 9424 61898 9480
rect 72956 11450 73012 11452
rect 73036 11450 73092 11452
rect 73116 11450 73172 11452
rect 73196 11450 73252 11452
rect 72956 11398 72982 11450
rect 72982 11398 73012 11450
rect 73036 11398 73046 11450
rect 73046 11398 73092 11450
rect 73116 11398 73162 11450
rect 73162 11398 73172 11450
rect 73196 11398 73226 11450
rect 73226 11398 73252 11450
rect 72956 11396 73012 11398
rect 73036 11396 73092 11398
rect 73116 11396 73172 11398
rect 73196 11396 73252 11398
rect 77574 10920 77630 10976
rect 72956 10362 73012 10364
rect 73036 10362 73092 10364
rect 73116 10362 73172 10364
rect 73196 10362 73252 10364
rect 72956 10310 72982 10362
rect 72982 10310 73012 10362
rect 73036 10310 73046 10362
rect 73046 10310 73092 10362
rect 73116 10310 73162 10362
rect 73162 10310 73172 10362
rect 73196 10310 73226 10362
rect 73226 10310 73252 10362
rect 72956 10308 73012 10310
rect 73036 10308 73092 10310
rect 73116 10308 73172 10310
rect 73196 10308 73252 10310
rect 79874 10104 79930 10160
rect 75182 9696 75238 9752
rect 89074 10648 89130 10704
rect 84290 9696 84346 9752
rect 90956 10906 91012 10908
rect 91036 10906 91092 10908
rect 91116 10906 91172 10908
rect 91196 10906 91252 10908
rect 90956 10854 90982 10906
rect 90982 10854 91012 10906
rect 91036 10854 91046 10906
rect 91046 10854 91092 10906
rect 91116 10854 91162 10906
rect 91162 10854 91172 10906
rect 91196 10854 91226 10906
rect 91226 10854 91252 10906
rect 90956 10852 91012 10854
rect 91036 10852 91092 10854
rect 91116 10852 91172 10854
rect 91196 10852 91252 10854
rect 97814 10648 97870 10704
rect 90730 10104 90786 10160
rect 90956 9818 91012 9820
rect 91036 9818 91092 9820
rect 91116 9818 91172 9820
rect 91196 9818 91252 9820
rect 90956 9766 90982 9818
rect 90982 9766 91012 9818
rect 91036 9766 91046 9818
rect 91046 9766 91092 9818
rect 91116 9766 91162 9818
rect 91162 9766 91172 9818
rect 91196 9766 91226 9818
rect 91226 9766 91252 9818
rect 90956 9764 91012 9766
rect 91036 9764 91092 9766
rect 91116 9764 91172 9766
rect 91196 9764 91252 9766
rect 88246 9424 88302 9480
rect 104530 9424 104586 9480
rect 54956 8730 55012 8732
rect 55036 8730 55092 8732
rect 55116 8730 55172 8732
rect 55196 8730 55252 8732
rect 54956 8678 54982 8730
rect 54982 8678 55012 8730
rect 55036 8678 55046 8730
rect 55046 8678 55092 8730
rect 55116 8678 55162 8730
rect 55162 8678 55172 8730
rect 55196 8678 55226 8730
rect 55226 8678 55252 8730
rect 54956 8676 55012 8678
rect 55036 8676 55092 8678
rect 55116 8676 55172 8678
rect 55196 8676 55252 8678
rect 72956 9274 73012 9276
rect 73036 9274 73092 9276
rect 73116 9274 73172 9276
rect 73196 9274 73252 9276
rect 72956 9222 72982 9274
rect 72982 9222 73012 9274
rect 73036 9222 73046 9274
rect 73046 9222 73092 9274
rect 73116 9222 73162 9274
rect 73162 9222 73172 9274
rect 73196 9222 73226 9274
rect 73226 9222 73252 9274
rect 72956 9220 73012 9222
rect 73036 9220 73092 9222
rect 73116 9220 73172 9222
rect 73196 9220 73252 9222
rect 75458 8880 75514 8936
rect 66258 8200 66314 8256
rect 71870 8200 71926 8256
rect 54956 7642 55012 7644
rect 55036 7642 55092 7644
rect 55116 7642 55172 7644
rect 55196 7642 55252 7644
rect 54956 7590 54982 7642
rect 54982 7590 55012 7642
rect 55036 7590 55046 7642
rect 55046 7590 55092 7642
rect 55116 7590 55162 7642
rect 55162 7590 55172 7642
rect 55196 7590 55226 7642
rect 55226 7590 55252 7642
rect 54956 7588 55012 7590
rect 55036 7588 55092 7590
rect 55116 7588 55172 7590
rect 55196 7588 55252 7590
rect 54956 6554 55012 6556
rect 55036 6554 55092 6556
rect 55116 6554 55172 6556
rect 55196 6554 55252 6556
rect 54956 6502 54982 6554
rect 54982 6502 55012 6554
rect 55036 6502 55046 6554
rect 55046 6502 55092 6554
rect 55116 6502 55162 6554
rect 55162 6502 55172 6554
rect 55196 6502 55226 6554
rect 55226 6502 55252 6554
rect 54956 6500 55012 6502
rect 55036 6500 55092 6502
rect 55116 6500 55172 6502
rect 55196 6500 55252 6502
rect 52366 6160 52422 6216
rect 60830 6160 60886 6216
rect 54956 5466 55012 5468
rect 55036 5466 55092 5468
rect 55116 5466 55172 5468
rect 55196 5466 55252 5468
rect 54956 5414 54982 5466
rect 54982 5414 55012 5466
rect 55036 5414 55046 5466
rect 55046 5414 55092 5466
rect 55116 5414 55162 5466
rect 55162 5414 55172 5466
rect 55196 5414 55226 5466
rect 55226 5414 55252 5466
rect 54956 5412 55012 5414
rect 55036 5412 55092 5414
rect 55116 5412 55172 5414
rect 55196 5412 55252 5414
rect 54956 4378 55012 4380
rect 55036 4378 55092 4380
rect 55116 4378 55172 4380
rect 55196 4378 55252 4380
rect 54956 4326 54982 4378
rect 54982 4326 55012 4378
rect 55036 4326 55046 4378
rect 55046 4326 55092 4378
rect 55116 4326 55162 4378
rect 55162 4326 55172 4378
rect 55196 4326 55226 4378
rect 55226 4326 55252 4378
rect 54956 4324 55012 4326
rect 55036 4324 55092 4326
rect 55116 4324 55172 4326
rect 55196 4324 55252 4326
rect 54956 3290 55012 3292
rect 55036 3290 55092 3292
rect 55116 3290 55172 3292
rect 55196 3290 55252 3292
rect 54956 3238 54982 3290
rect 54982 3238 55012 3290
rect 55036 3238 55046 3290
rect 55046 3238 55092 3290
rect 55116 3238 55162 3290
rect 55162 3238 55172 3290
rect 55196 3238 55226 3290
rect 55226 3238 55252 3290
rect 54956 3236 55012 3238
rect 55036 3236 55092 3238
rect 55116 3236 55172 3238
rect 55196 3236 55252 3238
rect 54956 2202 55012 2204
rect 55036 2202 55092 2204
rect 55116 2202 55172 2204
rect 55196 2202 55252 2204
rect 54956 2150 54982 2202
rect 54982 2150 55012 2202
rect 55036 2150 55046 2202
rect 55046 2150 55092 2202
rect 55116 2150 55162 2202
rect 55162 2150 55172 2202
rect 55196 2150 55226 2202
rect 55226 2150 55252 2202
rect 54956 2148 55012 2150
rect 55036 2148 55092 2150
rect 55116 2148 55172 2150
rect 55196 2148 55252 2150
rect 72956 8186 73012 8188
rect 73036 8186 73092 8188
rect 73116 8186 73172 8188
rect 73196 8186 73252 8188
rect 72956 8134 72982 8186
rect 72982 8134 73012 8186
rect 73036 8134 73046 8186
rect 73046 8134 73092 8186
rect 73116 8134 73162 8186
rect 73162 8134 73172 8186
rect 73196 8134 73226 8186
rect 73226 8134 73252 8186
rect 72956 8132 73012 8134
rect 73036 8132 73092 8134
rect 73116 8132 73172 8134
rect 73196 8132 73252 8134
rect 72956 7098 73012 7100
rect 73036 7098 73092 7100
rect 73116 7098 73172 7100
rect 73196 7098 73252 7100
rect 72956 7046 72982 7098
rect 72982 7046 73012 7098
rect 73036 7046 73046 7098
rect 73046 7046 73092 7098
rect 73116 7046 73162 7098
rect 73162 7046 73172 7098
rect 73196 7046 73226 7098
rect 73226 7046 73252 7098
rect 72956 7044 73012 7046
rect 73036 7044 73092 7046
rect 73116 7044 73172 7046
rect 73196 7044 73252 7046
rect 72956 6010 73012 6012
rect 73036 6010 73092 6012
rect 73116 6010 73172 6012
rect 73196 6010 73252 6012
rect 72956 5958 72982 6010
rect 72982 5958 73012 6010
rect 73036 5958 73046 6010
rect 73046 5958 73092 6010
rect 73116 5958 73162 6010
rect 73162 5958 73172 6010
rect 73196 5958 73226 6010
rect 73226 5958 73252 6010
rect 72956 5956 73012 5958
rect 73036 5956 73092 5958
rect 73116 5956 73172 5958
rect 73196 5956 73252 5958
rect 72956 4922 73012 4924
rect 73036 4922 73092 4924
rect 73116 4922 73172 4924
rect 73196 4922 73252 4924
rect 72956 4870 72982 4922
rect 72982 4870 73012 4922
rect 73036 4870 73046 4922
rect 73046 4870 73092 4922
rect 73116 4870 73162 4922
rect 73162 4870 73172 4922
rect 73196 4870 73226 4922
rect 73226 4870 73252 4922
rect 72956 4868 73012 4870
rect 73036 4868 73092 4870
rect 73116 4868 73172 4870
rect 73196 4868 73252 4870
rect 72956 3834 73012 3836
rect 73036 3834 73092 3836
rect 73116 3834 73172 3836
rect 73196 3834 73252 3836
rect 72956 3782 72982 3834
rect 72982 3782 73012 3834
rect 73036 3782 73046 3834
rect 73046 3782 73092 3834
rect 73116 3782 73162 3834
rect 73162 3782 73172 3834
rect 73196 3782 73226 3834
rect 73226 3782 73252 3834
rect 72956 3780 73012 3782
rect 73036 3780 73092 3782
rect 73116 3780 73172 3782
rect 73196 3780 73252 3782
rect 87878 8336 87934 8392
rect 90956 8730 91012 8732
rect 91036 8730 91092 8732
rect 91116 8730 91172 8732
rect 91196 8730 91252 8732
rect 90956 8678 90982 8730
rect 90982 8678 91012 8730
rect 91036 8678 91046 8730
rect 91046 8678 91092 8730
rect 91116 8678 91162 8730
rect 91162 8678 91172 8730
rect 91196 8678 91226 8730
rect 91226 8678 91252 8730
rect 90956 8676 91012 8678
rect 91036 8676 91092 8678
rect 91116 8676 91172 8678
rect 91196 8676 91252 8678
rect 88706 8200 88762 8256
rect 101310 8200 101366 8256
rect 90956 7642 91012 7644
rect 91036 7642 91092 7644
rect 91116 7642 91172 7644
rect 91196 7642 91252 7644
rect 90956 7590 90982 7642
rect 90982 7590 91012 7642
rect 91036 7590 91046 7642
rect 91046 7590 91092 7642
rect 91116 7590 91162 7642
rect 91162 7590 91172 7642
rect 91196 7590 91226 7642
rect 91226 7590 91252 7642
rect 90956 7588 91012 7590
rect 91036 7588 91092 7590
rect 91116 7588 91172 7590
rect 91196 7588 91252 7590
rect 90956 6554 91012 6556
rect 91036 6554 91092 6556
rect 91116 6554 91172 6556
rect 91196 6554 91252 6556
rect 90956 6502 90982 6554
rect 90982 6502 91012 6554
rect 91036 6502 91046 6554
rect 91046 6502 91092 6554
rect 91116 6502 91162 6554
rect 91162 6502 91172 6554
rect 91196 6502 91226 6554
rect 91226 6502 91252 6554
rect 90956 6500 91012 6502
rect 91036 6500 91092 6502
rect 91116 6500 91172 6502
rect 91196 6500 91252 6502
rect 90956 5466 91012 5468
rect 91036 5466 91092 5468
rect 91116 5466 91172 5468
rect 91196 5466 91252 5468
rect 90956 5414 90982 5466
rect 90982 5414 91012 5466
rect 91036 5414 91046 5466
rect 91046 5414 91092 5466
rect 91116 5414 91162 5466
rect 91162 5414 91172 5466
rect 91196 5414 91226 5466
rect 91226 5414 91252 5466
rect 90956 5412 91012 5414
rect 91036 5412 91092 5414
rect 91116 5412 91172 5414
rect 91196 5412 91252 5414
rect 90956 4378 91012 4380
rect 91036 4378 91092 4380
rect 91116 4378 91172 4380
rect 91196 4378 91252 4380
rect 90956 4326 90982 4378
rect 90982 4326 91012 4378
rect 91036 4326 91046 4378
rect 91046 4326 91092 4378
rect 91116 4326 91162 4378
rect 91162 4326 91172 4378
rect 91196 4326 91226 4378
rect 91226 4326 91252 4378
rect 90956 4324 91012 4326
rect 91036 4324 91092 4326
rect 91116 4324 91172 4326
rect 91196 4324 91252 4326
rect 90956 3290 91012 3292
rect 91036 3290 91092 3292
rect 91116 3290 91172 3292
rect 91196 3290 91252 3292
rect 90956 3238 90982 3290
rect 90982 3238 91012 3290
rect 91036 3238 91046 3290
rect 91046 3238 91092 3290
rect 91116 3238 91162 3290
rect 91162 3238 91172 3290
rect 91196 3238 91226 3290
rect 91226 3238 91252 3290
rect 90956 3236 91012 3238
rect 91036 3236 91092 3238
rect 91116 3236 91172 3238
rect 91196 3236 91252 3238
rect 78586 2760 78642 2816
rect 87418 2760 87474 2816
rect 72956 2746 73012 2748
rect 73036 2746 73092 2748
rect 73116 2746 73172 2748
rect 73196 2746 73252 2748
rect 72956 2694 72982 2746
rect 72982 2694 73012 2746
rect 73036 2694 73046 2746
rect 73046 2694 73092 2746
rect 73116 2694 73162 2746
rect 73162 2694 73172 2746
rect 73196 2694 73226 2746
rect 73226 2694 73252 2746
rect 72956 2692 73012 2694
rect 73036 2692 73092 2694
rect 73116 2692 73172 2694
rect 73196 2692 73252 2694
rect 90956 2202 91012 2204
rect 91036 2202 91092 2204
rect 91116 2202 91172 2204
rect 91196 2202 91252 2204
rect 90956 2150 90982 2202
rect 90982 2150 91012 2202
rect 91036 2150 91046 2202
rect 91046 2150 91092 2202
rect 91116 2150 91162 2202
rect 91162 2150 91172 2202
rect 91196 2150 91226 2202
rect 91226 2150 91252 2202
rect 90956 2148 91012 2150
rect 91036 2148 91092 2150
rect 91116 2148 91172 2150
rect 91196 2148 91252 2150
<< metal3 >>
rect 0 12656 480 12776
rect 62 12202 122 12656
rect 1485 12202 1551 12205
rect 62 12200 1551 12202
rect 62 12144 1490 12200
rect 1546 12144 1551 12200
rect 62 12142 1551 12144
rect 1485 12139 1551 12142
rect 36944 11456 37264 11457
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 11391 37264 11392
rect 72944 11456 73264 11457
rect 72944 11392 72952 11456
rect 73016 11392 73032 11456
rect 73096 11392 73112 11456
rect 73176 11392 73192 11456
rect 73256 11392 73264 11456
rect 72944 11391 73264 11392
rect 1669 10978 1735 10981
rect 10041 10978 10107 10981
rect 1669 10976 10107 10978
rect 1669 10920 1674 10976
rect 1730 10920 10046 10976
rect 10102 10920 10107 10976
rect 1669 10918 10107 10920
rect 1669 10915 1735 10918
rect 10041 10915 10107 10918
rect 21817 10978 21883 10981
rect 30281 10978 30347 10981
rect 21817 10976 30347 10978
rect 21817 10920 21822 10976
rect 21878 10920 30286 10976
rect 30342 10920 30347 10976
rect 21817 10918 30347 10920
rect 21817 10915 21883 10918
rect 30281 10915 30347 10918
rect 66345 10978 66411 10981
rect 77569 10978 77635 10981
rect 66345 10976 77635 10978
rect 66345 10920 66350 10976
rect 66406 10920 77574 10976
rect 77630 10920 77635 10976
rect 66345 10918 77635 10920
rect 66345 10915 66411 10918
rect 77569 10915 77635 10918
rect 18944 10912 19264 10913
rect 18944 10848 18952 10912
rect 19016 10848 19032 10912
rect 19096 10848 19112 10912
rect 19176 10848 19192 10912
rect 19256 10848 19264 10912
rect 18944 10847 19264 10848
rect 54944 10912 55264 10913
rect 54944 10848 54952 10912
rect 55016 10848 55032 10912
rect 55096 10848 55112 10912
rect 55176 10848 55192 10912
rect 55256 10848 55264 10912
rect 54944 10847 55264 10848
rect 90944 10912 91264 10913
rect 90944 10848 90952 10912
rect 91016 10848 91032 10912
rect 91096 10848 91112 10912
rect 91176 10848 91192 10912
rect 91256 10848 91264 10912
rect 90944 10847 91264 10848
rect 89069 10706 89135 10709
rect 97809 10706 97875 10709
rect 89069 10704 97875 10706
rect 89069 10648 89074 10704
rect 89130 10648 97814 10704
rect 97870 10648 97875 10704
rect 89069 10646 97875 10648
rect 89069 10643 89135 10646
rect 97809 10643 97875 10646
rect 0 10432 480 10464
rect 0 10376 110 10432
rect 166 10376 480 10432
rect 0 10344 480 10376
rect 36944 10368 37264 10369
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 10303 37264 10304
rect 72944 10368 73264 10369
rect 72944 10304 72952 10368
rect 73016 10304 73032 10368
rect 73096 10304 73112 10368
rect 73176 10304 73192 10368
rect 73256 10304 73264 10368
rect 72944 10303 73264 10304
rect 12893 10162 12959 10165
rect 26693 10162 26759 10165
rect 36813 10162 36879 10165
rect 12893 10160 13830 10162
rect 12893 10104 12898 10160
rect 12954 10104 13830 10160
rect 12893 10102 13830 10104
rect 12893 10099 12959 10102
rect 13770 10026 13830 10102
rect 26693 10160 36879 10162
rect 26693 10104 26698 10160
rect 26754 10104 36818 10160
rect 36874 10104 36879 10160
rect 26693 10102 36879 10104
rect 26693 10099 26759 10102
rect 36813 10099 36879 10102
rect 39389 10162 39455 10165
rect 50521 10162 50587 10165
rect 39389 10160 50587 10162
rect 39389 10104 39394 10160
rect 39450 10104 50526 10160
rect 50582 10104 50587 10160
rect 39389 10102 50587 10104
rect 39389 10099 39455 10102
rect 50521 10099 50587 10102
rect 79869 10162 79935 10165
rect 90725 10162 90791 10165
rect 79869 10160 90791 10162
rect 79869 10104 79874 10160
rect 79930 10104 90730 10160
rect 90786 10104 90791 10160
rect 79869 10102 90791 10104
rect 79869 10099 79935 10102
rect 90725 10099 90791 10102
rect 23565 10026 23631 10029
rect 13770 10024 23631 10026
rect 13770 9968 23570 10024
rect 23626 9968 23631 10024
rect 13770 9966 23631 9968
rect 23565 9963 23631 9966
rect 61469 10026 61535 10029
rect 64045 10026 64111 10029
rect 61469 10024 64111 10026
rect 61469 9968 61474 10024
rect 61530 9968 64050 10024
rect 64106 9968 64111 10024
rect 61469 9966 64111 9968
rect 61469 9963 61535 9966
rect 64045 9963 64111 9966
rect 18944 9824 19264 9825
rect 18944 9760 18952 9824
rect 19016 9760 19032 9824
rect 19096 9760 19112 9824
rect 19176 9760 19192 9824
rect 19256 9760 19264 9824
rect 18944 9759 19264 9760
rect 54944 9824 55264 9825
rect 54944 9760 54952 9824
rect 55016 9760 55032 9824
rect 55096 9760 55112 9824
rect 55176 9760 55192 9824
rect 55256 9760 55264 9824
rect 54944 9759 55264 9760
rect 90944 9824 91264 9825
rect 90944 9760 90952 9824
rect 91016 9760 91032 9824
rect 91096 9760 91112 9824
rect 91176 9760 91192 9824
rect 91256 9760 91264 9824
rect 90944 9759 91264 9760
rect 35157 9754 35223 9757
rect 43805 9754 43871 9757
rect 35157 9752 43871 9754
rect 35157 9696 35162 9752
rect 35218 9696 43810 9752
rect 43866 9696 43871 9752
rect 35157 9694 43871 9696
rect 35157 9691 35223 9694
rect 43805 9691 43871 9694
rect 75177 9754 75243 9757
rect 84285 9754 84351 9757
rect 75177 9752 84351 9754
rect 75177 9696 75182 9752
rect 75238 9696 84290 9752
rect 84346 9696 84351 9752
rect 75177 9694 84351 9696
rect 75177 9691 75243 9694
rect 84285 9691 84351 9694
rect 61837 9482 61903 9485
rect 42750 9480 61903 9482
rect 42750 9424 61842 9480
rect 61898 9424 61903 9480
rect 42750 9422 61903 9424
rect 39941 9346 40007 9349
rect 42750 9346 42810 9422
rect 61837 9419 61903 9422
rect 88241 9482 88307 9485
rect 104525 9482 104591 9485
rect 88241 9480 104591 9482
rect 88241 9424 88246 9480
rect 88302 9424 104530 9480
rect 104586 9424 104591 9480
rect 88241 9422 104591 9424
rect 88241 9419 88307 9422
rect 104525 9419 104591 9422
rect 39941 9344 42810 9346
rect 39941 9288 39946 9344
rect 40002 9288 42810 9344
rect 39941 9286 42810 9288
rect 39941 9283 40007 9286
rect 36944 9280 37264 9281
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 9215 37264 9216
rect 72944 9280 73264 9281
rect 72944 9216 72952 9280
rect 73016 9216 73032 9280
rect 73096 9216 73112 9280
rect 73176 9216 73192 9280
rect 73256 9216 73264 9280
rect 72944 9215 73264 9216
rect 1485 9210 1551 9213
rect 11421 9210 11487 9213
rect 1485 9208 11487 9210
rect 1485 9152 1490 9208
rect 1546 9152 11426 9208
rect 11482 9152 11487 9208
rect 1485 9150 11487 9152
rect 1485 9147 1551 9150
rect 11421 9147 11487 9150
rect 23197 9074 23263 9077
rect 36169 9074 36235 9077
rect 23197 9072 36235 9074
rect 23197 9016 23202 9072
rect 23258 9016 36174 9072
rect 36230 9016 36235 9072
rect 23197 9014 36235 9016
rect 23197 9011 23263 9014
rect 36169 9011 36235 9014
rect 105 8938 171 8941
rect 15285 8938 15351 8941
rect 105 8936 15351 8938
rect 105 8880 110 8936
rect 166 8880 15290 8936
rect 15346 8880 15351 8936
rect 105 8878 15351 8880
rect 105 8875 171 8878
rect 15285 8875 15351 8878
rect 39757 8938 39823 8941
rect 75453 8938 75519 8941
rect 39757 8936 75519 8938
rect 39757 8880 39762 8936
rect 39818 8880 75458 8936
rect 75514 8880 75519 8936
rect 39757 8878 75519 8880
rect 39757 8875 39823 8878
rect 75453 8875 75519 8878
rect 18944 8736 19264 8737
rect 18944 8672 18952 8736
rect 19016 8672 19032 8736
rect 19096 8672 19112 8736
rect 19176 8672 19192 8736
rect 19256 8672 19264 8736
rect 18944 8671 19264 8672
rect 54944 8736 55264 8737
rect 54944 8672 54952 8736
rect 55016 8672 55032 8736
rect 55096 8672 55112 8736
rect 55176 8672 55192 8736
rect 55256 8672 55264 8736
rect 54944 8671 55264 8672
rect 90944 8736 91264 8737
rect 90944 8672 90952 8736
rect 91016 8672 91032 8736
rect 91096 8672 91112 8736
rect 91176 8672 91192 8736
rect 91256 8672 91264 8736
rect 90944 8671 91264 8672
rect 21265 8530 21331 8533
rect 32489 8530 32555 8533
rect 21265 8528 32555 8530
rect 21265 8472 21270 8528
rect 21326 8472 32494 8528
rect 32550 8472 32555 8528
rect 21265 8470 32555 8472
rect 21265 8467 21331 8470
rect 32489 8467 32555 8470
rect 105 8394 171 8397
rect 9121 8394 9187 8397
rect 21909 8394 21975 8397
rect 35433 8394 35499 8397
rect 87873 8394 87939 8397
rect 105 8392 9690 8394
rect 105 8336 110 8392
rect 166 8336 9126 8392
rect 9182 8336 9690 8392
rect 105 8334 9690 8336
rect 105 8331 171 8334
rect 9121 8331 9187 8334
rect 9630 8258 9690 8334
rect 21909 8392 35499 8394
rect 21909 8336 21914 8392
rect 21970 8336 35438 8392
rect 35494 8336 35499 8392
rect 21909 8334 35499 8336
rect 21909 8331 21975 8334
rect 35433 8331 35499 8334
rect 42750 8392 87939 8394
rect 42750 8336 87878 8392
rect 87934 8336 87939 8392
rect 42750 8334 87939 8336
rect 10777 8258 10843 8261
rect 9630 8256 10843 8258
rect 9630 8200 10782 8256
rect 10838 8200 10843 8256
rect 9630 8198 10843 8200
rect 10777 8195 10843 8198
rect 23657 8258 23723 8261
rect 36813 8258 36879 8261
rect 23657 8256 36879 8258
rect 23657 8200 23662 8256
rect 23718 8200 36818 8256
rect 36874 8200 36879 8256
rect 23657 8198 36879 8200
rect 23657 8195 23723 8198
rect 36813 8195 36879 8198
rect 40033 8258 40099 8261
rect 42750 8258 42810 8334
rect 87873 8331 87939 8334
rect 40033 8256 42810 8258
rect 40033 8200 40038 8256
rect 40094 8200 42810 8256
rect 40033 8198 42810 8200
rect 66253 8258 66319 8261
rect 71865 8258 71931 8261
rect 66253 8256 71931 8258
rect 66253 8200 66258 8256
rect 66314 8200 71870 8256
rect 71926 8200 71931 8256
rect 66253 8198 71931 8200
rect 40033 8195 40099 8198
rect 66253 8195 66319 8198
rect 71865 8195 71931 8198
rect 88701 8258 88767 8261
rect 101305 8258 101371 8261
rect 88701 8256 101371 8258
rect 88701 8200 88706 8256
rect 88762 8200 101310 8256
rect 101366 8200 101371 8256
rect 88701 8198 101371 8200
rect 88701 8195 88767 8198
rect 101305 8195 101371 8198
rect 36944 8192 37264 8193
rect 0 8120 480 8152
rect 36944 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37264 8192
rect 36944 8127 37264 8128
rect 72944 8192 73264 8193
rect 72944 8128 72952 8192
rect 73016 8128 73032 8192
rect 73096 8128 73112 8192
rect 73176 8128 73192 8192
rect 73256 8128 73264 8192
rect 72944 8127 73264 8128
rect 0 8064 110 8120
rect 166 8064 480 8120
rect 0 8032 480 8064
rect 19793 8122 19859 8125
rect 32121 8122 32187 8125
rect 19793 8120 32187 8122
rect 19793 8064 19798 8120
rect 19854 8064 32126 8120
rect 32182 8064 32187 8120
rect 19793 8062 32187 8064
rect 19793 8059 19859 8062
rect 32121 8059 32187 8062
rect 23105 7986 23171 7989
rect 36353 7986 36419 7989
rect 23105 7984 36419 7986
rect 23105 7928 23110 7984
rect 23166 7928 36358 7984
rect 36414 7928 36419 7984
rect 23105 7926 36419 7928
rect 23105 7923 23171 7926
rect 36353 7923 36419 7926
rect 18944 7648 19264 7649
rect 18944 7584 18952 7648
rect 19016 7584 19032 7648
rect 19096 7584 19112 7648
rect 19176 7584 19192 7648
rect 19256 7584 19264 7648
rect 18944 7583 19264 7584
rect 54944 7648 55264 7649
rect 54944 7584 54952 7648
rect 55016 7584 55032 7648
rect 55096 7584 55112 7648
rect 55176 7584 55192 7648
rect 55256 7584 55264 7648
rect 54944 7583 55264 7584
rect 90944 7648 91264 7649
rect 90944 7584 90952 7648
rect 91016 7584 91032 7648
rect 91096 7584 91112 7648
rect 91176 7584 91192 7648
rect 91256 7584 91264 7648
rect 90944 7583 91264 7584
rect 36944 7104 37264 7105
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 7039 37264 7040
rect 72944 7104 73264 7105
rect 72944 7040 72952 7104
rect 73016 7040 73032 7104
rect 73096 7040 73112 7104
rect 73176 7040 73192 7104
rect 73256 7040 73264 7104
rect 72944 7039 73264 7040
rect 39297 6898 39363 6901
rect 46933 6898 46999 6901
rect 39297 6896 46999 6898
rect 39297 6840 39302 6896
rect 39358 6840 46938 6896
rect 46994 6840 46999 6896
rect 39297 6838 46999 6840
rect 39297 6835 39363 6838
rect 46933 6835 46999 6838
rect 18944 6560 19264 6561
rect 18944 6496 18952 6560
rect 19016 6496 19032 6560
rect 19096 6496 19112 6560
rect 19176 6496 19192 6560
rect 19256 6496 19264 6560
rect 18944 6495 19264 6496
rect 54944 6560 55264 6561
rect 54944 6496 54952 6560
rect 55016 6496 55032 6560
rect 55096 6496 55112 6560
rect 55176 6496 55192 6560
rect 55256 6496 55264 6560
rect 54944 6495 55264 6496
rect 90944 6560 91264 6561
rect 90944 6496 90952 6560
rect 91016 6496 91032 6560
rect 91096 6496 91112 6560
rect 91176 6496 91192 6560
rect 91256 6496 91264 6560
rect 90944 6495 91264 6496
rect 9489 6354 9555 6357
rect 62 6352 9555 6354
rect 62 6296 9494 6352
rect 9550 6296 9555 6352
rect 62 6294 9555 6296
rect 62 5840 122 6294
rect 9489 6291 9555 6294
rect 52361 6218 52427 6221
rect 60825 6218 60891 6221
rect 52361 6216 60891 6218
rect 52361 6160 52366 6216
rect 52422 6160 60830 6216
rect 60886 6160 60891 6216
rect 52361 6158 60891 6160
rect 52361 6155 52427 6158
rect 60825 6155 60891 6158
rect 36944 6016 37264 6017
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 5951 37264 5952
rect 72944 6016 73264 6017
rect 72944 5952 72952 6016
rect 73016 5952 73032 6016
rect 73096 5952 73112 6016
rect 73176 5952 73192 6016
rect 73256 5952 73264 6016
rect 72944 5951 73264 5952
rect 0 5720 480 5840
rect 18944 5472 19264 5473
rect 18944 5408 18952 5472
rect 19016 5408 19032 5472
rect 19096 5408 19112 5472
rect 19176 5408 19192 5472
rect 19256 5408 19264 5472
rect 18944 5407 19264 5408
rect 54944 5472 55264 5473
rect 54944 5408 54952 5472
rect 55016 5408 55032 5472
rect 55096 5408 55112 5472
rect 55176 5408 55192 5472
rect 55256 5408 55264 5472
rect 54944 5407 55264 5408
rect 90944 5472 91264 5473
rect 90944 5408 90952 5472
rect 91016 5408 91032 5472
rect 91096 5408 91112 5472
rect 91176 5408 91192 5472
rect 91256 5408 91264 5472
rect 90944 5407 91264 5408
rect 36944 4928 37264 4929
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 4863 37264 4864
rect 72944 4928 73264 4929
rect 72944 4864 72952 4928
rect 73016 4864 73032 4928
rect 73096 4864 73112 4928
rect 73176 4864 73192 4928
rect 73256 4864 73264 4928
rect 72944 4863 73264 4864
rect 26601 4858 26667 4861
rect 33777 4858 33843 4861
rect 26601 4856 33843 4858
rect 26601 4800 26606 4856
rect 26662 4800 33782 4856
rect 33838 4800 33843 4856
rect 26601 4798 33843 4800
rect 26601 4795 26667 4798
rect 33777 4795 33843 4798
rect 18944 4384 19264 4385
rect 18944 4320 18952 4384
rect 19016 4320 19032 4384
rect 19096 4320 19112 4384
rect 19176 4320 19192 4384
rect 19256 4320 19264 4384
rect 18944 4319 19264 4320
rect 54944 4384 55264 4385
rect 54944 4320 54952 4384
rect 55016 4320 55032 4384
rect 55096 4320 55112 4384
rect 55176 4320 55192 4384
rect 55256 4320 55264 4384
rect 54944 4319 55264 4320
rect 90944 4384 91264 4385
rect 90944 4320 90952 4384
rect 91016 4320 91032 4384
rect 91096 4320 91112 4384
rect 91176 4320 91192 4384
rect 91256 4320 91264 4384
rect 90944 4319 91264 4320
rect 36944 3840 37264 3841
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 3775 37264 3776
rect 72944 3840 73264 3841
rect 72944 3776 72952 3840
rect 73016 3776 73032 3840
rect 73096 3776 73112 3840
rect 73176 3776 73192 3840
rect 73256 3776 73264 3840
rect 72944 3775 73264 3776
rect 0 3408 480 3528
rect 18944 3296 19264 3297
rect 18944 3232 18952 3296
rect 19016 3232 19032 3296
rect 19096 3232 19112 3296
rect 19176 3232 19192 3296
rect 19256 3232 19264 3296
rect 18944 3231 19264 3232
rect 54944 3296 55264 3297
rect 54944 3232 54952 3296
rect 55016 3232 55032 3296
rect 55096 3232 55112 3296
rect 55176 3232 55192 3296
rect 55256 3232 55264 3296
rect 54944 3231 55264 3232
rect 90944 3296 91264 3297
rect 90944 3232 90952 3296
rect 91016 3232 91032 3296
rect 91096 3232 91112 3296
rect 91176 3232 91192 3296
rect 91256 3232 91264 3296
rect 90944 3231 91264 3232
rect 12709 2818 12775 2821
rect 19885 2818 19951 2821
rect 12709 2816 19951 2818
rect 12709 2760 12714 2816
rect 12770 2760 19890 2816
rect 19946 2760 19951 2816
rect 12709 2758 19951 2760
rect 12709 2755 12775 2758
rect 19885 2755 19951 2758
rect 78581 2818 78647 2821
rect 87413 2818 87479 2821
rect 78581 2816 87479 2818
rect 78581 2760 78586 2816
rect 78642 2760 87418 2816
rect 87474 2760 87479 2816
rect 78581 2758 87479 2760
rect 78581 2755 78647 2758
rect 87413 2755 87479 2758
rect 36944 2752 37264 2753
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2687 37264 2688
rect 72944 2752 73264 2753
rect 72944 2688 72952 2752
rect 73016 2688 73032 2752
rect 73096 2688 73112 2752
rect 73176 2688 73192 2752
rect 73256 2688 73264 2752
rect 72944 2687 73264 2688
rect 18944 2208 19264 2209
rect 18944 2144 18952 2208
rect 19016 2144 19032 2208
rect 19096 2144 19112 2208
rect 19176 2144 19192 2208
rect 19256 2144 19264 2208
rect 18944 2143 19264 2144
rect 54944 2208 55264 2209
rect 54944 2144 54952 2208
rect 55016 2144 55032 2208
rect 55096 2144 55112 2208
rect 55176 2144 55192 2208
rect 55256 2144 55264 2208
rect 54944 2143 55264 2144
rect 90944 2208 91264 2209
rect 90944 2144 90952 2208
rect 91016 2144 91032 2208
rect 91096 2144 91112 2208
rect 91176 2144 91192 2208
rect 91256 2144 91264 2208
rect 90944 2143 91264 2144
rect 54 1396 60 1460
rect 124 1458 130 1460
rect 124 1398 9690 1458
rect 124 1396 130 1398
rect 9630 1322 9690 1398
rect 18321 1322 18387 1325
rect 9630 1320 18387 1322
rect 9630 1264 18326 1320
rect 18382 1264 18387 1320
rect 9630 1262 18387 1264
rect 18321 1259 18387 1262
rect 0 1188 480 1216
rect 0 1124 60 1188
rect 124 1124 480 1188
rect 0 1096 480 1124
<< via3 >>
rect 36952 11452 37016 11456
rect 36952 11396 36956 11452
rect 36956 11396 37012 11452
rect 37012 11396 37016 11452
rect 36952 11392 37016 11396
rect 37032 11452 37096 11456
rect 37032 11396 37036 11452
rect 37036 11396 37092 11452
rect 37092 11396 37096 11452
rect 37032 11392 37096 11396
rect 37112 11452 37176 11456
rect 37112 11396 37116 11452
rect 37116 11396 37172 11452
rect 37172 11396 37176 11452
rect 37112 11392 37176 11396
rect 37192 11452 37256 11456
rect 37192 11396 37196 11452
rect 37196 11396 37252 11452
rect 37252 11396 37256 11452
rect 37192 11392 37256 11396
rect 72952 11452 73016 11456
rect 72952 11396 72956 11452
rect 72956 11396 73012 11452
rect 73012 11396 73016 11452
rect 72952 11392 73016 11396
rect 73032 11452 73096 11456
rect 73032 11396 73036 11452
rect 73036 11396 73092 11452
rect 73092 11396 73096 11452
rect 73032 11392 73096 11396
rect 73112 11452 73176 11456
rect 73112 11396 73116 11452
rect 73116 11396 73172 11452
rect 73172 11396 73176 11452
rect 73112 11392 73176 11396
rect 73192 11452 73256 11456
rect 73192 11396 73196 11452
rect 73196 11396 73252 11452
rect 73252 11396 73256 11452
rect 73192 11392 73256 11396
rect 18952 10908 19016 10912
rect 18952 10852 18956 10908
rect 18956 10852 19012 10908
rect 19012 10852 19016 10908
rect 18952 10848 19016 10852
rect 19032 10908 19096 10912
rect 19032 10852 19036 10908
rect 19036 10852 19092 10908
rect 19092 10852 19096 10908
rect 19032 10848 19096 10852
rect 19112 10908 19176 10912
rect 19112 10852 19116 10908
rect 19116 10852 19172 10908
rect 19172 10852 19176 10908
rect 19112 10848 19176 10852
rect 19192 10908 19256 10912
rect 19192 10852 19196 10908
rect 19196 10852 19252 10908
rect 19252 10852 19256 10908
rect 19192 10848 19256 10852
rect 54952 10908 55016 10912
rect 54952 10852 54956 10908
rect 54956 10852 55012 10908
rect 55012 10852 55016 10908
rect 54952 10848 55016 10852
rect 55032 10908 55096 10912
rect 55032 10852 55036 10908
rect 55036 10852 55092 10908
rect 55092 10852 55096 10908
rect 55032 10848 55096 10852
rect 55112 10908 55176 10912
rect 55112 10852 55116 10908
rect 55116 10852 55172 10908
rect 55172 10852 55176 10908
rect 55112 10848 55176 10852
rect 55192 10908 55256 10912
rect 55192 10852 55196 10908
rect 55196 10852 55252 10908
rect 55252 10852 55256 10908
rect 55192 10848 55256 10852
rect 90952 10908 91016 10912
rect 90952 10852 90956 10908
rect 90956 10852 91012 10908
rect 91012 10852 91016 10908
rect 90952 10848 91016 10852
rect 91032 10908 91096 10912
rect 91032 10852 91036 10908
rect 91036 10852 91092 10908
rect 91092 10852 91096 10908
rect 91032 10848 91096 10852
rect 91112 10908 91176 10912
rect 91112 10852 91116 10908
rect 91116 10852 91172 10908
rect 91172 10852 91176 10908
rect 91112 10848 91176 10852
rect 91192 10908 91256 10912
rect 91192 10852 91196 10908
rect 91196 10852 91252 10908
rect 91252 10852 91256 10908
rect 91192 10848 91256 10852
rect 36952 10364 37016 10368
rect 36952 10308 36956 10364
rect 36956 10308 37012 10364
rect 37012 10308 37016 10364
rect 36952 10304 37016 10308
rect 37032 10364 37096 10368
rect 37032 10308 37036 10364
rect 37036 10308 37092 10364
rect 37092 10308 37096 10364
rect 37032 10304 37096 10308
rect 37112 10364 37176 10368
rect 37112 10308 37116 10364
rect 37116 10308 37172 10364
rect 37172 10308 37176 10364
rect 37112 10304 37176 10308
rect 37192 10364 37256 10368
rect 37192 10308 37196 10364
rect 37196 10308 37252 10364
rect 37252 10308 37256 10364
rect 37192 10304 37256 10308
rect 72952 10364 73016 10368
rect 72952 10308 72956 10364
rect 72956 10308 73012 10364
rect 73012 10308 73016 10364
rect 72952 10304 73016 10308
rect 73032 10364 73096 10368
rect 73032 10308 73036 10364
rect 73036 10308 73092 10364
rect 73092 10308 73096 10364
rect 73032 10304 73096 10308
rect 73112 10364 73176 10368
rect 73112 10308 73116 10364
rect 73116 10308 73172 10364
rect 73172 10308 73176 10364
rect 73112 10304 73176 10308
rect 73192 10364 73256 10368
rect 73192 10308 73196 10364
rect 73196 10308 73252 10364
rect 73252 10308 73256 10364
rect 73192 10304 73256 10308
rect 18952 9820 19016 9824
rect 18952 9764 18956 9820
rect 18956 9764 19012 9820
rect 19012 9764 19016 9820
rect 18952 9760 19016 9764
rect 19032 9820 19096 9824
rect 19032 9764 19036 9820
rect 19036 9764 19092 9820
rect 19092 9764 19096 9820
rect 19032 9760 19096 9764
rect 19112 9820 19176 9824
rect 19112 9764 19116 9820
rect 19116 9764 19172 9820
rect 19172 9764 19176 9820
rect 19112 9760 19176 9764
rect 19192 9820 19256 9824
rect 19192 9764 19196 9820
rect 19196 9764 19252 9820
rect 19252 9764 19256 9820
rect 19192 9760 19256 9764
rect 54952 9820 55016 9824
rect 54952 9764 54956 9820
rect 54956 9764 55012 9820
rect 55012 9764 55016 9820
rect 54952 9760 55016 9764
rect 55032 9820 55096 9824
rect 55032 9764 55036 9820
rect 55036 9764 55092 9820
rect 55092 9764 55096 9820
rect 55032 9760 55096 9764
rect 55112 9820 55176 9824
rect 55112 9764 55116 9820
rect 55116 9764 55172 9820
rect 55172 9764 55176 9820
rect 55112 9760 55176 9764
rect 55192 9820 55256 9824
rect 55192 9764 55196 9820
rect 55196 9764 55252 9820
rect 55252 9764 55256 9820
rect 55192 9760 55256 9764
rect 90952 9820 91016 9824
rect 90952 9764 90956 9820
rect 90956 9764 91012 9820
rect 91012 9764 91016 9820
rect 90952 9760 91016 9764
rect 91032 9820 91096 9824
rect 91032 9764 91036 9820
rect 91036 9764 91092 9820
rect 91092 9764 91096 9820
rect 91032 9760 91096 9764
rect 91112 9820 91176 9824
rect 91112 9764 91116 9820
rect 91116 9764 91172 9820
rect 91172 9764 91176 9820
rect 91112 9760 91176 9764
rect 91192 9820 91256 9824
rect 91192 9764 91196 9820
rect 91196 9764 91252 9820
rect 91252 9764 91256 9820
rect 91192 9760 91256 9764
rect 36952 9276 37016 9280
rect 36952 9220 36956 9276
rect 36956 9220 37012 9276
rect 37012 9220 37016 9276
rect 36952 9216 37016 9220
rect 37032 9276 37096 9280
rect 37032 9220 37036 9276
rect 37036 9220 37092 9276
rect 37092 9220 37096 9276
rect 37032 9216 37096 9220
rect 37112 9276 37176 9280
rect 37112 9220 37116 9276
rect 37116 9220 37172 9276
rect 37172 9220 37176 9276
rect 37112 9216 37176 9220
rect 37192 9276 37256 9280
rect 37192 9220 37196 9276
rect 37196 9220 37252 9276
rect 37252 9220 37256 9276
rect 37192 9216 37256 9220
rect 72952 9276 73016 9280
rect 72952 9220 72956 9276
rect 72956 9220 73012 9276
rect 73012 9220 73016 9276
rect 72952 9216 73016 9220
rect 73032 9276 73096 9280
rect 73032 9220 73036 9276
rect 73036 9220 73092 9276
rect 73092 9220 73096 9276
rect 73032 9216 73096 9220
rect 73112 9276 73176 9280
rect 73112 9220 73116 9276
rect 73116 9220 73172 9276
rect 73172 9220 73176 9276
rect 73112 9216 73176 9220
rect 73192 9276 73256 9280
rect 73192 9220 73196 9276
rect 73196 9220 73252 9276
rect 73252 9220 73256 9276
rect 73192 9216 73256 9220
rect 18952 8732 19016 8736
rect 18952 8676 18956 8732
rect 18956 8676 19012 8732
rect 19012 8676 19016 8732
rect 18952 8672 19016 8676
rect 19032 8732 19096 8736
rect 19032 8676 19036 8732
rect 19036 8676 19092 8732
rect 19092 8676 19096 8732
rect 19032 8672 19096 8676
rect 19112 8732 19176 8736
rect 19112 8676 19116 8732
rect 19116 8676 19172 8732
rect 19172 8676 19176 8732
rect 19112 8672 19176 8676
rect 19192 8732 19256 8736
rect 19192 8676 19196 8732
rect 19196 8676 19252 8732
rect 19252 8676 19256 8732
rect 19192 8672 19256 8676
rect 54952 8732 55016 8736
rect 54952 8676 54956 8732
rect 54956 8676 55012 8732
rect 55012 8676 55016 8732
rect 54952 8672 55016 8676
rect 55032 8732 55096 8736
rect 55032 8676 55036 8732
rect 55036 8676 55092 8732
rect 55092 8676 55096 8732
rect 55032 8672 55096 8676
rect 55112 8732 55176 8736
rect 55112 8676 55116 8732
rect 55116 8676 55172 8732
rect 55172 8676 55176 8732
rect 55112 8672 55176 8676
rect 55192 8732 55256 8736
rect 55192 8676 55196 8732
rect 55196 8676 55252 8732
rect 55252 8676 55256 8732
rect 55192 8672 55256 8676
rect 90952 8732 91016 8736
rect 90952 8676 90956 8732
rect 90956 8676 91012 8732
rect 91012 8676 91016 8732
rect 90952 8672 91016 8676
rect 91032 8732 91096 8736
rect 91032 8676 91036 8732
rect 91036 8676 91092 8732
rect 91092 8676 91096 8732
rect 91032 8672 91096 8676
rect 91112 8732 91176 8736
rect 91112 8676 91116 8732
rect 91116 8676 91172 8732
rect 91172 8676 91176 8732
rect 91112 8672 91176 8676
rect 91192 8732 91256 8736
rect 91192 8676 91196 8732
rect 91196 8676 91252 8732
rect 91252 8676 91256 8732
rect 91192 8672 91256 8676
rect 36952 8188 37016 8192
rect 36952 8132 36956 8188
rect 36956 8132 37012 8188
rect 37012 8132 37016 8188
rect 36952 8128 37016 8132
rect 37032 8188 37096 8192
rect 37032 8132 37036 8188
rect 37036 8132 37092 8188
rect 37092 8132 37096 8188
rect 37032 8128 37096 8132
rect 37112 8188 37176 8192
rect 37112 8132 37116 8188
rect 37116 8132 37172 8188
rect 37172 8132 37176 8188
rect 37112 8128 37176 8132
rect 37192 8188 37256 8192
rect 37192 8132 37196 8188
rect 37196 8132 37252 8188
rect 37252 8132 37256 8188
rect 37192 8128 37256 8132
rect 72952 8188 73016 8192
rect 72952 8132 72956 8188
rect 72956 8132 73012 8188
rect 73012 8132 73016 8188
rect 72952 8128 73016 8132
rect 73032 8188 73096 8192
rect 73032 8132 73036 8188
rect 73036 8132 73092 8188
rect 73092 8132 73096 8188
rect 73032 8128 73096 8132
rect 73112 8188 73176 8192
rect 73112 8132 73116 8188
rect 73116 8132 73172 8188
rect 73172 8132 73176 8188
rect 73112 8128 73176 8132
rect 73192 8188 73256 8192
rect 73192 8132 73196 8188
rect 73196 8132 73252 8188
rect 73252 8132 73256 8188
rect 73192 8128 73256 8132
rect 18952 7644 19016 7648
rect 18952 7588 18956 7644
rect 18956 7588 19012 7644
rect 19012 7588 19016 7644
rect 18952 7584 19016 7588
rect 19032 7644 19096 7648
rect 19032 7588 19036 7644
rect 19036 7588 19092 7644
rect 19092 7588 19096 7644
rect 19032 7584 19096 7588
rect 19112 7644 19176 7648
rect 19112 7588 19116 7644
rect 19116 7588 19172 7644
rect 19172 7588 19176 7644
rect 19112 7584 19176 7588
rect 19192 7644 19256 7648
rect 19192 7588 19196 7644
rect 19196 7588 19252 7644
rect 19252 7588 19256 7644
rect 19192 7584 19256 7588
rect 54952 7644 55016 7648
rect 54952 7588 54956 7644
rect 54956 7588 55012 7644
rect 55012 7588 55016 7644
rect 54952 7584 55016 7588
rect 55032 7644 55096 7648
rect 55032 7588 55036 7644
rect 55036 7588 55092 7644
rect 55092 7588 55096 7644
rect 55032 7584 55096 7588
rect 55112 7644 55176 7648
rect 55112 7588 55116 7644
rect 55116 7588 55172 7644
rect 55172 7588 55176 7644
rect 55112 7584 55176 7588
rect 55192 7644 55256 7648
rect 55192 7588 55196 7644
rect 55196 7588 55252 7644
rect 55252 7588 55256 7644
rect 55192 7584 55256 7588
rect 90952 7644 91016 7648
rect 90952 7588 90956 7644
rect 90956 7588 91012 7644
rect 91012 7588 91016 7644
rect 90952 7584 91016 7588
rect 91032 7644 91096 7648
rect 91032 7588 91036 7644
rect 91036 7588 91092 7644
rect 91092 7588 91096 7644
rect 91032 7584 91096 7588
rect 91112 7644 91176 7648
rect 91112 7588 91116 7644
rect 91116 7588 91172 7644
rect 91172 7588 91176 7644
rect 91112 7584 91176 7588
rect 91192 7644 91256 7648
rect 91192 7588 91196 7644
rect 91196 7588 91252 7644
rect 91252 7588 91256 7644
rect 91192 7584 91256 7588
rect 36952 7100 37016 7104
rect 36952 7044 36956 7100
rect 36956 7044 37012 7100
rect 37012 7044 37016 7100
rect 36952 7040 37016 7044
rect 37032 7100 37096 7104
rect 37032 7044 37036 7100
rect 37036 7044 37092 7100
rect 37092 7044 37096 7100
rect 37032 7040 37096 7044
rect 37112 7100 37176 7104
rect 37112 7044 37116 7100
rect 37116 7044 37172 7100
rect 37172 7044 37176 7100
rect 37112 7040 37176 7044
rect 37192 7100 37256 7104
rect 37192 7044 37196 7100
rect 37196 7044 37252 7100
rect 37252 7044 37256 7100
rect 37192 7040 37256 7044
rect 72952 7100 73016 7104
rect 72952 7044 72956 7100
rect 72956 7044 73012 7100
rect 73012 7044 73016 7100
rect 72952 7040 73016 7044
rect 73032 7100 73096 7104
rect 73032 7044 73036 7100
rect 73036 7044 73092 7100
rect 73092 7044 73096 7100
rect 73032 7040 73096 7044
rect 73112 7100 73176 7104
rect 73112 7044 73116 7100
rect 73116 7044 73172 7100
rect 73172 7044 73176 7100
rect 73112 7040 73176 7044
rect 73192 7100 73256 7104
rect 73192 7044 73196 7100
rect 73196 7044 73252 7100
rect 73252 7044 73256 7100
rect 73192 7040 73256 7044
rect 18952 6556 19016 6560
rect 18952 6500 18956 6556
rect 18956 6500 19012 6556
rect 19012 6500 19016 6556
rect 18952 6496 19016 6500
rect 19032 6556 19096 6560
rect 19032 6500 19036 6556
rect 19036 6500 19092 6556
rect 19092 6500 19096 6556
rect 19032 6496 19096 6500
rect 19112 6556 19176 6560
rect 19112 6500 19116 6556
rect 19116 6500 19172 6556
rect 19172 6500 19176 6556
rect 19112 6496 19176 6500
rect 19192 6556 19256 6560
rect 19192 6500 19196 6556
rect 19196 6500 19252 6556
rect 19252 6500 19256 6556
rect 19192 6496 19256 6500
rect 54952 6556 55016 6560
rect 54952 6500 54956 6556
rect 54956 6500 55012 6556
rect 55012 6500 55016 6556
rect 54952 6496 55016 6500
rect 55032 6556 55096 6560
rect 55032 6500 55036 6556
rect 55036 6500 55092 6556
rect 55092 6500 55096 6556
rect 55032 6496 55096 6500
rect 55112 6556 55176 6560
rect 55112 6500 55116 6556
rect 55116 6500 55172 6556
rect 55172 6500 55176 6556
rect 55112 6496 55176 6500
rect 55192 6556 55256 6560
rect 55192 6500 55196 6556
rect 55196 6500 55252 6556
rect 55252 6500 55256 6556
rect 55192 6496 55256 6500
rect 90952 6556 91016 6560
rect 90952 6500 90956 6556
rect 90956 6500 91012 6556
rect 91012 6500 91016 6556
rect 90952 6496 91016 6500
rect 91032 6556 91096 6560
rect 91032 6500 91036 6556
rect 91036 6500 91092 6556
rect 91092 6500 91096 6556
rect 91032 6496 91096 6500
rect 91112 6556 91176 6560
rect 91112 6500 91116 6556
rect 91116 6500 91172 6556
rect 91172 6500 91176 6556
rect 91112 6496 91176 6500
rect 91192 6556 91256 6560
rect 91192 6500 91196 6556
rect 91196 6500 91252 6556
rect 91252 6500 91256 6556
rect 91192 6496 91256 6500
rect 36952 6012 37016 6016
rect 36952 5956 36956 6012
rect 36956 5956 37012 6012
rect 37012 5956 37016 6012
rect 36952 5952 37016 5956
rect 37032 6012 37096 6016
rect 37032 5956 37036 6012
rect 37036 5956 37092 6012
rect 37092 5956 37096 6012
rect 37032 5952 37096 5956
rect 37112 6012 37176 6016
rect 37112 5956 37116 6012
rect 37116 5956 37172 6012
rect 37172 5956 37176 6012
rect 37112 5952 37176 5956
rect 37192 6012 37256 6016
rect 37192 5956 37196 6012
rect 37196 5956 37252 6012
rect 37252 5956 37256 6012
rect 37192 5952 37256 5956
rect 72952 6012 73016 6016
rect 72952 5956 72956 6012
rect 72956 5956 73012 6012
rect 73012 5956 73016 6012
rect 72952 5952 73016 5956
rect 73032 6012 73096 6016
rect 73032 5956 73036 6012
rect 73036 5956 73092 6012
rect 73092 5956 73096 6012
rect 73032 5952 73096 5956
rect 73112 6012 73176 6016
rect 73112 5956 73116 6012
rect 73116 5956 73172 6012
rect 73172 5956 73176 6012
rect 73112 5952 73176 5956
rect 73192 6012 73256 6016
rect 73192 5956 73196 6012
rect 73196 5956 73252 6012
rect 73252 5956 73256 6012
rect 73192 5952 73256 5956
rect 18952 5468 19016 5472
rect 18952 5412 18956 5468
rect 18956 5412 19012 5468
rect 19012 5412 19016 5468
rect 18952 5408 19016 5412
rect 19032 5468 19096 5472
rect 19032 5412 19036 5468
rect 19036 5412 19092 5468
rect 19092 5412 19096 5468
rect 19032 5408 19096 5412
rect 19112 5468 19176 5472
rect 19112 5412 19116 5468
rect 19116 5412 19172 5468
rect 19172 5412 19176 5468
rect 19112 5408 19176 5412
rect 19192 5468 19256 5472
rect 19192 5412 19196 5468
rect 19196 5412 19252 5468
rect 19252 5412 19256 5468
rect 19192 5408 19256 5412
rect 54952 5468 55016 5472
rect 54952 5412 54956 5468
rect 54956 5412 55012 5468
rect 55012 5412 55016 5468
rect 54952 5408 55016 5412
rect 55032 5468 55096 5472
rect 55032 5412 55036 5468
rect 55036 5412 55092 5468
rect 55092 5412 55096 5468
rect 55032 5408 55096 5412
rect 55112 5468 55176 5472
rect 55112 5412 55116 5468
rect 55116 5412 55172 5468
rect 55172 5412 55176 5468
rect 55112 5408 55176 5412
rect 55192 5468 55256 5472
rect 55192 5412 55196 5468
rect 55196 5412 55252 5468
rect 55252 5412 55256 5468
rect 55192 5408 55256 5412
rect 90952 5468 91016 5472
rect 90952 5412 90956 5468
rect 90956 5412 91012 5468
rect 91012 5412 91016 5468
rect 90952 5408 91016 5412
rect 91032 5468 91096 5472
rect 91032 5412 91036 5468
rect 91036 5412 91092 5468
rect 91092 5412 91096 5468
rect 91032 5408 91096 5412
rect 91112 5468 91176 5472
rect 91112 5412 91116 5468
rect 91116 5412 91172 5468
rect 91172 5412 91176 5468
rect 91112 5408 91176 5412
rect 91192 5468 91256 5472
rect 91192 5412 91196 5468
rect 91196 5412 91252 5468
rect 91252 5412 91256 5468
rect 91192 5408 91256 5412
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 72952 4924 73016 4928
rect 72952 4868 72956 4924
rect 72956 4868 73012 4924
rect 73012 4868 73016 4924
rect 72952 4864 73016 4868
rect 73032 4924 73096 4928
rect 73032 4868 73036 4924
rect 73036 4868 73092 4924
rect 73092 4868 73096 4924
rect 73032 4864 73096 4868
rect 73112 4924 73176 4928
rect 73112 4868 73116 4924
rect 73116 4868 73172 4924
rect 73172 4868 73176 4924
rect 73112 4864 73176 4868
rect 73192 4924 73256 4928
rect 73192 4868 73196 4924
rect 73196 4868 73252 4924
rect 73252 4868 73256 4924
rect 73192 4864 73256 4868
rect 18952 4380 19016 4384
rect 18952 4324 18956 4380
rect 18956 4324 19012 4380
rect 19012 4324 19016 4380
rect 18952 4320 19016 4324
rect 19032 4380 19096 4384
rect 19032 4324 19036 4380
rect 19036 4324 19092 4380
rect 19092 4324 19096 4380
rect 19032 4320 19096 4324
rect 19112 4380 19176 4384
rect 19112 4324 19116 4380
rect 19116 4324 19172 4380
rect 19172 4324 19176 4380
rect 19112 4320 19176 4324
rect 19192 4380 19256 4384
rect 19192 4324 19196 4380
rect 19196 4324 19252 4380
rect 19252 4324 19256 4380
rect 19192 4320 19256 4324
rect 54952 4380 55016 4384
rect 54952 4324 54956 4380
rect 54956 4324 55012 4380
rect 55012 4324 55016 4380
rect 54952 4320 55016 4324
rect 55032 4380 55096 4384
rect 55032 4324 55036 4380
rect 55036 4324 55092 4380
rect 55092 4324 55096 4380
rect 55032 4320 55096 4324
rect 55112 4380 55176 4384
rect 55112 4324 55116 4380
rect 55116 4324 55172 4380
rect 55172 4324 55176 4380
rect 55112 4320 55176 4324
rect 55192 4380 55256 4384
rect 55192 4324 55196 4380
rect 55196 4324 55252 4380
rect 55252 4324 55256 4380
rect 55192 4320 55256 4324
rect 90952 4380 91016 4384
rect 90952 4324 90956 4380
rect 90956 4324 91012 4380
rect 91012 4324 91016 4380
rect 90952 4320 91016 4324
rect 91032 4380 91096 4384
rect 91032 4324 91036 4380
rect 91036 4324 91092 4380
rect 91092 4324 91096 4380
rect 91032 4320 91096 4324
rect 91112 4380 91176 4384
rect 91112 4324 91116 4380
rect 91116 4324 91172 4380
rect 91172 4324 91176 4380
rect 91112 4320 91176 4324
rect 91192 4380 91256 4384
rect 91192 4324 91196 4380
rect 91196 4324 91252 4380
rect 91252 4324 91256 4380
rect 91192 4320 91256 4324
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 72952 3836 73016 3840
rect 72952 3780 72956 3836
rect 72956 3780 73012 3836
rect 73012 3780 73016 3836
rect 72952 3776 73016 3780
rect 73032 3836 73096 3840
rect 73032 3780 73036 3836
rect 73036 3780 73092 3836
rect 73092 3780 73096 3836
rect 73032 3776 73096 3780
rect 73112 3836 73176 3840
rect 73112 3780 73116 3836
rect 73116 3780 73172 3836
rect 73172 3780 73176 3836
rect 73112 3776 73176 3780
rect 73192 3836 73256 3840
rect 73192 3780 73196 3836
rect 73196 3780 73252 3836
rect 73252 3780 73256 3836
rect 73192 3776 73256 3780
rect 18952 3292 19016 3296
rect 18952 3236 18956 3292
rect 18956 3236 19012 3292
rect 19012 3236 19016 3292
rect 18952 3232 19016 3236
rect 19032 3292 19096 3296
rect 19032 3236 19036 3292
rect 19036 3236 19092 3292
rect 19092 3236 19096 3292
rect 19032 3232 19096 3236
rect 19112 3292 19176 3296
rect 19112 3236 19116 3292
rect 19116 3236 19172 3292
rect 19172 3236 19176 3292
rect 19112 3232 19176 3236
rect 19192 3292 19256 3296
rect 19192 3236 19196 3292
rect 19196 3236 19252 3292
rect 19252 3236 19256 3292
rect 19192 3232 19256 3236
rect 54952 3292 55016 3296
rect 54952 3236 54956 3292
rect 54956 3236 55012 3292
rect 55012 3236 55016 3292
rect 54952 3232 55016 3236
rect 55032 3292 55096 3296
rect 55032 3236 55036 3292
rect 55036 3236 55092 3292
rect 55092 3236 55096 3292
rect 55032 3232 55096 3236
rect 55112 3292 55176 3296
rect 55112 3236 55116 3292
rect 55116 3236 55172 3292
rect 55172 3236 55176 3292
rect 55112 3232 55176 3236
rect 55192 3292 55256 3296
rect 55192 3236 55196 3292
rect 55196 3236 55252 3292
rect 55252 3236 55256 3292
rect 55192 3232 55256 3236
rect 90952 3292 91016 3296
rect 90952 3236 90956 3292
rect 90956 3236 91012 3292
rect 91012 3236 91016 3292
rect 90952 3232 91016 3236
rect 91032 3292 91096 3296
rect 91032 3236 91036 3292
rect 91036 3236 91092 3292
rect 91092 3236 91096 3292
rect 91032 3232 91096 3236
rect 91112 3292 91176 3296
rect 91112 3236 91116 3292
rect 91116 3236 91172 3292
rect 91172 3236 91176 3292
rect 91112 3232 91176 3236
rect 91192 3292 91256 3296
rect 91192 3236 91196 3292
rect 91196 3236 91252 3292
rect 91252 3236 91256 3292
rect 91192 3232 91256 3236
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 72952 2748 73016 2752
rect 72952 2692 72956 2748
rect 72956 2692 73012 2748
rect 73012 2692 73016 2748
rect 72952 2688 73016 2692
rect 73032 2748 73096 2752
rect 73032 2692 73036 2748
rect 73036 2692 73092 2748
rect 73092 2692 73096 2748
rect 73032 2688 73096 2692
rect 73112 2748 73176 2752
rect 73112 2692 73116 2748
rect 73116 2692 73172 2748
rect 73172 2692 73176 2748
rect 73112 2688 73176 2692
rect 73192 2748 73256 2752
rect 73192 2692 73196 2748
rect 73196 2692 73252 2748
rect 73252 2692 73256 2748
rect 73192 2688 73256 2692
rect 18952 2204 19016 2208
rect 18952 2148 18956 2204
rect 18956 2148 19012 2204
rect 19012 2148 19016 2204
rect 18952 2144 19016 2148
rect 19032 2204 19096 2208
rect 19032 2148 19036 2204
rect 19036 2148 19092 2204
rect 19092 2148 19096 2204
rect 19032 2144 19096 2148
rect 19112 2204 19176 2208
rect 19112 2148 19116 2204
rect 19116 2148 19172 2204
rect 19172 2148 19176 2204
rect 19112 2144 19176 2148
rect 19192 2204 19256 2208
rect 19192 2148 19196 2204
rect 19196 2148 19252 2204
rect 19252 2148 19256 2204
rect 19192 2144 19256 2148
rect 54952 2204 55016 2208
rect 54952 2148 54956 2204
rect 54956 2148 55012 2204
rect 55012 2148 55016 2204
rect 54952 2144 55016 2148
rect 55032 2204 55096 2208
rect 55032 2148 55036 2204
rect 55036 2148 55092 2204
rect 55092 2148 55096 2204
rect 55032 2144 55096 2148
rect 55112 2204 55176 2208
rect 55112 2148 55116 2204
rect 55116 2148 55172 2204
rect 55172 2148 55176 2204
rect 55112 2144 55176 2148
rect 55192 2204 55256 2208
rect 55192 2148 55196 2204
rect 55196 2148 55252 2204
rect 55252 2148 55256 2204
rect 55192 2144 55256 2148
rect 90952 2204 91016 2208
rect 90952 2148 90956 2204
rect 90956 2148 91012 2204
rect 91012 2148 91016 2204
rect 90952 2144 91016 2148
rect 91032 2204 91096 2208
rect 91032 2148 91036 2204
rect 91036 2148 91092 2204
rect 91092 2148 91096 2204
rect 91032 2144 91096 2148
rect 91112 2204 91176 2208
rect 91112 2148 91116 2204
rect 91116 2148 91172 2204
rect 91172 2148 91176 2204
rect 91112 2144 91176 2148
rect 91192 2204 91256 2208
rect 91192 2148 91196 2204
rect 91196 2148 91252 2204
rect 91252 2148 91256 2204
rect 91192 2144 91256 2148
rect 60 1396 124 1460
rect 60 1124 124 1188
<< metal4 >>
rect 18944 10912 19264 11472
rect 18944 10848 18952 10912
rect 19016 10848 19032 10912
rect 19096 10848 19112 10912
rect 19176 10848 19192 10912
rect 19256 10848 19264 10912
rect 18944 9824 19264 10848
rect 18944 9760 18952 9824
rect 19016 9760 19032 9824
rect 19096 9760 19112 9824
rect 19176 9760 19192 9824
rect 19256 9760 19264 9824
rect 18944 8736 19264 9760
rect 18944 8672 18952 8736
rect 19016 8672 19032 8736
rect 19096 8672 19112 8736
rect 19176 8672 19192 8736
rect 19256 8672 19264 8736
rect 18944 7648 19264 8672
rect 18944 7584 18952 7648
rect 19016 7584 19032 7648
rect 19096 7584 19112 7648
rect 19176 7584 19192 7648
rect 19256 7584 19264 7648
rect 18944 6560 19264 7584
rect 18944 6496 18952 6560
rect 19016 6496 19032 6560
rect 19096 6496 19112 6560
rect 19176 6496 19192 6560
rect 19256 6496 19264 6560
rect 18944 5472 19264 6496
rect 18944 5408 18952 5472
rect 19016 5408 19032 5472
rect 19096 5408 19112 5472
rect 19176 5408 19192 5472
rect 19256 5408 19264 5472
rect 18944 4384 19264 5408
rect 18944 4320 18952 4384
rect 19016 4320 19032 4384
rect 19096 4320 19112 4384
rect 19176 4320 19192 4384
rect 19256 4320 19264 4384
rect 18944 3296 19264 4320
rect 18944 3232 18952 3296
rect 19016 3232 19032 3296
rect 19096 3232 19112 3296
rect 19176 3232 19192 3296
rect 19256 3232 19264 3296
rect 18944 2208 19264 3232
rect 18944 2144 18952 2208
rect 19016 2144 19032 2208
rect 19096 2144 19112 2208
rect 19176 2144 19192 2208
rect 19256 2144 19264 2208
rect 18944 2128 19264 2144
rect 36944 11456 37264 11472
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 10368 37264 11392
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 9280 37264 10304
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 8192 37264 9216
rect 36944 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37264 8192
rect 36944 7104 37264 8128
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 6016 37264 7040
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 4928 37264 5952
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 2752 37264 3776
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2128 37264 2688
rect 54944 10912 55264 11472
rect 54944 10848 54952 10912
rect 55016 10848 55032 10912
rect 55096 10848 55112 10912
rect 55176 10848 55192 10912
rect 55256 10848 55264 10912
rect 54944 9824 55264 10848
rect 54944 9760 54952 9824
rect 55016 9760 55032 9824
rect 55096 9760 55112 9824
rect 55176 9760 55192 9824
rect 55256 9760 55264 9824
rect 54944 8736 55264 9760
rect 54944 8672 54952 8736
rect 55016 8672 55032 8736
rect 55096 8672 55112 8736
rect 55176 8672 55192 8736
rect 55256 8672 55264 8736
rect 54944 7648 55264 8672
rect 54944 7584 54952 7648
rect 55016 7584 55032 7648
rect 55096 7584 55112 7648
rect 55176 7584 55192 7648
rect 55256 7584 55264 7648
rect 54944 6560 55264 7584
rect 54944 6496 54952 6560
rect 55016 6496 55032 6560
rect 55096 6496 55112 6560
rect 55176 6496 55192 6560
rect 55256 6496 55264 6560
rect 54944 5472 55264 6496
rect 54944 5408 54952 5472
rect 55016 5408 55032 5472
rect 55096 5408 55112 5472
rect 55176 5408 55192 5472
rect 55256 5408 55264 5472
rect 54944 4384 55264 5408
rect 54944 4320 54952 4384
rect 55016 4320 55032 4384
rect 55096 4320 55112 4384
rect 55176 4320 55192 4384
rect 55256 4320 55264 4384
rect 54944 3296 55264 4320
rect 54944 3232 54952 3296
rect 55016 3232 55032 3296
rect 55096 3232 55112 3296
rect 55176 3232 55192 3296
rect 55256 3232 55264 3296
rect 54944 2208 55264 3232
rect 54944 2144 54952 2208
rect 55016 2144 55032 2208
rect 55096 2144 55112 2208
rect 55176 2144 55192 2208
rect 55256 2144 55264 2208
rect 54944 2128 55264 2144
rect 72944 11456 73264 11472
rect 72944 11392 72952 11456
rect 73016 11392 73032 11456
rect 73096 11392 73112 11456
rect 73176 11392 73192 11456
rect 73256 11392 73264 11456
rect 72944 10368 73264 11392
rect 72944 10304 72952 10368
rect 73016 10304 73032 10368
rect 73096 10304 73112 10368
rect 73176 10304 73192 10368
rect 73256 10304 73264 10368
rect 72944 9280 73264 10304
rect 72944 9216 72952 9280
rect 73016 9216 73032 9280
rect 73096 9216 73112 9280
rect 73176 9216 73192 9280
rect 73256 9216 73264 9280
rect 72944 8192 73264 9216
rect 72944 8128 72952 8192
rect 73016 8128 73032 8192
rect 73096 8128 73112 8192
rect 73176 8128 73192 8192
rect 73256 8128 73264 8192
rect 72944 7104 73264 8128
rect 72944 7040 72952 7104
rect 73016 7040 73032 7104
rect 73096 7040 73112 7104
rect 73176 7040 73192 7104
rect 73256 7040 73264 7104
rect 72944 6016 73264 7040
rect 72944 5952 72952 6016
rect 73016 5952 73032 6016
rect 73096 5952 73112 6016
rect 73176 5952 73192 6016
rect 73256 5952 73264 6016
rect 72944 4928 73264 5952
rect 72944 4864 72952 4928
rect 73016 4864 73032 4928
rect 73096 4864 73112 4928
rect 73176 4864 73192 4928
rect 73256 4864 73264 4928
rect 72944 3840 73264 4864
rect 72944 3776 72952 3840
rect 73016 3776 73032 3840
rect 73096 3776 73112 3840
rect 73176 3776 73192 3840
rect 73256 3776 73264 3840
rect 72944 2752 73264 3776
rect 72944 2688 72952 2752
rect 73016 2688 73032 2752
rect 73096 2688 73112 2752
rect 73176 2688 73192 2752
rect 73256 2688 73264 2752
rect 72944 2128 73264 2688
rect 90944 10912 91264 11472
rect 90944 10848 90952 10912
rect 91016 10848 91032 10912
rect 91096 10848 91112 10912
rect 91176 10848 91192 10912
rect 91256 10848 91264 10912
rect 90944 9824 91264 10848
rect 90944 9760 90952 9824
rect 91016 9760 91032 9824
rect 91096 9760 91112 9824
rect 91176 9760 91192 9824
rect 91256 9760 91264 9824
rect 90944 8736 91264 9760
rect 90944 8672 90952 8736
rect 91016 8672 91032 8736
rect 91096 8672 91112 8736
rect 91176 8672 91192 8736
rect 91256 8672 91264 8736
rect 90944 7648 91264 8672
rect 90944 7584 90952 7648
rect 91016 7584 91032 7648
rect 91096 7584 91112 7648
rect 91176 7584 91192 7648
rect 91256 7584 91264 7648
rect 90944 6560 91264 7584
rect 90944 6496 90952 6560
rect 91016 6496 91032 6560
rect 91096 6496 91112 6560
rect 91176 6496 91192 6560
rect 91256 6496 91264 6560
rect 90944 5472 91264 6496
rect 90944 5408 90952 5472
rect 91016 5408 91032 5472
rect 91096 5408 91112 5472
rect 91176 5408 91192 5472
rect 91256 5408 91264 5472
rect 90944 4384 91264 5408
rect 90944 4320 90952 4384
rect 91016 4320 91032 4384
rect 91096 4320 91112 4384
rect 91176 4320 91192 4384
rect 91256 4320 91264 4384
rect 90944 3296 91264 4320
rect 90944 3232 90952 3296
rect 91016 3232 91032 3296
rect 91096 3232 91112 3296
rect 91176 3232 91192 3296
rect 91256 3232 91264 3296
rect 90944 2208 91264 3232
rect 90944 2144 90952 2208
rect 91016 2144 91032 2208
rect 91096 2144 91112 2208
rect 91176 2144 91192 2208
rect 91256 2144 91264 2208
rect 90944 2128 91264 2144
rect 59 1460 125 1461
rect 59 1396 60 1460
rect 124 1396 125 1460
rect 59 1395 125 1396
rect 62 1189 122 1395
rect 59 1188 125 1189
rect 59 1124 60 1188
rect 124 1124 125 1188
rect 59 1123 125 1124
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_34 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_35
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_36
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_37
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_38
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_39
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_40
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_41
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_42
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_416
timestamp 1586364061
transform 1 0 39376 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_428
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_415
timestamp 1586364061
transform 1 0 39284 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_428
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_440
timestamp 1586364061
transform 1 0 41584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_447
timestamp 1586364061
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_459
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_452
timestamp 1586364061
transform 1 0 42688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_466
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_478
timestamp 1586364061
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_464
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_476
timestamp 1586364061
transform 1 0 44896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_490
timestamp 1586364061
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_521
timestamp 1586364061
transform 1 0 49036 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_528
timestamp 1586364061
transform 1 0 49680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_525
timestamp 1586364061
transform 1 0 49404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_540
timestamp 1586364061
transform 1 0 50784 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_552
timestamp 1586364061
transform 1 0 51888 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_537
timestamp 1586364061
transform 1 0 50508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_550
timestamp 1586364061
transform 1 0 51704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_559
timestamp 1586364061
transform 1 0 52532 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_562
timestamp 1586364061
transform 1 0 52808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_571
timestamp 1586364061
transform 1 0 53636 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_583
timestamp 1586364061
transform 1 0 54740 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_574
timestamp 1586364061
transform 1 0 53912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_586
timestamp 1586364061
transform 1 0 55016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 55292 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_590
timestamp 1586364061
transform 1 0 55384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_602
timestamp 1586364061
transform 1 0 56488 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_598
timestamp 1586364061
transform 1 0 56120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 58144 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_614
timestamp 1586364061
transform 1 0 57592 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_621
timestamp 1586364061
transform 1 0 58236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_611
timestamp 1586364061
transform 1 0 57316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_623
timestamp 1586364061
transform 1 0 58420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_633
timestamp 1586364061
transform 1 0 59340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_635
timestamp 1586364061
transform 1 0 59524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 60996 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_645
timestamp 1586364061
transform 1 0 60444 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_652
timestamp 1586364061
transform 1 0 61088 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_647
timestamp 1586364061
transform 1 0 60628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_659
timestamp 1586364061
transform 1 0 61732 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_664
timestamp 1586364061
transform 1 0 62192 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_676
timestamp 1586364061
transform 1 0 63296 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_672
timestamp 1586364061
transform 1 0 62928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 63848 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_683
timestamp 1586364061
transform 1 0 63940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_695
timestamp 1586364061
transform 1 0 65044 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_684
timestamp 1586364061
transform 1 0 64032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 66700 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_707
timestamp 1586364061
transform 1 0 66148 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_696
timestamp 1586364061
transform 1 0 65136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_708
timestamp 1586364061
transform 1 0 66240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_714
timestamp 1586364061
transform 1 0 66792 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_726
timestamp 1586364061
transform 1 0 67896 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_720
timestamp 1586364061
transform 1 0 67344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 69552 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 68448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_738
timestamp 1586364061
transform 1 0 69000 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_745
timestamp 1586364061
transform 1 0 69644 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_733
timestamp 1586364061
transform 1 0 68540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_745
timestamp 1586364061
transform 1 0 69644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_757
timestamp 1586364061
transform 1 0 70748 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_757
timestamp 1586364061
transform 1 0 70748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 72404 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_769
timestamp 1586364061
transform 1 0 71852 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_776
timestamp 1586364061
transform 1 0 72496 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_769
timestamp 1586364061
transform 1 0 71852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_781
timestamp 1586364061
transform 1 0 72956 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 74060 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_788
timestamp 1586364061
transform 1 0 73600 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_800
timestamp 1586364061
transform 1 0 74704 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_794
timestamp 1586364061
transform 1 0 74152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 75256 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_807
timestamp 1586364061
transform 1 0 75348 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_819
timestamp 1586364061
transform 1 0 76452 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_806
timestamp 1586364061
transform 1 0 75256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_818
timestamp 1586364061
transform 1 0 76360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 78108 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_831
timestamp 1586364061
transform 1 0 77556 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_838
timestamp 1586364061
transform 1 0 78200 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_830
timestamp 1586364061
transform 1 0 77464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 79672 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_850
timestamp 1586364061
transform 1 0 79304 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_842
timestamp 1586364061
transform 1 0 78568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_855
timestamp 1586364061
transform 1 0 79764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 80960 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_862
timestamp 1586364061
transform 1 0 80408 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_869
timestamp 1586364061
transform 1 0 81052 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_867
timestamp 1586364061
transform 1 0 80868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_881
timestamp 1586364061
transform 1 0 82156 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_879
timestamp 1586364061
transform 1 0 81972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_891
timestamp 1586364061
transform 1 0 83076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 83812 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_893
timestamp 1586364061
transform 1 0 83260 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_900
timestamp 1586364061
transform 1 0 83904 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_903
timestamp 1586364061
transform 1 0 84180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 85284 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_912
timestamp 1586364061
transform 1 0 85008 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_924
timestamp 1586364061
transform 1 0 86112 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_916
timestamp 1586364061
transform 1 0 85376 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 86664 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_931
timestamp 1586364061
transform 1 0 86756 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_943
timestamp 1586364061
transform 1 0 87860 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_928
timestamp 1586364061
transform 1 0 86480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_940
timestamp 1586364061
transform 1 0 87584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 89516 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_955
timestamp 1586364061
transform 1 0 88964 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_962
timestamp 1586364061
transform 1 0 89608 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_952
timestamp 1586364061
transform 1 0 88688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 90896 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_974
timestamp 1586364061
transform 1 0 90712 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_964
timestamp 1586364061
transform 1 0 89792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_977
timestamp 1586364061
transform 1 0 90988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 92368 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_986
timestamp 1586364061
transform 1 0 91816 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_993
timestamp 1586364061
transform 1 0 92460 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_989
timestamp 1586364061
transform 1 0 92092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1005
timestamp 1586364061
transform 1 0 93564 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1001
timestamp 1586364061
transform 1 0 93196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1013
timestamp 1586364061
transform 1 0 94300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 95220 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1017
timestamp 1586364061
transform 1 0 94668 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1024
timestamp 1586364061
transform 1 0 95312 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1025
timestamp 1586364061
transform 1 0 95404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 96508 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1036
timestamp 1586364061
transform 1 0 96416 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1048
timestamp 1586364061
transform 1 0 97520 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1038
timestamp 1586364061
transform 1 0 96600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1050
timestamp 1586364061
transform 1 0 97704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 98072 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1055
timestamp 1586364061
transform 1 0 98164 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1067
timestamp 1586364061
transform 1 0 99268 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1062
timestamp 1586364061
transform 1 0 98808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 100924 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1079
timestamp 1586364061
transform 1 0 100372 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1086
timestamp 1586364061
transform 1 0 101016 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1074
timestamp 1586364061
transform 1 0 99912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1086
timestamp 1586364061
transform 1 0 101016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 102120 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1098
timestamp 1586364061
transform 1 0 102120 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1099
timestamp 1586364061
transform 1 0 102212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 103776 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1110
timestamp 1586364061
transform 1 0 103224 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1117
timestamp 1586364061
transform 1 0 103868 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1111
timestamp 1586364061
transform 1 0 103316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1123
timestamp 1586364061
transform 1 0 104420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1129
timestamp 1586364061
transform 1 0 104972 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_1141
timestamp 1586364061
transform 1 0 106076 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_1135
timestamp 1586364061
transform 1 0 105524 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 106812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 106812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_1145 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 106444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_1143
timestamp 1586364061
transform 1 0 106260 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_410
timestamp 1586364061
transform 1 0 38824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_422
timestamp 1586364061
transform 1 0 39928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_434
timestamp 1586364061
transform 1 0 41032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_446
timestamp 1586364061
transform 1 0 42136 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_520
timestamp 1586364061
transform 1 0 48944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_532
timestamp 1586364061
transform 1 0 50048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_544
timestamp 1586364061
transform 1 0 51152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_556
timestamp 1586364061
transform 1 0 52256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_568
timestamp 1586364061
transform 1 0 53360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_581
timestamp 1586364061
transform 1 0 54556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_593
timestamp 1586364061
transform 1 0 55660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_605
timestamp 1586364061
transform 1 0 56764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_617
timestamp 1586364061
transform 1 0 57868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_629
timestamp 1586364061
transform 1 0 58972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_642
timestamp 1586364061
transform 1 0 60168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_654
timestamp 1586364061
transform 1 0 61272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_666
timestamp 1586364061
transform 1 0 62376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_678
timestamp 1586364061
transform 1 0 63480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_690
timestamp 1586364061
transform 1 0 64584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 65688 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_703
timestamp 1586364061
transform 1 0 65780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_715
timestamp 1586364061
transform 1 0 66884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_727
timestamp 1586364061
transform 1 0 67988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_739
timestamp 1586364061
transform 1 0 69092 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 71300 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_751
timestamp 1586364061
transform 1 0 70196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_764
timestamp 1586364061
transform 1 0 71392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_776
timestamp 1586364061
transform 1 0 72496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_788
timestamp 1586364061
transform 1 0 73600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_800
timestamp 1586364061
transform 1 0 74704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_812
timestamp 1586364061
transform 1 0 75808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 76912 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_825
timestamp 1586364061
transform 1 0 77004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_837
timestamp 1586364061
transform 1 0 78108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_849
timestamp 1586364061
transform 1 0 79212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_861
timestamp 1586364061
transform 1 0 80316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_873
timestamp 1586364061
transform 1 0 81420 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 82524 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_886
timestamp 1586364061
transform 1 0 82616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_898
timestamp 1586364061
transform 1 0 83720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_910
timestamp 1586364061
transform 1 0 84824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_922
timestamp 1586364061
transform 1 0 85928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_934
timestamp 1586364061
transform 1 0 87032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 88136 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_947
timestamp 1586364061
transform 1 0 88228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_959
timestamp 1586364061
transform 1 0 89332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_971
timestamp 1586364061
transform 1 0 90436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_983
timestamp 1586364061
transform 1 0 91540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_995
timestamp 1586364061
transform 1 0 92644 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 93748 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1008
timestamp 1586364061
transform 1 0 93840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1020
timestamp 1586364061
transform 1 0 94944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1032
timestamp 1586364061
transform 1 0 96048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1044
timestamp 1586364061
transform 1 0 97152 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 99360 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1056
timestamp 1586364061
transform 1 0 98256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1069
timestamp 1586364061
transform 1 0 99452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1081
timestamp 1586364061
transform 1 0 100556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1093
timestamp 1586364061
transform 1 0 101660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1105
timestamp 1586364061
transform 1 0 102764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1117
timestamp 1586364061
transform 1 0 103868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 104972 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1130
timestamp 1586364061
transform 1 0 105064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 106812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_1142
timestamp 1586364061
transform 1 0 106168 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_415
timestamp 1586364061
transform 1 0 39284 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_440
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_525
timestamp 1586364061
transform 1 0 49404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_537
timestamp 1586364061
transform 1 0 50508 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_550
timestamp 1586364061
transform 1 0 51704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_562
timestamp 1586364061
transform 1 0 52808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_574
timestamp 1586364061
transform 1 0 53912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_586
timestamp 1586364061
transform 1 0 55016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_598
timestamp 1586364061
transform 1 0 56120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_611
timestamp 1586364061
transform 1 0 57316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_623
timestamp 1586364061
transform 1 0 58420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_635
timestamp 1586364061
transform 1 0 59524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_647
timestamp 1586364061
transform 1 0 60628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_659
timestamp 1586364061
transform 1 0 61732 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 62836 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_672
timestamp 1586364061
transform 1 0 62928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_684
timestamp 1586364061
transform 1 0 64032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_696
timestamp 1586364061
transform 1 0 65136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_708
timestamp 1586364061
transform 1 0 66240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_720
timestamp 1586364061
transform 1 0 67344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 68448 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_733
timestamp 1586364061
transform 1 0 68540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_745
timestamp 1586364061
transform 1 0 69644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_757
timestamp 1586364061
transform 1 0 70748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_769
timestamp 1586364061
transform 1 0 71852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_781
timestamp 1586364061
transform 1 0 72956 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 74060 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_794
timestamp 1586364061
transform 1 0 74152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_806
timestamp 1586364061
transform 1 0 75256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_818
timestamp 1586364061
transform 1 0 76360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_830
timestamp 1586364061
transform 1 0 77464 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 79672 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_842
timestamp 1586364061
transform 1 0 78568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_855
timestamp 1586364061
transform 1 0 79764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_867
timestamp 1586364061
transform 1 0 80868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_879
timestamp 1586364061
transform 1 0 81972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_891
timestamp 1586364061
transform 1 0 83076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_903
timestamp 1586364061
transform 1 0 84180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 85284 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_916
timestamp 1586364061
transform 1 0 85376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_928
timestamp 1586364061
transform 1 0 86480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_940
timestamp 1586364061
transform 1 0 87584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_952
timestamp 1586364061
transform 1 0 88688 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 90896 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_964
timestamp 1586364061
transform 1 0 89792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_977
timestamp 1586364061
transform 1 0 90988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_989
timestamp 1586364061
transform 1 0 92092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1001
timestamp 1586364061
transform 1 0 93196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1013
timestamp 1586364061
transform 1 0 94300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1025
timestamp 1586364061
transform 1 0 95404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 96508 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1038
timestamp 1586364061
transform 1 0 96600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1050
timestamp 1586364061
transform 1 0 97704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1062
timestamp 1586364061
transform 1 0 98808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1074
timestamp 1586364061
transform 1 0 99912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1086
timestamp 1586364061
transform 1 0 101016 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 102120 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1099
timestamp 1586364061
transform 1 0 102212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1111
timestamp 1586364061
transform 1 0 103316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1123
timestamp 1586364061
transform 1 0 104420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_1135
timestamp 1586364061
transform 1 0 105524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 106812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_1143
timestamp 1586364061
transform 1 0 106260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_410
timestamp 1586364061
transform 1 0 38824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_422
timestamp 1586364061
transform 1 0 39928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_434
timestamp 1586364061
transform 1 0 41032 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_446
timestamp 1586364061
transform 1 0 42136 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_520
timestamp 1586364061
transform 1 0 48944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_532
timestamp 1586364061
transform 1 0 50048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_544
timestamp 1586364061
transform 1 0 51152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_556
timestamp 1586364061
transform 1 0 52256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_568
timestamp 1586364061
transform 1 0 53360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_581
timestamp 1586364061
transform 1 0 54556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_593
timestamp 1586364061
transform 1 0 55660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_605
timestamp 1586364061
transform 1 0 56764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_617
timestamp 1586364061
transform 1 0 57868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_629
timestamp 1586364061
transform 1 0 58972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_642
timestamp 1586364061
transform 1 0 60168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_654
timestamp 1586364061
transform 1 0 61272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_666
timestamp 1586364061
transform 1 0 62376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_678
timestamp 1586364061
transform 1 0 63480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_690
timestamp 1586364061
transform 1 0 64584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 65688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_703
timestamp 1586364061
transform 1 0 65780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_715
timestamp 1586364061
transform 1 0 66884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_727
timestamp 1586364061
transform 1 0 67988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_739
timestamp 1586364061
transform 1 0 69092 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 71300 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_751
timestamp 1586364061
transform 1 0 70196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_764
timestamp 1586364061
transform 1 0 71392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_776
timestamp 1586364061
transform 1 0 72496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_788
timestamp 1586364061
transform 1 0 73600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_800
timestamp 1586364061
transform 1 0 74704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_812
timestamp 1586364061
transform 1 0 75808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 76912 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_825
timestamp 1586364061
transform 1 0 77004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_837
timestamp 1586364061
transform 1 0 78108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_849
timestamp 1586364061
transform 1 0 79212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_861
timestamp 1586364061
transform 1 0 80316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_873
timestamp 1586364061
transform 1 0 81420 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 82524 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_886
timestamp 1586364061
transform 1 0 82616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_898
timestamp 1586364061
transform 1 0 83720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_910
timestamp 1586364061
transform 1 0 84824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_922
timestamp 1586364061
transform 1 0 85928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_934
timestamp 1586364061
transform 1 0 87032 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 88136 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_947
timestamp 1586364061
transform 1 0 88228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_959
timestamp 1586364061
transform 1 0 89332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_971
timestamp 1586364061
transform 1 0 90436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_983
timestamp 1586364061
transform 1 0 91540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_995
timestamp 1586364061
transform 1 0 92644 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 93748 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1008
timestamp 1586364061
transform 1 0 93840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1020
timestamp 1586364061
transform 1 0 94944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1032
timestamp 1586364061
transform 1 0 96048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1044
timestamp 1586364061
transform 1 0 97152 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 99360 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1056
timestamp 1586364061
transform 1 0 98256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1069
timestamp 1586364061
transform 1 0 99452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1081
timestamp 1586364061
transform 1 0 100556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1093
timestamp 1586364061
transform 1 0 101660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1105
timestamp 1586364061
transform 1 0 102764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1117
timestamp 1586364061
transform 1 0 103868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 104972 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1130
timestamp 1586364061
transform 1 0 105064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 106812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_1142
timestamp 1586364061
transform 1 0 106168 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_415
timestamp 1586364061
transform 1 0 39284 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_440
timestamp 1586364061
transform 1 0 41584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_464
timestamp 1586364061
transform 1 0 43792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_476
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_525
timestamp 1586364061
transform 1 0 49404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_537
timestamp 1586364061
transform 1 0 50508 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_550
timestamp 1586364061
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_562
timestamp 1586364061
transform 1 0 52808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_574
timestamp 1586364061
transform 1 0 53912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_586
timestamp 1586364061
transform 1 0 55016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_598
timestamp 1586364061
transform 1 0 56120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_611
timestamp 1586364061
transform 1 0 57316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_623
timestamp 1586364061
transform 1 0 58420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_635
timestamp 1586364061
transform 1 0 59524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_647
timestamp 1586364061
transform 1 0 60628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_659
timestamp 1586364061
transform 1 0 61732 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 62836 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_672
timestamp 1586364061
transform 1 0 62928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_684
timestamp 1586364061
transform 1 0 64032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_696
timestamp 1586364061
transform 1 0 65136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_708
timestamp 1586364061
transform 1 0 66240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_720
timestamp 1586364061
transform 1 0 67344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 68448 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_733
timestamp 1586364061
transform 1 0 68540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_745
timestamp 1586364061
transform 1 0 69644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_757
timestamp 1586364061
transform 1 0 70748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_769
timestamp 1586364061
transform 1 0 71852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_781
timestamp 1586364061
transform 1 0 72956 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 74060 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_794
timestamp 1586364061
transform 1 0 74152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_806
timestamp 1586364061
transform 1 0 75256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_818
timestamp 1586364061
transform 1 0 76360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_830
timestamp 1586364061
transform 1 0 77464 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 79672 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_842
timestamp 1586364061
transform 1 0 78568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_855
timestamp 1586364061
transform 1 0 79764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_867
timestamp 1586364061
transform 1 0 80868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_879
timestamp 1586364061
transform 1 0 81972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_891
timestamp 1586364061
transform 1 0 83076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_903
timestamp 1586364061
transform 1 0 84180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 85284 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_916
timestamp 1586364061
transform 1 0 85376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_928
timestamp 1586364061
transform 1 0 86480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_940
timestamp 1586364061
transform 1 0 87584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_952
timestamp 1586364061
transform 1 0 88688 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 90896 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_964
timestamp 1586364061
transform 1 0 89792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_977
timestamp 1586364061
transform 1 0 90988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_989
timestamp 1586364061
transform 1 0 92092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1001
timestamp 1586364061
transform 1 0 93196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1013
timestamp 1586364061
transform 1 0 94300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1025
timestamp 1586364061
transform 1 0 95404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 96508 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1038
timestamp 1586364061
transform 1 0 96600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1050
timestamp 1586364061
transform 1 0 97704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1062
timestamp 1586364061
transform 1 0 98808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1074
timestamp 1586364061
transform 1 0 99912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1086
timestamp 1586364061
transform 1 0 101016 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 102120 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1099
timestamp 1586364061
transform 1 0 102212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1111
timestamp 1586364061
transform 1 0 103316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1123
timestamp 1586364061
transform 1 0 104420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_1135
timestamp 1586364061
transform 1 0 105524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 106812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_1143
timestamp 1586364061
transform 1 0 106260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__11__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_189
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_410
timestamp 1586364061
transform 1 0 38824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_422
timestamp 1586364061
transform 1 0 39928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_415
timestamp 1586364061
transform 1 0 39284 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_434
timestamp 1586364061
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_446
timestamp 1586364061
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_452
timestamp 1586364061
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_471
timestamp 1586364061
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_464
timestamp 1586364061
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_476
timestamp 1586364061
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_483
timestamp 1586364061
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_495
timestamp 1586364061
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_507
timestamp 1586364061
transform 1 0 47748 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_501
timestamp 1586364061
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_520
timestamp 1586364061
transform 1 0 48944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_532
timestamp 1586364061
transform 1 0 50048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_525
timestamp 1586364061
transform 1 0 49404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_544
timestamp 1586364061
transform 1 0 51152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_537
timestamp 1586364061
transform 1 0 50508 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_550
timestamp 1586364061
transform 1 0 51704 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_556
timestamp 1586364061
transform 1 0 52256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_568
timestamp 1586364061
transform 1 0 53360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_562
timestamp 1586364061
transform 1 0 52808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_581
timestamp 1586364061
transform 1 0 54556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_574
timestamp 1586364061
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_586
timestamp 1586364061
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_593
timestamp 1586364061
transform 1 0 55660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_605
timestamp 1586364061
transform 1 0 56764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_598
timestamp 1586364061
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_617
timestamp 1586364061
transform 1 0 57868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_611
timestamp 1586364061
transform 1 0 57316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_623
timestamp 1586364061
transform 1 0 58420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_629
timestamp 1586364061
transform 1 0 58972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_642
timestamp 1586364061
transform 1 0 60168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_635
timestamp 1586364061
transform 1 0 59524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_654
timestamp 1586364061
transform 1 0 61272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_647
timestamp 1586364061
transform 1 0 60628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_659
timestamp 1586364061
transform 1 0 61732 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_666
timestamp 1586364061
transform 1 0 62376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_672
timestamp 1586364061
transform 1 0 62928 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_678
timestamp 1586364061
transform 1 0 63480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_690
timestamp 1586364061
transform 1 0 64584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_684
timestamp 1586364061
transform 1 0 64032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 65688 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_703
timestamp 1586364061
transform 1 0 65780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_696
timestamp 1586364061
transform 1 0 65136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_708
timestamp 1586364061
transform 1 0 66240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_715
timestamp 1586364061
transform 1 0 66884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_727
timestamp 1586364061
transform 1 0 67988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_720
timestamp 1586364061
transform 1 0 67344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 68448 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_739
timestamp 1586364061
transform 1 0 69092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_733
timestamp 1586364061
transform 1 0 68540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_745
timestamp 1586364061
transform 1 0 69644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 71300 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_751
timestamp 1586364061
transform 1 0 70196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_764
timestamp 1586364061
transform 1 0 71392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_757
timestamp 1586364061
transform 1 0 70748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_776
timestamp 1586364061
transform 1 0 72496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_769
timestamp 1586364061
transform 1 0 71852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_781
timestamp 1586364061
transform 1 0 72956 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 74060 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_788
timestamp 1586364061
transform 1 0 73600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_800
timestamp 1586364061
transform 1 0 74704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_794
timestamp 1586364061
transform 1 0 74152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_812
timestamp 1586364061
transform 1 0 75808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_806
timestamp 1586364061
transform 1 0 75256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_818
timestamp 1586364061
transform 1 0 76360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_825
timestamp 1586364061
transform 1 0 77004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_837
timestamp 1586364061
transform 1 0 78108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_830
timestamp 1586364061
transform 1 0 77464 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 79672 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_849
timestamp 1586364061
transform 1 0 79212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_842
timestamp 1586364061
transform 1 0 78568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_855
timestamp 1586364061
transform 1 0 79764 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_861
timestamp 1586364061
transform 1 0 80316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_873
timestamp 1586364061
transform 1 0 81420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_867
timestamp 1586364061
transform 1 0 80868 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 82524 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_886
timestamp 1586364061
transform 1 0 82616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_879
timestamp 1586364061
transform 1 0 81972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_891
timestamp 1586364061
transform 1 0 83076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_898
timestamp 1586364061
transform 1 0 83720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_903
timestamp 1586364061
transform 1 0 84180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 85284 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_910
timestamp 1586364061
transform 1 0 84824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_922
timestamp 1586364061
transform 1 0 85928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_916
timestamp 1586364061
transform 1 0 85376 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_934
timestamp 1586364061
transform 1 0 87032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_928
timestamp 1586364061
transform 1 0 86480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_940
timestamp 1586364061
transform 1 0 87584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 88136 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_947
timestamp 1586364061
transform 1 0 88228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_959
timestamp 1586364061
transform 1 0 89332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_952
timestamp 1586364061
transform 1 0 88688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 90896 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_971
timestamp 1586364061
transform 1 0 90436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_964
timestamp 1586364061
transform 1 0 89792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_977
timestamp 1586364061
transform 1 0 90988 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_983
timestamp 1586364061
transform 1 0 91540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_995
timestamp 1586364061
transform 1 0 92644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_989
timestamp 1586364061
transform 1 0 92092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 93748 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1008
timestamp 1586364061
transform 1 0 93840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1001
timestamp 1586364061
transform 1 0 93196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1013
timestamp 1586364061
transform 1 0 94300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1020
timestamp 1586364061
transform 1 0 94944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1032
timestamp 1586364061
transform 1 0 96048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1025
timestamp 1586364061
transform 1 0 95404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 96508 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1044
timestamp 1586364061
transform 1 0 97152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1038
timestamp 1586364061
transform 1 0 96600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1050
timestamp 1586364061
transform 1 0 97704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 99360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1056
timestamp 1586364061
transform 1 0 98256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1069
timestamp 1586364061
transform 1 0 99452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1062
timestamp 1586364061
transform 1 0 98808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1081
timestamp 1586364061
transform 1 0 100556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1074
timestamp 1586364061
transform 1 0 99912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1086
timestamp 1586364061
transform 1 0 101016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 102120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1093
timestamp 1586364061
transform 1 0 101660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1105
timestamp 1586364061
transform 1 0 102764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1099
timestamp 1586364061
transform 1 0 102212 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1117
timestamp 1586364061
transform 1 0 103868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1111
timestamp 1586364061
transform 1 0 103316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1123
timestamp 1586364061
transform 1 0 104420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 104972 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1130
timestamp 1586364061
transform 1 0 105064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_1135
timestamp 1586364061
transform 1 0 105524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 106812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 106812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_1142
timestamp 1586364061
transform 1 0 106168 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_1143
timestamp 1586364061
transform 1 0 106260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _11_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _08_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_255
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_410
timestamp 1586364061
transform 1 0 38824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_422
timestamp 1586364061
transform 1 0 39928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_434
timestamp 1586364061
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_446
timestamp 1586364061
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_459
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_471
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_483
timestamp 1586364061
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_495
timestamp 1586364061
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_507
timestamp 1586364061
transform 1 0 47748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_520
timestamp 1586364061
transform 1 0 48944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_532
timestamp 1586364061
transform 1 0 50048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_544
timestamp 1586364061
transform 1 0 51152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_556
timestamp 1586364061
transform 1 0 52256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_568
timestamp 1586364061
transform 1 0 53360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_581
timestamp 1586364061
transform 1 0 54556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_593
timestamp 1586364061
transform 1 0 55660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_605
timestamp 1586364061
transform 1 0 56764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_617
timestamp 1586364061
transform 1 0 57868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_629
timestamp 1586364061
transform 1 0 58972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_642
timestamp 1586364061
transform 1 0 60168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_654
timestamp 1586364061
transform 1 0 61272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_666
timestamp 1586364061
transform 1 0 62376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_678
timestamp 1586364061
transform 1 0 63480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_690
timestamp 1586364061
transform 1 0 64584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 65688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_703
timestamp 1586364061
transform 1 0 65780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_715
timestamp 1586364061
transform 1 0 66884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_727
timestamp 1586364061
transform 1 0 67988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_739
timestamp 1586364061
transform 1 0 69092 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 71300 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_751
timestamp 1586364061
transform 1 0 70196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_764
timestamp 1586364061
transform 1 0 71392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_776
timestamp 1586364061
transform 1 0 72496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_788
timestamp 1586364061
transform 1 0 73600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_800
timestamp 1586364061
transform 1 0 74704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_812
timestamp 1586364061
transform 1 0 75808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_825
timestamp 1586364061
transform 1 0 77004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_837
timestamp 1586364061
transform 1 0 78108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_849
timestamp 1586364061
transform 1 0 79212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_861
timestamp 1586364061
transform 1 0 80316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_873
timestamp 1586364061
transform 1 0 81420 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 82524 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_886
timestamp 1586364061
transform 1 0 82616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_898
timestamp 1586364061
transform 1 0 83720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_910
timestamp 1586364061
transform 1 0 84824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_922
timestamp 1586364061
transform 1 0 85928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_934
timestamp 1586364061
transform 1 0 87032 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 88136 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_947
timestamp 1586364061
transform 1 0 88228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_959
timestamp 1586364061
transform 1 0 89332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_971
timestamp 1586364061
transform 1 0 90436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_983
timestamp 1586364061
transform 1 0 91540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_995
timestamp 1586364061
transform 1 0 92644 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 93748 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1008
timestamp 1586364061
transform 1 0 93840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1020
timestamp 1586364061
transform 1 0 94944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1032
timestamp 1586364061
transform 1 0 96048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1044
timestamp 1586364061
transform 1 0 97152 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 99360 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1056
timestamp 1586364061
transform 1 0 98256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1069
timestamp 1586364061
transform 1 0 99452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1081
timestamp 1586364061
transform 1 0 100556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1093
timestamp 1586364061
transform 1 0 101660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1105
timestamp 1586364061
transform 1 0 102764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1117
timestamp 1586364061
transform 1 0 103868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 104972 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1130
timestamp 1586364061
transform 1 0 105064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 106812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_1142
timestamp 1586364061
transform 1 0 106168 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_and4_4  _07_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_415
timestamp 1586364061
transform 1 0 39284 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_440
timestamp 1586364061
transform 1 0 41584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_452
timestamp 1586364061
transform 1 0 42688 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_464
timestamp 1586364061
transform 1 0 43792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_476
timestamp 1586364061
transform 1 0 44896 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_489
timestamp 1586364061
transform 1 0 46092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_501
timestamp 1586364061
transform 1 0 47196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_513
timestamp 1586364061
transform 1 0 48300 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_525
timestamp 1586364061
transform 1 0 49404 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 51612 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_537
timestamp 1586364061
transform 1 0 50508 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_550
timestamp 1586364061
transform 1 0 51704 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_562
timestamp 1586364061
transform 1 0 52808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_574
timestamp 1586364061
transform 1 0 53912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_586
timestamp 1586364061
transform 1 0 55016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_598
timestamp 1586364061
transform 1 0 56120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 57224 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_611
timestamp 1586364061
transform 1 0 57316 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_623
timestamp 1586364061
transform 1 0 58420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_635
timestamp 1586364061
transform 1 0 59524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_647
timestamp 1586364061
transform 1 0 60628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_659
timestamp 1586364061
transform 1 0 61732 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 62836 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_672
timestamp 1586364061
transform 1 0 62928 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_684
timestamp 1586364061
transform 1 0 64032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_696
timestamp 1586364061
transform 1 0 65136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_708
timestamp 1586364061
transform 1 0 66240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_720
timestamp 1586364061
transform 1 0 67344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 68448 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_733
timestamp 1586364061
transform 1 0 68540 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_745
timestamp 1586364061
transform 1 0 69644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_757
timestamp 1586364061
transform 1 0 70748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_769
timestamp 1586364061
transform 1 0 71852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_781
timestamp 1586364061
transform 1 0 72956 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 74060 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_794
timestamp 1586364061
transform 1 0 74152 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_806
timestamp 1586364061
transform 1 0 75256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_818
timestamp 1586364061
transform 1 0 76360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_830
timestamp 1586364061
transform 1 0 77464 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 79672 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_842
timestamp 1586364061
transform 1 0 78568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_855
timestamp 1586364061
transform 1 0 79764 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_867
timestamp 1586364061
transform 1 0 80868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_879
timestamp 1586364061
transform 1 0 81972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_891
timestamp 1586364061
transform 1 0 83076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_903
timestamp 1586364061
transform 1 0 84180 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 85284 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_916
timestamp 1586364061
transform 1 0 85376 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_928
timestamp 1586364061
transform 1 0 86480 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_940
timestamp 1586364061
transform 1 0 87584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_952
timestamp 1586364061
transform 1 0 88688 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 90896 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_964
timestamp 1586364061
transform 1 0 89792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_977
timestamp 1586364061
transform 1 0 90988 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_989
timestamp 1586364061
transform 1 0 92092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1001
timestamp 1586364061
transform 1 0 93196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1013
timestamp 1586364061
transform 1 0 94300 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1025
timestamp 1586364061
transform 1 0 95404 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 96508 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1038
timestamp 1586364061
transform 1 0 96600 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1050
timestamp 1586364061
transform 1 0 97704 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1062
timestamp 1586364061
transform 1 0 98808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1074
timestamp 1586364061
transform 1 0 99912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1086
timestamp 1586364061
transform 1 0 101016 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 102120 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1099
timestamp 1586364061
transform 1 0 102212 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1111
timestamp 1586364061
transform 1 0 103316 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1123
timestamp 1586364061
transform 1 0 104420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_1135
timestamp 1586364061
transform 1 0 105524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 106812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_1143
timestamp 1586364061
transform 1 0 106260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 774 592
use scs8hd_nor4_4  _13_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 1602 592
use scs8hd_fill_1  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_and4_4  _05_
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_229
timestamp 1586364061
transform 1 0 22172 0 -1 8160
box -38 -48 774 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 22908 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_373
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36340 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_381
timestamp 1586364061
transform 1 0 36156 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_385
timestamp 1586364061
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_410
timestamp 1586364061
transform 1 0 38824 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_422
timestamp 1586364061
transform 1 0 39928 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_434
timestamp 1586364061
transform 1 0 41032 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_446
timestamp 1586364061
transform 1 0 42136 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_459
timestamp 1586364061
transform 1 0 43332 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_471
timestamp 1586364061
transform 1 0 44436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_483
timestamp 1586364061
transform 1 0 45540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_495
timestamp 1586364061
transform 1 0 46644 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_507
timestamp 1586364061
transform 1 0 47748 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 48852 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_520
timestamp 1586364061
transform 1 0 48944 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_532
timestamp 1586364061
transform 1 0 50048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_544
timestamp 1586364061
transform 1 0 51152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_556
timestamp 1586364061
transform 1 0 52256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_568
timestamp 1586364061
transform 1 0 53360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 54464 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_581
timestamp 1586364061
transform 1 0 54556 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_593
timestamp 1586364061
transform 1 0 55660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_605
timestamp 1586364061
transform 1 0 56764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_617
timestamp 1586364061
transform 1 0 57868 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 60076 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_629
timestamp 1586364061
transform 1 0 58972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_642
timestamp 1586364061
transform 1 0 60168 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_654
timestamp 1586364061
transform 1 0 61272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_666
timestamp 1586364061
transform 1 0 62376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_678
timestamp 1586364061
transform 1 0 63480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_690
timestamp 1586364061
transform 1 0 64584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 65688 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_703
timestamp 1586364061
transform 1 0 65780 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_715
timestamp 1586364061
transform 1 0 66884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_727
timestamp 1586364061
transform 1 0 67988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_739
timestamp 1586364061
transform 1 0 69092 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 71300 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_751
timestamp 1586364061
transform 1 0 70196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_764
timestamp 1586364061
transform 1 0 71392 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_776
timestamp 1586364061
transform 1 0 72496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_788
timestamp 1586364061
transform 1 0 73600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_800
timestamp 1586364061
transform 1 0 74704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_812
timestamp 1586364061
transform 1 0 75808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 76912 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_825
timestamp 1586364061
transform 1 0 77004 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_837
timestamp 1586364061
transform 1 0 78108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_849
timestamp 1586364061
transform 1 0 79212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_861
timestamp 1586364061
transform 1 0 80316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_873
timestamp 1586364061
transform 1 0 81420 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 82524 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_886
timestamp 1586364061
transform 1 0 82616 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_898
timestamp 1586364061
transform 1 0 83720 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_910
timestamp 1586364061
transform 1 0 84824 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_922
timestamp 1586364061
transform 1 0 85928 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_934
timestamp 1586364061
transform 1 0 87032 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 88136 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_947
timestamp 1586364061
transform 1 0 88228 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_959
timestamp 1586364061
transform 1 0 89332 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_971
timestamp 1586364061
transform 1 0 90436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_983
timestamp 1586364061
transform 1 0 91540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_995
timestamp 1586364061
transform 1 0 92644 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 93748 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_1008
timestamp 1586364061
transform 1 0 93840 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1020
timestamp 1586364061
transform 1 0 94944 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1032
timestamp 1586364061
transform 1 0 96048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1044
timestamp 1586364061
transform 1 0 97152 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 99360 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_1056
timestamp 1586364061
transform 1 0 98256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1069
timestamp 1586364061
transform 1 0 99452 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1081
timestamp 1586364061
transform 1 0 100556 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1093
timestamp 1586364061
transform 1 0 101660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1105
timestamp 1586364061
transform 1 0 102764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_1117
timestamp 1586364061
transform 1 0 103868 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 104972 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_1130
timestamp 1586364061
transform 1 0 105064 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 106812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_1142
timestamp 1586364061
transform 1 0 106168 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _15_
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 590 592
use scs8hd_decap_4  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _14_
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 130 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_336
timestamp 1586364061
transform 1 0 32016 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_339
timestamp 1586364061
transform 1 0 32292 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_343
timestamp 1586364061
transform 1 0 32660 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_355
timestamp 1586364061
transform 1 0 33764 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35420 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_363
timestamp 1586364061
transform 1 0 34500 0 1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36340 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 36156 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35788 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_375
timestamp 1586364061
transform 1 0 35604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_379
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_394
timestamp 1586364061
transform 1 0 37352 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_400
timestamp 1586364061
transform 1 0 37904 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_404
timestamp 1586364061
transform 1 0 38272 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_416
timestamp 1586364061
transform 1 0 39376 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_424
timestamp 1586364061
transform 1 0 40112 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_428
timestamp 1586364061
transform 1 0 40480 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_440
timestamp 1586364061
transform 1 0 41584 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_452
timestamp 1586364061
transform 1 0 42688 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_464
timestamp 1586364061
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_476
timestamp 1586364061
transform 1 0 44896 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_489
timestamp 1586364061
transform 1 0 46092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_501
timestamp 1586364061
transform 1 0 47196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_513
timestamp 1586364061
transform 1 0 48300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_525
timestamp 1586364061
transform 1 0 49404 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 51612 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_537
timestamp 1586364061
transform 1 0 50508 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_550
timestamp 1586364061
transform 1 0 51704 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_562
timestamp 1586364061
transform 1 0 52808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_574
timestamp 1586364061
transform 1 0 53912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_586
timestamp 1586364061
transform 1 0 55016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_598
timestamp 1586364061
transform 1 0 56120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 57224 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_611
timestamp 1586364061
transform 1 0 57316 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_623
timestamp 1586364061
transform 1 0 58420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_635
timestamp 1586364061
transform 1 0 59524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_647
timestamp 1586364061
transform 1 0 60628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_659
timestamp 1586364061
transform 1 0 61732 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 62836 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_672
timestamp 1586364061
transform 1 0 62928 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_684
timestamp 1586364061
transform 1 0 64032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_696
timestamp 1586364061
transform 1 0 65136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_708
timestamp 1586364061
transform 1 0 66240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_720
timestamp 1586364061
transform 1 0 67344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 68448 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_733
timestamp 1586364061
transform 1 0 68540 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_745
timestamp 1586364061
transform 1 0 69644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_757
timestamp 1586364061
transform 1 0 70748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_769
timestamp 1586364061
transform 1 0 71852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_781
timestamp 1586364061
transform 1 0 72956 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 74060 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_794
timestamp 1586364061
transform 1 0 74152 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_806
timestamp 1586364061
transform 1 0 75256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_818
timestamp 1586364061
transform 1 0 76360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_830
timestamp 1586364061
transform 1 0 77464 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 79672 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_842
timestamp 1586364061
transform 1 0 78568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_855
timestamp 1586364061
transform 1 0 79764 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_867
timestamp 1586364061
transform 1 0 80868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_879
timestamp 1586364061
transform 1 0 81972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_891
timestamp 1586364061
transform 1 0 83076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_903
timestamp 1586364061
transform 1 0 84180 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 85284 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_916
timestamp 1586364061
transform 1 0 85376 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_928
timestamp 1586364061
transform 1 0 86480 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_940
timestamp 1586364061
transform 1 0 87584 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_952
timestamp 1586364061
transform 1 0 88688 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 90896 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_964
timestamp 1586364061
transform 1 0 89792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_977
timestamp 1586364061
transform 1 0 90988 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_989
timestamp 1586364061
transform 1 0 92092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1001
timestamp 1586364061
transform 1 0 93196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1013
timestamp 1586364061
transform 1 0 94300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1025
timestamp 1586364061
transform 1 0 95404 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 96508 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_1038
timestamp 1586364061
transform 1 0 96600 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1050
timestamp 1586364061
transform 1 0 97704 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1062
timestamp 1586364061
transform 1 0 98808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1074
timestamp 1586364061
transform 1 0 99912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1086
timestamp 1586364061
transform 1 0 101016 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 102120 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_1099
timestamp 1586364061
transform 1 0 102212 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1111
timestamp 1586364061
transform 1 0 103316 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_1123
timestamp 1586364061
transform 1 0 104420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_1135
timestamp 1586364061
transform 1 0 105524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 106812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_1143
timestamp 1586364061
transform 1 0 106260 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_14
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_26
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_and4_4  _09_
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_244
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_256
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_268
timestamp 1586364061
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_348
timestamp 1586364061
transform 1 0 33120 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_360
timestamp 1586364061
transform 1 0 34224 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_372
timestamp 1586364061
transform 1 0 35328 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 35880 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_389
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_409
timestamp 1586364061
transform 1 0 38732 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_421
timestamp 1586364061
transform 1 0 39836 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_433
timestamp 1586364061
transform 1 0 40940 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_445
timestamp 1586364061
transform 1 0 42044 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_457
timestamp 1586364061
transform 1 0 43148 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_459
timestamp 1586364061
transform 1 0 43332 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_471
timestamp 1586364061
transform 1 0 44436 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_483
timestamp 1586364061
transform 1 0 45540 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_495
timestamp 1586364061
transform 1 0 46644 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_507
timestamp 1586364061
transform 1 0 47748 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 48852 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_520
timestamp 1586364061
transform 1 0 48944 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_532
timestamp 1586364061
transform 1 0 50048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_544
timestamp 1586364061
transform 1 0 51152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_556
timestamp 1586364061
transform 1 0 52256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_568
timestamp 1586364061
transform 1 0 53360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 54464 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_581
timestamp 1586364061
transform 1 0 54556 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_593
timestamp 1586364061
transform 1 0 55660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_605
timestamp 1586364061
transform 1 0 56764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_617
timestamp 1586364061
transform 1 0 57868 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 60076 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_629
timestamp 1586364061
transform 1 0 58972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_642
timestamp 1586364061
transform 1 0 60168 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_654
timestamp 1586364061
transform 1 0 61272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_666
timestamp 1586364061
transform 1 0 62376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_678
timestamp 1586364061
transform 1 0 63480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_690
timestamp 1586364061
transform 1 0 64584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 65688 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_703
timestamp 1586364061
transform 1 0 65780 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_715
timestamp 1586364061
transform 1 0 66884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_727
timestamp 1586364061
transform 1 0 67988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_739
timestamp 1586364061
transform 1 0 69092 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 71300 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_751
timestamp 1586364061
transform 1 0 70196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_764
timestamp 1586364061
transform 1 0 71392 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_776
timestamp 1586364061
transform 1 0 72496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_788
timestamp 1586364061
transform 1 0 73600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_800
timestamp 1586364061
transform 1 0 74704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_812
timestamp 1586364061
transform 1 0 75808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 76912 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_825
timestamp 1586364061
transform 1 0 77004 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_837
timestamp 1586364061
transform 1 0 78108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_849
timestamp 1586364061
transform 1 0 79212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_861
timestamp 1586364061
transform 1 0 80316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_873
timestamp 1586364061
transform 1 0 81420 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 82524 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_886
timestamp 1586364061
transform 1 0 82616 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_898
timestamp 1586364061
transform 1 0 83720 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_910
timestamp 1586364061
transform 1 0 84824 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_922
timestamp 1586364061
transform 1 0 85928 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_934
timestamp 1586364061
transform 1 0 87032 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 88136 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_947
timestamp 1586364061
transform 1 0 88228 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_959
timestamp 1586364061
transform 1 0 89332 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_971
timestamp 1586364061
transform 1 0 90436 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_983
timestamp 1586364061
transform 1 0 91540 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_995
timestamp 1586364061
transform 1 0 92644 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 93748 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_1008
timestamp 1586364061
transform 1 0 93840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1020
timestamp 1586364061
transform 1 0 94944 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1032
timestamp 1586364061
transform 1 0 96048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1044
timestamp 1586364061
transform 1 0 97152 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 99360 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_1056
timestamp 1586364061
transform 1 0 98256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1069
timestamp 1586364061
transform 1 0 99452 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1081
timestamp 1586364061
transform 1 0 100556 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1093
timestamp 1586364061
transform 1 0 101660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1105
timestamp 1586364061
transform 1 0 102764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_1117
timestamp 1586364061
transform 1 0 103868 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 104972 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_1130
timestamp 1586364061
transform 1 0 105064 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 106812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_1142
timestamp 1586364061
transform 1 0 106168 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _19_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_128
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 21804 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_222
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_223
timestamp 1586364061
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_233
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_245
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_257
timestamp 1586364061
transform 1 0 24748 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_278
timestamp 1586364061
transform 1 0 26680 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_269
timestamp 1586364061
transform 1 0 25852 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_280
timestamp 1586364061
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_290
timestamp 1586364061
transform 1 0 27784 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_13_302
timestamp 1586364061
transform 1 0 28888 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_292
timestamp 1586364061
transform 1 0 27968 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_304
timestamp 1586364061
transform 1 0 29072 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_316
timestamp 1586364061
transform 1 0 30176 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_328
timestamp 1586364061
transform 1 0 31280 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 34960 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 35052 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 35420 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_371
timestamp 1586364061
transform 1 0 35236 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_367
timestamp 1586364061
transform 1 0 34868 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 36156 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36156 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_375
timestamp 1586364061
transform 1 0 35604 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_392
timestamp 1586364061
transform 1 0 37168 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_376
timestamp 1586364061
transform 1 0 35696 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_380
timestamp 1586364061
transform 1 0 36064 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_383
timestamp 1586364061
transform 1 0 36340 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_404
timestamp 1586364061
transform 1 0 38272 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_395
timestamp 1586364061
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_410
timestamp 1586364061
transform 1 0 38824 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 39192 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 39192 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_412
timestamp 1586364061
transform 1 0 39008 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_416
timestamp 1586364061
transform 1 0 39376 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_424
timestamp 1586364061
transform 1 0 40112 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_428
timestamp 1586364061
transform 1 0 40480 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_418
timestamp 1586364061
transform 1 0 39560 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_440
timestamp 1586364061
transform 1 0 41584 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_430
timestamp 1586364061
transform 1 0 40664 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_442
timestamp 1586364061
transform 1 0 41768 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_452
timestamp 1586364061
transform 1 0 42688 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_454
timestamp 1586364061
transform 1 0 42872 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_459
timestamp 1586364061
transform 1 0 43332 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_464
timestamp 1586364061
transform 1 0 43792 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_476
timestamp 1586364061
transform 1 0 44896 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_471
timestamp 1586364061
transform 1 0 44436 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_489
timestamp 1586364061
transform 1 0 46092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_483
timestamp 1586364061
transform 1 0 45540 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_495
timestamp 1586364061
transform 1 0 46644 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_501
timestamp 1586364061
transform 1 0 47196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_513
timestamp 1586364061
transform 1 0 48300 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_507
timestamp 1586364061
transform 1 0 47748 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 48944 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 48852 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 48944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 49312 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_519
timestamp 1586364061
transform 1 0 48852 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_522
timestamp 1586364061
transform 1 0 49128 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_526
timestamp 1586364061
transform 1 0 49496 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_528
timestamp 1586364061
transform 1 0 49680 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 51612 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_538
timestamp 1586364061
transform 1 0 50600 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_546
timestamp 1586364061
transform 1 0 51336 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_13_550
timestamp 1586364061
transform 1 0 51704 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_540
timestamp 1586364061
transform 1 0 50784 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_552
timestamp 1586364061
transform 1 0 51888 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 52716 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 52716 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_558
timestamp 1586364061
transform 1 0 52440 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_563
timestamp 1586364061
transform 1 0 52900 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_560
timestamp 1586364061
transform 1 0 52624 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_565
timestamp 1586364061
transform 1 0 53084 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 54464 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_575
timestamp 1586364061
transform 1 0 54004 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_587
timestamp 1586364061
transform 1 0 55108 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_577
timestamp 1586364061
transform 1 0 54188 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_581
timestamp 1586364061
transform 1 0 54556 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_599
timestamp 1586364061
transform 1 0 56212 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_593
timestamp 1586364061
transform 1 0 55660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_605
timestamp 1586364061
transform 1 0 56764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 57224 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_607
timestamp 1586364061
transform 1 0 56948 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_611
timestamp 1586364061
transform 1 0 57316 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_623
timestamp 1586364061
transform 1 0 58420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_617
timestamp 1586364061
transform 1 0 57868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 60076 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_635
timestamp 1586364061
transform 1 0 59524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_629
timestamp 1586364061
transform 1 0 58972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_642
timestamp 1586364061
transform 1 0 60168 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 61456 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 61456 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_647
timestamp 1586364061
transform 1 0 60628 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_655
timestamp 1586364061
transform 1 0 61364 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_658
timestamp 1586364061
transform 1 0 61640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_654
timestamp 1586364061
transform 1 0 61272 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 62836 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 61824 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_662
timestamp 1586364061
transform 1 0 62008 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_670
timestamp 1586364061
transform 1 0 62744 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_672
timestamp 1586364061
transform 1 0 62928 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_664
timestamp 1586364061
transform 1 0 62192 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_676
timestamp 1586364061
transform 1 0 63296 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_684
timestamp 1586364061
transform 1 0 64032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_688
timestamp 1586364061
transform 1 0 64400 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 66148 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 65688 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 66148 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_696
timestamp 1586364061
transform 1 0 65136 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_704
timestamp 1586364061
transform 1 0 65872 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_709
timestamp 1586364061
transform 1 0 66332 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_700
timestamp 1586364061
transform 1 0 65504 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_703
timestamp 1586364061
transform 1 0 65780 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_711
timestamp 1586364061
transform 1 0 66516 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_721
timestamp 1586364061
transform 1 0 67436 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_729
timestamp 1586364061
transform 1 0 68172 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_723
timestamp 1586364061
transform 1 0 67620 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 68448 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_733
timestamp 1586364061
transform 1 0 68540 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_745
timestamp 1586364061
transform 1 0 69644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_735
timestamp 1586364061
transform 1 0 68724 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_747
timestamp 1586364061
transform 1 0 69828 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 71300 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_757
timestamp 1586364061
transform 1 0 70748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_759
timestamp 1586364061
transform 1 0 70932 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_764
timestamp 1586364061
transform 1 0 71392 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_769
timestamp 1586364061
transform 1 0 71852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_781
timestamp 1586364061
transform 1 0 72956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_776
timestamp 1586364061
transform 1 0 72496 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 74060 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_794
timestamp 1586364061
transform 1 0 74152 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_802
timestamp 1586364061
transform 1 0 74888 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_788
timestamp 1586364061
transform 1 0 73600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_800
timestamp 1586364061
transform 1 0 74704 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 75072 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 75072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 75440 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_806
timestamp 1586364061
transform 1 0 75256 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_810
timestamp 1586364061
transform 1 0 75624 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_812
timestamp 1586364061
transform 1 0 75808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 76912 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_822
timestamp 1586364061
transform 1 0 76728 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_834
timestamp 1586364061
transform 1 0 77832 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_825
timestamp 1586364061
transform 1 0 77004 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_837
timestamp 1586364061
transform 1 0 78108 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 79672 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 79672 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_846
timestamp 1586364061
transform 1 0 78936 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_855
timestamp 1586364061
transform 1 0 79764 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_849
timestamp 1586364061
transform 1 0 79212 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_853
timestamp 1586364061
transform 1 0 79580 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 79948 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_859
timestamp 1586364061
transform 1 0 80132 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_871
timestamp 1586364061
transform 1 0 81236 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_858
timestamp 1586364061
transform 1 0 80040 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_870
timestamp 1586364061
transform 1 0 81144 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 82524 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_883
timestamp 1586364061
transform 1 0 82340 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_882
timestamp 1586364061
transform 1 0 82248 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_886
timestamp 1586364061
transform 1 0 82616 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_895
timestamp 1586364061
transform 1 0 83444 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_907
timestamp 1586364061
transform 1 0 84548 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_898
timestamp 1586364061
transform 1 0 83720 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 85284 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_916
timestamp 1586364061
transform 1 0 85376 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_910
timestamp 1586364061
transform 1 0 84824 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_922
timestamp 1586364061
transform 1 0 85928 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 88044 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 87860 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_928
timestamp 1586364061
transform 1 0 86480 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_13_940
timestamp 1586364061
transform 1 0 87584 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_934
timestamp 1586364061
transform 1 0 87032 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 88228 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 88136 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 88596 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 88964 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_949
timestamp 1586364061
transform 1 0 88412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_953
timestamp 1586364061
transform 1 0 88780 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_957
timestamp 1586364061
transform 1 0 89148 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_955
timestamp 1586364061
transform 1 0 88964 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 90896 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_969
timestamp 1586364061
transform 1 0 90252 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_975
timestamp 1586364061
transform 1 0 90804 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_977
timestamp 1586364061
transform 1 0 90988 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_967
timestamp 1586364061
transform 1 0 90068 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_979
timestamp 1586364061
transform 1 0 91172 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_989
timestamp 1586364061
transform 1 0 92092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_991
timestamp 1586364061
transform 1 0 92276 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 93748 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1001
timestamp 1586364061
transform 1 0 93196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1013
timestamp 1586364061
transform 1 0 94300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_1003
timestamp 1586364061
transform 1 0 93380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_1008
timestamp 1586364061
transform 1 0 93840 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1025
timestamp 1586364061
transform 1 0 95404 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1020
timestamp 1586364061
transform 1 0 94944 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1032
timestamp 1586364061
transform 1 0 96048 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 96508 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1038
timestamp 1586364061
transform 1 0 96600 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1050
timestamp 1586364061
transform 1 0 97704 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1044
timestamp 1586364061
transform 1 0 97152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 99360 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1062
timestamp 1586364061
transform 1 0 98808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1056
timestamp 1586364061
transform 1 0 98256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1069
timestamp 1586364061
transform 1 0 99452 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1074
timestamp 1586364061
transform 1 0 99912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1086
timestamp 1586364061
transform 1 0 101016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1081
timestamp 1586364061
transform 1 0 100556 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 102120 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_1099
timestamp 1586364061
transform 1 0 102212 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1093
timestamp 1586364061
transform 1 0 101660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1105
timestamp 1586364061
transform 1 0 102764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1111
timestamp 1586364061
transform 1 0 103316 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_1123
timestamp 1586364061
transform 1 0 104420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_1117
timestamp 1586364061
transform 1 0 103868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 104972 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_1135
timestamp 1586364061
transform 1 0 105524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_1130
timestamp 1586364061
transform 1 0 105064 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 106812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 106812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_1143
timestamp 1586364061
transform 1 0 106260 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_1142
timestamp 1586364061
transform 1 0 106168 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_415
timestamp 1586364061
transform 1 0 39284 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_428
timestamp 1586364061
transform 1 0 40480 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_440
timestamp 1586364061
transform 1 0 41584 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_452
timestamp 1586364061
transform 1 0 42688 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_464
timestamp 1586364061
transform 1 0 43792 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_476
timestamp 1586364061
transform 1 0 44896 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_489
timestamp 1586364061
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_501
timestamp 1586364061
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_513
timestamp 1586364061
transform 1 0 48300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_525
timestamp 1586364061
transform 1 0 49404 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 51612 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_537
timestamp 1586364061
transform 1 0 50508 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_550
timestamp 1586364061
transform 1 0 51704 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_562
timestamp 1586364061
transform 1 0 52808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_574
timestamp 1586364061
transform 1 0 53912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_586
timestamp 1586364061
transform 1 0 55016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_598
timestamp 1586364061
transform 1 0 56120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 57224 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_611
timestamp 1586364061
transform 1 0 57316 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_623
timestamp 1586364061
transform 1 0 58420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_635
timestamp 1586364061
transform 1 0 59524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_647
timestamp 1586364061
transform 1 0 60628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_659
timestamp 1586364061
transform 1 0 61732 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 62836 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_672
timestamp 1586364061
transform 1 0 62928 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_684
timestamp 1586364061
transform 1 0 64032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_696
timestamp 1586364061
transform 1 0 65136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_708
timestamp 1586364061
transform 1 0 66240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_720
timestamp 1586364061
transform 1 0 67344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 68448 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_733
timestamp 1586364061
transform 1 0 68540 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_745
timestamp 1586364061
transform 1 0 69644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_757
timestamp 1586364061
transform 1 0 70748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_769
timestamp 1586364061
transform 1 0 71852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_781
timestamp 1586364061
transform 1 0 72956 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 74060 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_794
timestamp 1586364061
transform 1 0 74152 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_806
timestamp 1586364061
transform 1 0 75256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_818
timestamp 1586364061
transform 1 0 76360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_830
timestamp 1586364061
transform 1 0 77464 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 79672 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_842
timestamp 1586364061
transform 1 0 78568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_855
timestamp 1586364061
transform 1 0 79764 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_867
timestamp 1586364061
transform 1 0 80868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_879
timestamp 1586364061
transform 1 0 81972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_891
timestamp 1586364061
transform 1 0 83076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_903
timestamp 1586364061
transform 1 0 84180 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 85284 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_916
timestamp 1586364061
transform 1 0 85376 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_928
timestamp 1586364061
transform 1 0 86480 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_940
timestamp 1586364061
transform 1 0 87584 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_952
timestamp 1586364061
transform 1 0 88688 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 90896 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_964
timestamp 1586364061
transform 1 0 89792 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_977
timestamp 1586364061
transform 1 0 90988 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_989
timestamp 1586364061
transform 1 0 92092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1001
timestamp 1586364061
transform 1 0 93196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1013
timestamp 1586364061
transform 1 0 94300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1025
timestamp 1586364061
transform 1 0 95404 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 96508 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_1038
timestamp 1586364061
transform 1 0 96600 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1050
timestamp 1586364061
transform 1 0 97704 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1062
timestamp 1586364061
transform 1 0 98808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1074
timestamp 1586364061
transform 1 0 99912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1086
timestamp 1586364061
transform 1 0 101016 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 102120 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_1099
timestamp 1586364061
transform 1 0 102212 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1111
timestamp 1586364061
transform 1 0 103316 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_1123
timestamp 1586364061
transform 1 0 104420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_1135
timestamp 1586364061
transform 1 0 105524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 106812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_1143
timestamp 1586364061
transform 1 0 106260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_94
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_118
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 15364 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_156
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_249
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 26772 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_273
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_280
timestamp 1586364061
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_292
timestamp 1586364061
transform 1 0 27968 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 29624 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_304
timestamp 1586364061
transform 1 0 29072 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_311
timestamp 1586364061
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_323
timestamp 1586364061
transform 1 0 30820 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_335
timestamp 1586364061
transform 1 0 31924 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 32476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_342
timestamp 1586364061
transform 1 0 32568 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_354
timestamp 1586364061
transform 1 0 33672 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 35328 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_366
timestamp 1586364061
transform 1 0 34776 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 38180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_397
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_404
timestamp 1586364061
transform 1 0 38272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_416
timestamp 1586364061
transform 1 0 39376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_428
timestamp 1586364061
transform 1 0 40480 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 41032 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_435
timestamp 1586364061
transform 1 0 41124 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_447
timestamp 1586364061
transform 1 0 42228 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_459
timestamp 1586364061
transform 1 0 43332 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 43884 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_466
timestamp 1586364061
transform 1 0 43976 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_478
timestamp 1586364061
transform 1 0 45080 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 46736 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_490
timestamp 1586364061
transform 1 0 46184 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_497
timestamp 1586364061
transform 1 0 46828 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_509
timestamp 1586364061
transform 1 0 47932 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 49588 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_521
timestamp 1586364061
transform 1 0 49036 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_528
timestamp 1586364061
transform 1 0 49680 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_540
timestamp 1586364061
transform 1 0 50784 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_552
timestamp 1586364061
transform 1 0 51888 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 52440 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_559
timestamp 1586364061
transform 1 0 52532 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_571
timestamp 1586364061
transform 1 0 53636 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_583
timestamp 1586364061
transform 1 0 54740 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 55292 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_590
timestamp 1586364061
transform 1 0 55384 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_602
timestamp 1586364061
transform 1 0 56488 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 58144 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_614
timestamp 1586364061
transform 1 0 57592 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_621
timestamp 1586364061
transform 1 0 58236 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_633
timestamp 1586364061
transform 1 0 59340 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 60996 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_645
timestamp 1586364061
transform 1 0 60444 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_652
timestamp 1586364061
transform 1 0 61088 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_664
timestamp 1586364061
transform 1 0 62192 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_676
timestamp 1586364061
transform 1 0 63296 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 63848 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_683
timestamp 1586364061
transform 1 0 63940 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_695
timestamp 1586364061
transform 1 0 65044 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 66700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_707
timestamp 1586364061
transform 1 0 66148 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_714
timestamp 1586364061
transform 1 0 66792 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_726
timestamp 1586364061
transform 1 0 67896 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 69552 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_738
timestamp 1586364061
transform 1 0 69000 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_745
timestamp 1586364061
transform 1 0 69644 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_757
timestamp 1586364061
transform 1 0 70748 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 72404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_769
timestamp 1586364061
transform 1 0 71852 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_776
timestamp 1586364061
transform 1 0 72496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_788
timestamp 1586364061
transform 1 0 73600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_800
timestamp 1586364061
transform 1 0 74704 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 75256 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_807
timestamp 1586364061
transform 1 0 75348 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_819
timestamp 1586364061
transform 1 0 76452 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 78108 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_831
timestamp 1586364061
transform 1 0 77556 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_838
timestamp 1586364061
transform 1 0 78200 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_850
timestamp 1586364061
transform 1 0 79304 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 80960 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_862
timestamp 1586364061
transform 1 0 80408 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_869
timestamp 1586364061
transform 1 0 81052 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_881
timestamp 1586364061
transform 1 0 82156 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 83812 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_893
timestamp 1586364061
transform 1 0 83260 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_900
timestamp 1586364061
transform 1 0 83904 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_912
timestamp 1586364061
transform 1 0 85008 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_924
timestamp 1586364061
transform 1 0 86112 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 86664 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_931
timestamp 1586364061
transform 1 0 86756 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_943
timestamp 1586364061
transform 1 0 87860 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 89516 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_955
timestamp 1586364061
transform 1 0 88964 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_962
timestamp 1586364061
transform 1 0 89608 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_974
timestamp 1586364061
transform 1 0 90712 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 92368 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_986
timestamp 1586364061
transform 1 0 91816 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_993
timestamp 1586364061
transform 1 0 92460 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1005
timestamp 1586364061
transform 1 0 93564 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 95220 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_1017
timestamp 1586364061
transform 1 0 94668 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_1024
timestamp 1586364061
transform 1 0 95312 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1036
timestamp 1586364061
transform 1 0 96416 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_1048
timestamp 1586364061
transform 1 0 97520 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 98072 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_1055
timestamp 1586364061
transform 1 0 98164 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1067
timestamp 1586364061
transform 1 0 99268 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 100924 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_1079
timestamp 1586364061
transform 1 0 100372 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_1086
timestamp 1586364061
transform 1 0 101016 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1098
timestamp 1586364061
transform 1 0 102120 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 103776 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_1110
timestamp 1586364061
transform 1 0 103224 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_1117
timestamp 1586364061
transform 1 0 103868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_1129
timestamp 1586364061
transform 1 0 104972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_1141
timestamp 1586364061
transform 1 0 106076 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 106812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_1145
timestamp 1586364061
transform 1 0 106444 0 -1 11424
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 3408 480 3528 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 5720 480 5840 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 8032 480 8152 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 10344 480 10464 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 12656 480 12776 6 data_in
port 4 nsew default input
rlabel metal3 s 0 1096 480 1216 6 enable
port 5 nsew default input
rlabel metal2 s 6734 0 6790 480 6 gfpga_pad_GPIO_PAD[0]
port 6 nsew default bidirectional
rlabel metal2 s 20166 0 20222 480 6 gfpga_pad_GPIO_PAD[1]
port 7 nsew default bidirectional
rlabel metal2 s 33690 0 33746 480 6 gfpga_pad_GPIO_PAD[2]
port 8 nsew default bidirectional
rlabel metal2 s 47214 0 47270 480 6 gfpga_pad_GPIO_PAD[3]
port 9 nsew default bidirectional
rlabel metal2 s 60738 0 60794 480 6 gfpga_pad_GPIO_PAD[4]
port 10 nsew default bidirectional
rlabel metal2 s 74170 0 74226 480 6 gfpga_pad_GPIO_PAD[5]
port 11 nsew default bidirectional
rlabel metal2 s 87694 0 87750 480 6 gfpga_pad_GPIO_PAD[6]
port 12 nsew default bidirectional
rlabel metal2 s 101218 0 101274 480 6 gfpga_pad_GPIO_PAD[7]
port 13 nsew default bidirectional
rlabel metal2 s 3330 13520 3386 14000 6 top_width_0_height_0__pin_0_
port 14 nsew default input
rlabel metal2 s 70766 13520 70822 14000 6 top_width_0_height_0__pin_10_
port 15 nsew default input
rlabel metal2 s 77574 13520 77630 14000 6 top_width_0_height_0__pin_11_
port 16 nsew default tristate
rlabel metal2 s 84290 13520 84346 14000 6 top_width_0_height_0__pin_12_
port 17 nsew default input
rlabel metal2 s 91006 13520 91062 14000 6 top_width_0_height_0__pin_13_
port 18 nsew default tristate
rlabel metal2 s 97814 13520 97870 14000 6 top_width_0_height_0__pin_14_
port 19 nsew default input
rlabel metal2 s 104530 13520 104586 14000 6 top_width_0_height_0__pin_15_
port 20 nsew default tristate
rlabel metal2 s 10046 13520 10102 14000 6 top_width_0_height_0__pin_1_
port 21 nsew default tristate
rlabel metal2 s 16762 13520 16818 14000 6 top_width_0_height_0__pin_2_
port 22 nsew default input
rlabel metal2 s 23570 13520 23626 14000 6 top_width_0_height_0__pin_3_
port 23 nsew default tristate
rlabel metal2 s 30286 13520 30342 14000 6 top_width_0_height_0__pin_4_
port 24 nsew default input
rlabel metal2 s 37002 13520 37058 14000 6 top_width_0_height_0__pin_5_
port 25 nsew default tristate
rlabel metal2 s 43810 13520 43866 14000 6 top_width_0_height_0__pin_6_
port 26 nsew default input
rlabel metal2 s 50526 13520 50582 14000 6 top_width_0_height_0__pin_7_
port 27 nsew default tristate
rlabel metal2 s 57334 13520 57390 14000 6 top_width_0_height_0__pin_8_
port 28 nsew default input
rlabel metal2 s 64050 13520 64106 14000 6 top_width_0_height_0__pin_9_
port 29 nsew default tristate
rlabel metal4 s 18944 2128 19264 11472 6 vpwr
port 30 nsew default input
rlabel metal4 s 36944 2128 37264 11472 6 vgnd
port 31 nsew default input
<< end >>
